* NGSPICE file created from wishbone_nn.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt wishbone_nn vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XANTENNA__0674__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold340 _0992_/Q vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _1042_/Q vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _0653_/X vssd1 vssd1 vccd1 vccd1 _0943_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0422__B _0424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0849__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 _0627_/X vssd1 vssd1 vccd1 vccd1 _0918_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _0821_/X vssd1 vssd1 vccd1 vccd1 _1086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _0559_/X vssd1 vssd1 vccd1 vccd1 _0855_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0584__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0985_ _1017_/CLK _0985_/D vssd1 vssd1 vccd1 vccd1 _0985_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout127 _1076_/Q vssd1 vssd1 vccd1 vccd1 _0546_/S1 sky130_fd_sc_hd__buf_4
X_0419_ _0419_/A _0419_/B _0419_/C _0419_/D vssd1 vssd1 vccd1 vccd1 _0424_/B sky130_fd_sc_hd__or4_2
XANTENNA__0669__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 _0850_/S vssd1 vssd1 vccd1 vccd1 _0580_/S sky130_fd_sc_hd__buf_8
Xfanout105 _0836_/S vssd1 vssd1 vccd1 vccd1 _0827_/S sky130_fd_sc_hd__buf_8
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold170 _0748_/X vssd1 vssd1 vccd1 vccd1 _1036_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0579__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 _1025_/Q vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _0634_/X vssd1 vssd1 vccd1 vccd1 _0925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0770_ hold512/X hold590/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0968_ _1104_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout125_A _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0899_ _1100_/CLK _0899_/D vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0482__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0822_ hold411/X hold394/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0822_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0772__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0684_ hold432/X hold463/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0753_ _0802_/B _0759_/B vssd1 vssd1 vccd1 vccd1 _0755_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0473__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0682__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1098_ _1098_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0592__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0767__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1021_ _1096_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0805_ input1/X _0809_/C vssd1 vssd1 vccd1 vccd1 _0805_/Y sky130_fd_sc_hd__nor2_1
X_0736_ hold358/X hold267/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0736_/X sky130_fd_sc_hd__mux2_1
X_0598_ hold245/X hold195/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0667_ hold43/X hold23/X _0682_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
XANTENNA__0446__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0677__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0437__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0587__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1109_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ _0901_/Q _0869_/Q _1102_/Q _1064_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0521_/X sky130_fd_sc_hd__mux4_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0452_ _0496_/A _0452_/B vssd1 vssd1 vccd1 vccd1 _0452_/X sky130_fd_sc_hd__and2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _1101_/CLK _1004_/D vssd1 vssd1 vccd1 vccd1 _1004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 _0583_/X vssd1 vssd1 vccd1 vccd1 _0877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _0663_/X vssd1 vssd1 vccd1 vccd1 _0953_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _0776_/X vssd1 vssd1 vccd1 vccd1 _1052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _0883_/Q vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold577 _0998_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
X_0719_ hold370/X hold308/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0719_/X sky130_fd_sc_hd__mux2_1
Xhold566 _1023_/Q vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold555 _1072_/Q vssd1 vssd1 vccd1 vccd1 _0615_/B sky130_fd_sc_hd__buf_1
Xhold588 _0920_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput75 _0484_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 _0524_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput97 _0448_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0780__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0435_ _0434_/X _0433_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0436_/B sky130_fd_sc_hd__mux2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0504_ _0552_/A _0504_/B vssd1 vssd1 vccd1 vccd1 _0504_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0690__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 _0703_/X vssd1 vssd1 vccd1 vccd1 _0992_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _0960_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _1079_/Q vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _0766_/X vssd1 vssd1 vccd1 vccd1 _1042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold396 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input46/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold352 _0919_/Q vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0775__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0984_ _1090_/CLK _0984_/D vssd1 vssd1 vccd1 vccd1 _0984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0685__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 hold561/X vssd1 vssd1 vccd1 vccd1 _0804_/D sky130_fd_sc_hd__buf_6
X_0418_ _0418_/A input9/X _0418_/C _0418_/D vssd1 vssd1 vccd1 vccd1 _0419_/D sky130_fd_sc_hd__or4_1
Xfanout117 _0572_/S vssd1 vssd1 vccd1 vccd1 _0850_/S sky130_fd_sc_hd__buf_8
Xfanout106 _0778_/S vssd1 vssd1 vccd1 vccd1 _0795_/S sky130_fd_sc_hd__buf_8
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold171 _0908_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _1028_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _0579_/X vssd1 vssd1 vccd1 vccd1 _0875_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _0737_/X vssd1 vssd1 vccd1 vccd1 _1025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0549__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0595__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0967_ _1104_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _0967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0898_ _1109_/CLK _0898_/D vssd1 vssd1 vccd1 vccd1 _0898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0428__B _0428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0821_ hold372/X hold291/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0752_ _0759_/B _0802_/B vssd1 vssd1 vccd1 vccd1 _0755_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0683_ _1074_/Q _1073_/Q input1/X _0797_/B vssd1 vssd1 vccd1 vccd1 _0714_/S sky130_fd_sc_hd__or4_4
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097_ _1100_/CLK _1097_/D vssd1 vssd1 vccd1 vccd1 _1097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1020_ _1093_/CLK _1020_/D vssd1 vssd1 vccd1 vccd1 _1020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0783__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0735_ hold566/X hold5/X _0748_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
X_0804_ _0759_/B _0804_/B _0804_/C _0804_/D vssd1 vssd1 vccd1 vccd1 _0809_/C sky130_fd_sc_hd__and4b_2
X_0597_ hold572/X hold198/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0597_/X sky130_fd_sc_hd__mux2_1
X_0666_ hold204/X hold195/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0666_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0693__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkbuf_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__clkbuf_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0778__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0451_ _0450_/X _0449_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0452_/B sky130_fd_sc_hd__mux2_1
X_0520_ _0552_/A _0520_/B vssd1 vssd1 vccd1 vccd1 _0520_/X sky130_fd_sc_hd__and2_1
X_1003_ _1109_/CLK _1003_/D vssd1 vssd1 vccd1 vccd1 _1003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold501 _1014_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_0718_ hold399/X hold375/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0718_/X sky130_fd_sc_hd__mux2_1
Xhold578 _0975_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 input63/X vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__clkbuf_2
Xhold534 _0589_/X vssd1 vssd1 vccd1 vccd1 _0883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _0851_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold556 _0796_/X vssd1 vssd1 vccd1 vccd1 _0797_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _1074_/Q vssd1 vssd1 vccd1 vccd1 _0800_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 _1095_/Q vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0688__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0649_ hold147/X hold163/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0649_/X sky130_fd_sc_hd__mux2_1
Xhold589 _0983_/Q vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0598__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 _0528_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput98 _0452_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
Xoutput76 _0488_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0503_ _0502_/X _0501_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0504_/B sky130_fd_sc_hd__mux2_1
X_0434_ _1007_/Q _0975_/Q _0943_/Q _0911_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0434_/X sky130_fd_sc_hd__mux4_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold320 _0937_/Q vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _0670_/X vssd1 vssd1 vccd1 vccd1 _0960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _0814_/X vssd1 vssd1 vccd1 vccd1 _1079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _0885_/Q vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 input61/X vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__clkbuf_2
Xhold375 input46/X vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__clkbuf_2
Xhold364 _0917_/Q vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _0628_/X vssd1 vssd1 vccd1 vccd1 _0919_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0791__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0983_ _1098_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 _0983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout129 _1075_/Q vssd1 vssd1 vccd1 vccd1 _0482_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout107 _0787_/S vssd1 vssd1 vccd1 vccd1 _0778_/S sky130_fd_sc_hd__buf_8
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0417_ input6/X input5/X input8/X input7/X vssd1 vssd1 vccd1 vccd1 _0419_/C sky130_fd_sc_hd__or4_1
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0494__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold161 _0876_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _0614_/X vssd1 vssd1 vccd1 vccd1 _0908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _0740_/X vssd1 vssd1 vccd1 vccd1 _1028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 input41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _0588_/X vssd1 vssd1 vccd1 vccd1 _0882_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0549__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0485__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0786__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0966_ _1103_/CLK _0966_/D vssd1 vssd1 vccd1 vccd1 _0966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1093_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0897_ _1108_/CLK hold89/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0696__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0444__B _0444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0820_ hold473/X hold407/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0458__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0751_ _0802_/C _0761_/B hold551/X _0811_/A vssd1 vssd1 vccd1 vccd1 _0751_/X sky130_fd_sc_hd__o211a_1
X_0682_ hold173/X hold147/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0682_/X sky130_fd_sc_hd__mux2_1
X_1096_ _1096_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout130_A _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0449__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0949_ _1115_/CLK _0949_/D vssd1 vssd1 vccd1 vccd1 _0949_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0665_ hold444/X hold198/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0734_ hold219/X hold96/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0734_/X sky130_fd_sc_hd__mux2_1
X_0803_ _0759_/B _0804_/B _0804_/C vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0596_ hold427/X hold404/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0596_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1079_ _1111_/CLK _1079_/D vssd1 vssd1 vccd1 vccd1 _1079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ _1011_/Q _0979_/Q _0947_/Q _0915_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0450_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1098_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0794__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1002_ _1107_/CLK hold77/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold502 _0726_/X vssd1 vssd1 vccd1 vccd1 _1014_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0717_ hold465/X hold432/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0717_/X sky130_fd_sc_hd__mux2_1
Xhold579 _1053_/Q vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_0648_ hold101/X hold120/X _0648_/S vssd1 vssd1 vccd1 vccd1 _0648_/X sky130_fd_sc_hd__mux2_1
Xhold568 _0967_/Q vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _0555_/X vssd1 vssd1 vccd1 vccd1 _0851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _0857_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _0770_/X vssd1 vssd1 vccd1 vccd1 _1046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _0797_/X vssd1 vssd1 vccd1 vccd1 _1072_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _0800_/Y vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0579_ hold101/X hold159/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0579_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput88 _0532_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput99 _0456_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
Xoutput77 _0492_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0789__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0502_ _1024_/Q _0992_/Q _0960_/Q _0928_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0502_/X sky130_fd_sc_hd__mux4_1
X_0433_ _0879_/Q _1112_/Q _1080_/Q _1042_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0433_/X sky130_fd_sc_hd__mux4_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0699__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 _1050_/Q vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold321 _0646_/X vssd1 vssd1 vccd1 vccd1 _0937_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _0688_/X vssd1 vssd1 vccd1 vccd1 _0977_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _1027_/Q vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _0619_/X vssd1 vssd1 vccd1 vccd1 _0910_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _1111_/Q vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _0591_/X vssd1 vssd1 vccd1 vccd1 _0885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _0949_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _0626_/X vssd1 vssd1 vccd1 vccd1 _0917_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0982_ _1092_/CLK _0982_/D vssd1 vssd1 vccd1 vccd1 _0982_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout108 _0731_/S vssd1 vssd1 vccd1 vccd1 _0748_/S sky130_fd_sc_hd__buf_8
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0416_ _0416_/A _0416_/B _0416_/C _0416_/D vssd1 vssd1 vccd1 vccd1 _0419_/B sky130_fd_sc_hd__or4_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold162 _0580_/X vssd1 vssd1 vccd1 vccd1 _0876_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0494__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold151 _0990_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _0933_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _0972_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _0907_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 input41/X vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0485__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0896_ _1100_/CLK _0896_/D vssd1 vssd1 vccd1 vccd1 _0896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0965_ _1108_/CLK _0965_/D vssd1 vssd1 vccd1 vccd1 _0965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0681_ hold118/X hold101/X _0681_/S vssd1 vssd1 vccd1 vccd1 _0681_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0458__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0750_ _0802_/C _0804_/B vssd1 vssd1 vccd1 vccd1 _0750_/Y sky130_fd_sc_hd__nand2_1
X_1095_ _1098_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 _1095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0948_ _1111_/CLK _0948_/D vssd1 vssd1 vccd1 vccd1 _0948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout123_A _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0449__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0879_ _1112_/CLK _0879_/D vssd1 vssd1 vccd1 vccd1 _0879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0802_ _0802_/A _0802_/B _0802_/C vssd1 vssd1 vccd1 vccd1 _0804_/C sky130_fd_sc_hd__or3_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0664_ hold507/X hold404/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0733_ hold27/X hold23/X _0748_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0595_ hold537/X hold521/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1078_ _1110_/CLK _1078_/D vssd1 vssd1 vccd1 vccd1 _1078_/Q sky130_fd_sc_hd__dfxtp_1
Xhold22 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0530__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _1106_/CLK _1001_/D vssd1 vssd1 vccd1 vccd1 _1001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0521__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 _0945_/Q vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
X_0578_ hold60/X hold70/X _0580_/S vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
Xhold514 _0915_/Q vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _0561_/X vssd1 vssd1 vccd1 vccd1 _0857_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _1090_/Q vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _1094_/Q vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
X_0716_ _1074_/Q _1073_/Q _0812_/C vssd1 vssd1 vccd1 vccd1 _0747_/S sky130_fd_sc_hd__nor3b_4
X_0647_ hold60/X hold83/X _0649_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
Xhold558 _1073_/Q vssd1 vssd1 vccd1 vccd1 _0615_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _0801_/Y vssd1 vssd1 vccd1 vccd1 _1074_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput89 _0536_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput78 _0496_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0501_ _0896_/Q _0864_/Q _1097_/Q _1059_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0501_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0432_ _0444_/A _0432_/B vssd1 vssd1 vccd1 vccd1 _0432_/X sky130_fd_sc_hd__and2_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold322 _1001_/Q vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _0774_/X vssd1 vssd1 vccd1 vccd1 _1050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 _0775_/X vssd1 vssd1 vccd1 vccd1 _1051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _0888_/Q vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _0659_/X vssd1 vssd1 vccd1 vccd1 _0949_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _0739_/X vssd1 vssd1 vccd1 vccd1 _1027_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _0846_/X vssd1 vssd1 vccd1 vccd1 _1111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _1006_/Q vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _1041_/Q vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _0951_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0810__B1 _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0981_ _1115_/CLK _0981_/D vssd1 vssd1 vccd1 vccd1 _0981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0804__D _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout109 _0747_/S vssd1 vssd1 vccd1 vccd1 _0731_/S sky130_fd_sc_hd__buf_8
X_0415_ _0415_/A _0415_/B input4/X input3/X vssd1 vssd1 vccd1 vccd1 _0419_/A sky130_fd_sc_hd__or4_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0503__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 _0682_/X vssd1 vssd1 vccd1 vccd1 _0972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _0940_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _0613_/X vssd1 vssd1 vccd1 vccd1 _0907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _0701_/X vssd1 vssd1 vccd1 vccd1 _0990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 _1057_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _0642_/X vssd1 vssd1 vccd1 vccd1 _0933_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 _0732_/X vssd1 vssd1 vccd1 vccd1 _1020_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0964_ _1101_/CLK _0964_/D vssd1 vssd1 vccd1 vccd1 _0964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0895_ _1104_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1108_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0680_ hold64/X hold60/X _0682_/S vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__mux2_1
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1094_ _1096_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _1094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0947_ _1084_/CLK _0947_/D vssd1 vssd1 vccd1 vccd1 _0947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0878_ _1111_/CLK _0878_/D vssd1 vssd1 vccd1 vccd1 _0878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout116_A _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _0617_/B hold546/X input1/X vssd1 vssd1 vccd1 vccd1 _0801_/Y sky130_fd_sc_hd__a21oi_1
X_0732_ hold564/X hold195/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0732_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0663_ hold543/X hold521/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0663_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0601__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0594_ hold344/X hold237/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0594_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1077_ _1084_/CLK _1077_/D vssd1 vssd1 vccd1 vccd1 _1077_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0511__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkbuf_2
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0530__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ _1104_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold504 _0655_/X vssd1 vssd1 vccd1 vccd1 _0945_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0715_ hold147/X hold226/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0715_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0521__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold515 _0624_/X vssd1 vssd1 vccd1 vccd1 _0915_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold526 _0825_/X vssd1 vssd1 vccd1 vccd1 _1090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0577_ hold288/X hold303/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0577_/X sky130_fd_sc_hd__mux2_1
X_0646_ hold288/X hold320/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0646_/X sky130_fd_sc_hd__mux2_1
Xhold548 _1038_/Q vssd1 vssd1 vccd1 vccd1 _0802_/B sky130_fd_sc_hd__buf_1
Xhold537 _0889_/Q vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _0798_/X vssd1 vssd1 vccd1 vccd1 _0799_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput79 _0500_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
XFILLER_0_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0431_ _0430_/X _0429_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0432_/B sky130_fd_sc_hd__mux2_1
X_0500_ _0552_/A _0500_/B vssd1 vssd1 vccd1 vccd1 _0500_/X sky130_fd_sc_hd__and2_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 _0899_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _0712_/X vssd1 vssd1 vccd1 vccd1 _1001_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _1026_/Q vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _0765_/X vssd1 vssd1 vccd1 vccd1 _1041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold301 _0981_/Q vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _0661_/X vssd1 vssd1 vccd1 vccd1 _0951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold312 _0952_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _0594_/X vssd1 vssd1 vccd1 vccd1 _0888_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0430__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 _0853_/Q vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_0629_ hold237/X hold588/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0810__A1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0497__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0980_ _1012_/CLK _0980_/D vssd1 vssd1 vccd1 vccd1 _0980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0414_ _0414_/A _0414_/B _0414_/C vssd1 vssd1 vccd1 vccd1 _0424_/A sky130_fd_sc_hd__or3_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold164 _0649_/X vssd1 vssd1 vccd1 vccd1 _0940_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _0939_/Q vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _0929_/Q vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _1115_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 input40/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 input50/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold131 _0781_/X vssd1 vssd1 vccd1 vccd1 _1057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _1045_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0963_ _1100_/CLK _0963_/D vssd1 vssd1 vccd1 vccd1 _0963_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0604__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0894_ _1098_/CLK _0894_/D vssd1 vssd1 vccd1 vccd1 _0894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1093_ _1093_/CLK _1093_/D vssd1 vssd1 vccd1 vccd1 _1093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0877_ _1110_/CLK _0877_/D vssd1 vssd1 vccd1 vccd1 _0877_/Q sky130_fd_sc_hd__dfxtp_1
X_0946_ _1084_/CLK _0946_/D vssd1 vssd1 vccd1 vccd1 _0946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout109_A _0747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0731_ hold262/X hold198/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__mux2_1
X_0800_ _0800_/A _0800_/B vssd1 vssd1 vccd1 vccd1 _0800_/Y sky130_fd_sc_hd__nand2_1
X_0593_ hold391/X hold93/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0593_/X sky130_fd_sc_hd__mux2_1
X_0662_ hold312/X hold237/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1076_ _1084_/CLK _1076_/D vssd1 vssd1 vccd1 vccd1 _1076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0929_ _1025_/CLK _0929_/D vssd1 vssd1 vccd1 vccd1 _0929_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1012_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0702__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold505 _1043_/Q vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
X_0714_ hold101/X hold108/X _0714_/S vssd1 vssd1 vccd1 vccd1 _0714_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0612__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold516 _0947_/Q vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
X_0645_ hold20/X hold35/X _0649_/S vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__mux2_1
Xhold549 _0757_/X vssd1 vssd1 vccd1 vccd1 _1038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _0979_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold538 _0595_/X vssd1 vssd1 vccd1 vccd1 _0889_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0576_ hold20/X hold62/X _0580_/S vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1059_ _1100_/CLK _1059_/D vssd1 vssd1 vccd1 vccd1 _1059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput69 wire120/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0430_ _1006_/Q _0974_/Q _0942_/Q _0910_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0430_/X sky130_fd_sc_hd__mux4_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0607__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold346 _1068_/Q vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _0605_/X vssd1 vssd1 vccd1 vccd1 _0899_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 _0738_/X vssd1 vssd1 vccd1 vccd1 _1026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _0942_/Q vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _1088_/Q vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _0879_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold302 _0692_/X vssd1 vssd1 vccd1 vccd1 _0981_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 _0662_/X vssd1 vssd1 vccd1 vccd1 _0952_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0628_ hold93/X hold352/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0628_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0430__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0559_ hold93/X hold383/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0559_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0497__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0427__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0413_ _0413_/A _0413_/B _0413_/C _0413_/D vssd1 vssd1 vccd1 vccd1 _0414_/C sky130_fd_sc_hd__or4_1
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 _0958_/Q vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold121 _0648_/X vssd1 vssd1 vccd1 vccd1 _0939_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 input40/X vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__clkbuf_2
Xhold132 _1015_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _0638_/X vssd1 vssd1 vccd1 vccd1 _0929_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _0946_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 input50/X vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__clkbuf_2
Xhold187 _0850_/X vssd1 vssd1 vccd1 vccd1 _1115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _0769_/X vssd1 vssd1 vccd1 vccd1 _1045_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0710__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ _1093_/CLK _0962_/D vssd1 vssd1 vccd1 vccd1 _0962_/Q sky130_fd_sc_hd__dfxtp_1
X_0893_ _1096_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0620__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0705__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1092_ _1092_/CLK _1092_/D vssd1 vssd1 vccd1 vccd1 _1092_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1084_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0945_ _1110_/CLK _0945_/D vssd1 vssd1 vccd1 vccd1 _0945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0876_ _1109_/CLK _0876_/D vssd1 vssd1 vccd1 vccd1 _0876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0542__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0435__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0533__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0730_ hold425/X hold404/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0730_/X sky130_fd_sc_hd__mux2_1
X_0661_ hold366/X hold93/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0592_ hold413/X hold394/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1075_ _1084_/CLK _1075_/D vssd1 vssd1 vccd1 vccd1 _1075_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0859_ _1092_/CLK _0859_/D vssd1 vssd1 vccd1 vccd1 _0859_/Q sky130_fd_sc_hd__dfxtp_1
X_0928_ _1061_/CLK _0928_/D vssd1 vssd1 vccd1 vccd1 _0928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0506__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 _0767_/X vssd1 vssd1 vccd1 vccd1 _1043_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0644_ hold2/X hold15/X _0649_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
Xhold528 _0690_/X vssd1 vssd1 vccd1 vccd1 _0979_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 _0657_/X vssd1 vssd1 vccd1 vccd1 _0947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _0985_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_0713_ hold60/X hold76/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__mux2_1
X_0575_ hold2/X hold9/X _0580_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1058_ _1096_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0713__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0623__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold347 _0792_/X vssd1 vssd1 vccd1 vccd1 _1068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 _0873_/Q vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _0896_/Q vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
X_0558_ hold394/X hold409/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0558_/X sky130_fd_sc_hd__mux2_1
Xhold358 _1024_/Q vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
X_0627_ hold394/X hold586/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0627_/X sky130_fd_sc_hd__mux2_1
Xhold336 _1033_/Q vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold325 _0823_/X vssd1 vssd1 vccd1 vccd1 _1088_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _0585_/X vssd1 vssd1 vccd1 vccd1 _0879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0489_ hold37/A hold31/A _1094_/Q hold49/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0489_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0708__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0443__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0412_ _0412_/A _0412_/B _0412_/C _0412_/D vssd1 vssd1 vccd1 vccd1 _0414_/B sky130_fd_sc_hd__or4_1
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0618__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold144 _0926_/Q vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _0727_/X vssd1 vssd1 vccd1 vccd1 _1015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _0668_/X vssd1 vssd1 vccd1 vccd1 _0958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _1102_/Q vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 input58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _0597_/X vssd1 vssd1 vccd1 vccd1 _0891_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold155 _1109_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _0707_/X vssd1 vssd1 vccd1 vccd1 _0996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _1070_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _0656_/X vssd1 vssd1 vccd1 vccd1 _0946_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ _1025_/CLK _0961_/D vssd1 vssd1 vccd1 vccd1 _0961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0892_ _1093_/CLK _0892_/D vssd1 vssd1 vccd1 vccd1 _0892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0721__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1091_ _1091_/CLK _1091_/D vssd1 vssd1 vccd1 vccd1 _1091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0944_ _1113_/CLK _0944_/D vssd1 vssd1 vccd1 vccd1 _0944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0631__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0875_ _1107_/CLK _0875_/D vssd1 vssd1 vccd1 vccd1 _0875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0542__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0533__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0660_ hold487/X hold394/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0660_/X sky130_fd_sc_hd__mux2_1
X_0591_ hold342/X hold291/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0591_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0451__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1074_ _1112_/CLK _1074_/D vssd1 vssd1 vccd1 vccd1 _1074_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0626__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0927_ _1066_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0789_ hold209/X hold243/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0789_/X sky130_fd_sc_hd__mux2_1
X_0858_ _1092_/CLK _0858_/D vssd1 vssd1 vccd1 vccd1 _0858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0506__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0574_ hold209/X hold230/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0574_/X sky130_fd_sc_hd__mux2_1
X_0712_ hold288/X hold322/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0712_/X sky130_fd_sc_hd__mux2_1
X_0643_ hold209/X hold256/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0643_/X sky130_fd_sc_hd__mux2_1
Xhold507 _0954_/Q vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _1011_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _1084_/Q vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0442__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1057_ _1098_/CLK _1057_/D vssd1 vssd1 vccd1 vccd1 _1057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0433__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold315 _0602_/X vssd1 vssd1 vccd1 vccd1 _0896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _0577_/X vssd1 vssd1 vccd1 vccd1 _0873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold326 _1112_/Q vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _0736_/X vssd1 vssd1 vccd1 vccd1 _1024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _0745_/X vssd1 vssd1 vccd1 vccd1 _1033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _1080_/Q vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_0557_ hold291/X hold389/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0626_ hold291/X hold364/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0626_/X sky130_fd_sc_hd__mux2_1
X_1109_ _1109_/CLK _1109_/D vssd1 vssd1 vccd1 vccd1 _1109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0488_ _0496_/A _0488_/B vssd1 vssd1 vccd1 vccd1 _0488_/X sky130_fd_sc_hd__and2_1
XANTENNA__0814__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0724__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0411_ _0411_/A _0411_/B input23/X input22/X vssd1 vssd1 vccd1 vccd1 _0414_/A sky130_fd_sc_hd__or4bb_1
XFILLER_0_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0634__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 _0844_/X vssd1 vssd1 vccd1 vccd1 _1109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _0635_/X vssd1 vssd1 vccd1 vccd1 _0926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _1064_/Q vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _0837_/X vssd1 vssd1 vccd1 vccd1 _1102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 input58/X vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__buf_2
Xhold112 _0862_/Q vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _0894_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 _0868_/Q vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _0794_/X vssd1 vssd1 vccd1 vccd1 _1070_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0609_ hold53/X hold2/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0719__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0960_ _1061_/CLK _0960_/D vssd1 vssd1 vccd1 vccd1 _0960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0891_ _1100_/CLK _0891_/D vssd1 vssd1 vccd1 vccd1 _0891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0629__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0539__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ _1090_/CLK _1090_/D vssd1 vssd1 vccd1 vccd1 _1090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0874_ _1107_/CLK hold71/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
X_0943_ _1112_/CLK _0943_/D vssd1 vssd1 vccd1 vccd1 _0943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0822__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0732__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0590_ hold440/X hold407/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0590_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1073_ _1112_/CLK _1073_/D vssd1 vssd1 vccd1 vccd1 _1073_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0926_ _1025_/CLK _0926_/D vssd1 vssd1 vccd1 vccd1 _0926_/Q sky130_fd_sc_hd__dfxtp_1
X_0857_ _1090_/CLK _0857_/D vssd1 vssd1 vccd1 vccd1 _0857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0642__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0788_ hold81/X hold134/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__mux2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout107_A _0787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0817__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0727__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold508 _0664_/X vssd1 vssd1 vccd1 vccd1 _0954_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0711_ hold20/X hold33/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0442__S1 _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0573_ hold81/X hold128/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0573_/X sky130_fd_sc_hd__mux2_1
Xhold519 _0819_/X vssd1 vssd1 vccd1 vccd1 _1084_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0642_ hold81/X hold140/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0642_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0637__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1056_ _1096_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
X_0909_ _1110_/CLK _0909_/D vssd1 vssd1 vccd1 vccd1 _0909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0433__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0547__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold316 _0905_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _0928_/Q vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 _0969_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0625_ hold407/X hold467/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0625_/X sky130_fd_sc_hd__mux2_1
Xhold327 _0847_/X vssd1 vssd1 vccd1 vccd1 _1112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _0815_/X vssd1 vssd1 vccd1 vccd1 _1080_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0556_ hold407/X hold593/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0556_/X sky130_fd_sc_hd__mux2_1
X_0487_ _0486_/X _0485_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0488_/B sky130_fd_sc_hd__mux2_1
X_1108_ _1108_/CLK _1108_/D vssd1 vssd1 vccd1 vccd1 _1108_/Q sky130_fd_sc_hd__dfxtp_1
X_1039_ _1084_/CLK _1039_/D vssd1 vssd1 vccd1 vccd1 _1039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0830__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0740__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0410_ _0410_/A vssd1 vssd1 vccd1 vccd1 _0422_/A sky130_fd_sc_hd__inv_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0608_ hold277/X hold209/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0608_/X sky130_fd_sc_hd__mux2_1
Xhold179 _0572_/X vssd1 vssd1 vccd1 vccd1 _0868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _0747_/X vssd1 vssd1 vccd1 vccd1 _1035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _0788_/X vssd1 vssd1 vccd1 vccd1 _1064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _1034_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _0914_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold146 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _0566_/X vssd1 vssd1 vccd1 vccd1 _0862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _0600_/X vssd1 vssd1 vccd1 vccd1 _0894_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0538_/X _0537_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0540_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0825__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0560__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0735__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0890_ _1091_/CLK _0890_/D vssd1 vssd1 vccd1 vccd1 _0890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0645__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1110_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0545__S0 _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0555__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0873_ _1106_/CLK _0873_/D vssd1 vssd1 vccd1 vccd1 _0873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0942_ _1113_/CLK _0942_/D vssd1 vssd1 vccd1 vccd1 _0942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0518__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0509__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ _1112_/CLK _1072_/D vssd1 vssd1 vccd1 vccd1 _1072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0787_ hold176/X hold190/X _0787_/S vssd1 vssd1 vccd1 vccd1 _0787_/X sky130_fd_sc_hd__mux2_1
X_0925_ _1017_/CLK _0925_/D vssd1 vssd1 vccd1 vccd1 _0925_/Q sky130_fd_sc_hd__dfxtp_1
X_0856_ _1090_/CLK _0856_/D vssd1 vssd1 vccd1 vccd1 _0856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0833__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0743__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold509 _1078_/Q vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_0641_ hold176/X hold200/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0710_ hold2/X hold7/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
X_0572_ hold176/X hold178/X _0572_/S vssd1 vssd1 vccd1 vccd1 _0572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055_ _1091_/CLK _1055_/D vssd1 vssd1 vccd1 vccd1 _1055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0653__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0908_ _1109_/CLK _0908_/D vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0839_ hold13/X hold2/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XANTENNA__0828__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0563__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0738__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold317 _0611_/X vssd1 vssd1 vccd1 vccd1 _0905_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _0637_/X vssd1 vssd1 vccd1 vccd1 _0928_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 _0679_/X vssd1 vssd1 vccd1 vccd1 _0969_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0624_ hold512/X hold514/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0624_/X sky130_fd_sc_hd__mux2_1
Xhold328 _1016_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0648__S _0648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0486_ _1020_/Q _0988_/Q _0956_/Q _0924_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0486_/X sky130_fd_sc_hd__mux4_1
X_0555_ hold512/X hold523/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0555_/X sky130_fd_sc_hd__mux2_1
X_1107_ _1107_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
X_1038_ _1084_/CLK _1038_/D vssd1 vssd1 vccd1 vccd1 _1038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0558__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0538_ _1033_/Q _1001_/Q _0969_/Q _0937_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0538_/X sky130_fd_sc_hd__mux4_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold169 _1036_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _0993_/Q vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
X_0607_ hold213/X hold81/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0607_/X sky130_fd_sc_hd__mux2_1
Xhold103 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _1010_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _0623_/X vssd1 vssd1 vccd1 vccd1 _0914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold125 _0746_/X vssd1 vssd1 vccd1 vccd1 _1034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 input59/X vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__clkbuf_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0469_ _0888_/Q _0856_/Q _1089_/Q _1051_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0469_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0841__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0661__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0490__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0836__S _0836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0545__S1 _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0571__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0481__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0746__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0941_ _1110_/CLK _0941_/D vssd1 vssd1 vccd1 vccd1 _0941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ _1105_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0656__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0566__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0518__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0454__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1071_ _1109_/CLK _1071_/D vssd1 vssd1 vccd1 vccd1 _1071_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0509__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0924_ _1093_/CLK _0924_/D vssd1 vssd1 vccd1 vccd1 _0924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0786_ hold222/X hold583/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__mux2_1
X_0855_ _1012_/CLK _0855_/D vssd1 vssd1 vccd1 vccd1 _0855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0445__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_0571_ hold222/X hold224/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0571_/X sky130_fd_sc_hd__mux2_1
X_0640_ hold222/X hold228/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1054_ _1092_/CLK _1054_/D vssd1 vssd1 vccd1 vccd1 _1054_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0807__A1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0907_ _1107_/CLK _0907_/D vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0838_ hold239/X hold209/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0838_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout112_A _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0769_ hold104/X hold153/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0769_/X sky130_fd_sc_hd__mux2_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0844__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold318 _0911_/Q vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold307 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
X_0623_ hold104/X hold157/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0623_/X sky130_fd_sc_hd__mux2_1
Xhold329 _0728_/X vssd1 vssd1 vccd1 vccd1 _1016_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0554_ _1073_/Q input1/X _0797_/B _1074_/Q vssd1 vssd1 vccd1 vccd1 _0572_/S sky130_fd_sc_hd__or4b_4
X_1106_ _1106_/CLK _1106_/D vssd1 vssd1 vccd1 vccd1 _1106_/Q sky130_fd_sc_hd__dfxtp_1
X_0485_ _0892_/Q _0860_/Q _1093_/Q _1055_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0485_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0664__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1037_ _1084_/CLK _1037_/D vssd1 vssd1 vccd1 vccd1 _1037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0839__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0574__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold115 _0704_/X vssd1 vssd1 vccd1 vccd1 _0993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 input62/X vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold126 _0965_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_0537_ _0905_/Q _0873_/Q _1106_/Q _1068_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0537_/X sky130_fd_sc_hd__mux4_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold148 _0795_/X vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ hold232/X hold176/X _0606_/S vssd1 vssd1 vccd1 vccd1 _0606_/X sky130_fd_sc_hd__mux2_1
Xhold159 _0875_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0659__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 _0722_/X vssd1 vssd1 vccd1 vccd1 _1010_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0468_ _0496_/A _0468_/B vssd1 vssd1 vccd1 vccd1 _0468_/X sky130_fd_sc_hd__and2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0569__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0479__S _1077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0490__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0481__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 _0768_/X vssd1 vssd1 vccd1 vccd1 _1044_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0940_ _1109_/CLK _0940_/D vssd1 vssd1 vccd1 vccd1 _0940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0871_ _1104_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1106_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0672__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0847__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0454__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1108_/CLK _1070_/D vssd1 vssd1 vccd1 vccd1 _1070_/Q sky130_fd_sc_hd__dfxtp_1
X_0854_ _1114_/CLK _0854_/D vssd1 vssd1 vccd1 vccd1 _0854_/Q sky130_fd_sc_hd__dfxtp_1
X_0923_ _1092_/CLK _0923_/D vssd1 vssd1 vccd1 vccd1 _0923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0785_ hold250/X hold281/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0785_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0445__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0667__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0577__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0570_ hold250/X hold275/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0570_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0487__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ _1091_/CLK _1053_/D vssd1 vssd1 vccd1 vccd1 _1053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0837_ hold122/X hold81/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__mux2_1
X_0906_ _1107_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0768_ hold397/X hold489/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0768_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0699_ hold195/X hold254/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0699_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout105_A _0836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold308 input57/X vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0770__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0622_ hold397/X hold450/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0622_/X sky130_fd_sc_hd__mux2_1
Xhold319 _0620_/X vssd1 vssd1 vccd1 vccd1 _0911_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0484_ _0496_/A _0484_/B vssd1 vssd1 vccd1 vccd1 _0484_/X sky130_fd_sc_hd__and2_1
XFILLER_0_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0553_ _0615_/B _0759_/B _0804_/B vssd1 vssd1 vccd1 vccd1 _0797_/B sky130_fd_sc_hd__nand3_2
X_1105_ _1105_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1036_ _1109_/CLK _1036_/D vssd1 vssd1 vccd1 vccd1 _1036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0680__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0590__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0765__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 _0961_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 _0689_/X vssd1 vssd1 vccd1 vccd1 _0978_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold116 _1083_/Q vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _0882_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _0675_/X vssd1 vssd1 vccd1 vccd1 _0965_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0605_ hold334/X hold222/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0605_/X sky130_fd_sc_hd__mux2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0467_ _0466_/X _0465_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0468_/B sky130_fd_sc_hd__mux2_1
X_0536_ _0552_/A _0536_/B vssd1 vssd1 vccd1 vccd1 _0536_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1019_ _1061_/CLK _1019_/D vssd1 vssd1 vccd1 vccd1 _1019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0675__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0585__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0495__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0519_ _0518_/X _0517_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0520_/B sky130_fd_sc_hd__mux2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold491 _0880_/Q vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold480 _0724_/X vssd1 vssd1 vccd1 vccd1 _1012_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0870_ _1103_/CLK _0870_/D vssd1 vssd1 vccd1 vccd1 _0870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0999_ _1104_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0773__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0922_ _1012_/CLK _0922_/D vssd1 vssd1 vccd1 vccd1 _0922_/Q sky130_fd_sc_hd__dfxtp_1
X_0853_ _1012_/CLK _0853_/D vssd1 vssd1 vccd1 vccd1 _0853_/Q sky130_fd_sc_hd__dfxtp_1
X_0784_ hold86/X hold595/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__mux2_1
Xinput1 wb_rst_i vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0593__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0768__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1052_ _1090_/CLK _1052_/D vssd1 vssd1 vccd1 vccd1 _1052_/Q sky130_fd_sc_hd__dfxtp_1
X_0905_ _1106_/CLK _0905_/D vssd1 vssd1 vccd1 vccd1 _0905_/Q sky130_fd_sc_hd__dfxtp_1
X_0767_ hold457/X hold505/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0767_/X sky130_fd_sc_hd__mux2_1
X_0836_ hold241/X hold176/X _0836_/S vssd1 vssd1 vccd1 vccd1 _0836_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0698_ hold198/X hold252/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0678__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0588__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0621_ hold457/X hold483/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0621_/X sky130_fd_sc_hd__mux2_1
Xhold309 _0686_/X vssd1 vssd1 vccd1 vccd1 _0975_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0483_ _0482_/X _0481_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0484_/B sky130_fd_sc_hd__mux2_1
X_0552_ _0552_/A _0552_/B vssd1 vssd1 vccd1 vccd1 _0552_/X sky130_fd_sc_hd__and2_1
X_1035_ _1109_/CLK _1035_/D vssd1 vssd1 vccd1 vccd1 _1035_/Q sky130_fd_sc_hd__dfxtp_1
X_1104_ _1104_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0819_ hold518/X hold512/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1091_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0781__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0604_ hold264/X hold250/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0604_/X sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold139 _0671_/X vssd1 vssd1 vccd1 vccd1 _0961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _0869_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _0818_/X vssd1 vssd1 vccd1 vccd1 _1083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _0865_/Q vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0466_ _1015_/Q _0983_/Q _0951_/Q _0919_/Q _0804_/D _0482_/S1 vssd1 vssd1 vccd1 vccd1
+ _0466_/X sky130_fd_sc_hd__mux4_1
X_0535_ _0534_/X _0533_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0536_/B sky130_fd_sc_hd__mux2_1
X_1018_ _1091_/CLK _1018_/D vssd1 vssd1 vccd1 vccd1 _1018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0691__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0493__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0776__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0518_ _1028_/Q _0996_/Q _0964_/Q _0932_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0518_/X sky130_fd_sc_hd__mux4_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0686__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0449_ _0883_/Q _0851_/Q _1084_/Q _1046_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0449_/X sky130_fd_sc_hd__mux4_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0466__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 _0651_/X vssd1 vssd1 vccd1 vccd1 _0941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _0982_/Q vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _0586_/X vssd1 vssd1 vccd1 vccd1 _0880_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0596__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0457__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0998_ _1103_/CLK _0998_/D vssd1 vssd1 vccd1 vccd1 _0998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1096_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0921_ _1017_/CLK _0921_/D vssd1 vssd1 vccd1 vccd1 _0921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0783_ hold267/X hold594/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0783_/X sky130_fd_sc_hd__mux2_1
X_0852_ _1091_/CLK _0852_/D vssd1 vssd1 vccd1 vccd1 _0852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1051_ _1090_/CLK _1051_/D vssd1 vssd1 vccd1 vccd1 _1051_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0784__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0904_ _1104_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_0835_ hold273/X hold222/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0835_/X sky130_fd_sc_hd__mux2_1
X_0697_ hold404/X hold419/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0697_/X sky130_fd_sc_hd__mux2_1
X_0766_ hold308/X hold362/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0766_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0694__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0779__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0551_ _0550_/X _0549_/X _1077_/Q vssd1 vssd1 vccd1 vccd1 _0552_/B sky130_fd_sc_hd__mux2_1
X_0620_ hold308/X hold318/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0482_ _1019_/Q _0987_/Q _0955_/Q _0923_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0482_/X sky130_fd_sc_hd__mux4_1
X_1103_ _1103_/CLK _1103_/D vssd1 vssd1 vccd1 vccd1 _1103_/Q sky130_fd_sc_hd__dfxtp_1
X_1034_ _1105_/CLK _1034_/D vssd1 vssd1 vccd1 vccd1 _1034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0749_ _0802_/A _0802_/B _0802_/C _0759_/B _0804_/B vssd1 vssd1 vccd1 vccd1 _0761_/B
+ sky130_fd_sc_hd__o41a_2
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout110_A _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0689__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0818_ hold116/X hold104/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0818_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0599__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 _0971_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _0573_/X vssd1 vssd1 vccd1 vccd1 _0869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0534_ _1032_/Q hold33/A hold29/A hold35/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0534_/X sky130_fd_sc_hd__mux4_1
X_0603_ hold88/X hold86/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
Xhold107 _0569_/X vssd1 vssd1 vccd1 vccd1 _0865_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ _0887_/Q _0855_/Q _1088_/Q _1050_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0465_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1017_ _1017_/CLK _1017_/D vssd1 vssd1 vccd1 vccd1 _1017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0493__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0792__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0517_ _0900_/Q _0868_/Q _1101_/Q _1063_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0517_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0540__B _0540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0448_ _0496_/A _0448_/B vssd1 vssd1 vccd1 vccd1 _0448_/X sky130_fd_sc_hd__and2_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold471 _0980_/Q vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold460 _0631_/X vssd1 vssd1 vccd1 vccd1 _0922_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0466__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _0693_/X vssd1 vssd1 vccd1 vccd1 _0982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _0944_/Q vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0457__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0787__S _0787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0997_ _1107_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 _0997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0697__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold290 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0920_ _1115_/CLK _0920_/D vssd1 vssd1 vccd1 vccd1 _0920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0782_ hold5/X hold41/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
X_0851_ _1017_/CLK _0851_/D vssd1 vssd1 vccd1 vccd1 _0851_/Q sky130_fd_sc_hd__dfxtp_1
Xinput3 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ _1115_/CLK _1050_/D vssd1 vssd1 vccd1 vccd1 _1050_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0834_ hold283/X hold250/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0903_ _1105_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0765_ hold375/X hold377/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0765_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0696_ hold521/X hold539/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0696_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0502__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0550_ _1036_/Q _1004_/Q _0972_/Q _0940_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0550_/X sky130_fd_sc_hd__mux4_1
X_0481_ _0891_/Q _0859_/Q _1092_/Q _1054_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0481_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0795__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1102_ _1108_/CLK _1102_/D vssd1 vssd1 vccd1 vccd1 _1102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1033_ _1106_/CLK _1033_/D vssd1 vssd1 vccd1 vccd1 _1033_/Q sky130_fd_sc_hd__dfxtp_1
X_0817_ hold461/X hold397/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_1
Xinput50 input50/A vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
X_0679_ hold305/X hold288/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0679_/X sky130_fd_sc_hd__mux2_1
X_0748_ hold169/X hold147/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0748_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout103_A _0648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 _1003_/Q vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_0602_ hold314/X hold267/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0602_/X sky130_fd_sc_hd__mux2_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _0681_/X vssd1 vssd1 vccd1 vccd1 _0971_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0464_ _0496_/A _0464_/B vssd1 vssd1 vccd1 vccd1 _0464_/X sky130_fd_sc_hd__and2_1
X_0533_ hold39/A hold62/A hold68/A hold78/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0533_/X sky130_fd_sc_hd__mux4_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1025_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1016_ _1090_/CLK _1016_/D vssd1 vssd1 vccd1 vccd1 _1016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ _0552_/A _0516_/B vssd1 vssd1 vccd1 vccd1 _0516_/X sky130_fd_sc_hd__and2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0447_ _0446_/X _0445_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0448_/B sky130_fd_sc_hd__mux2_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold461 _1082_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _0913_/Q vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _0654_/X vssd1 vssd1 vccd1 vccd1 _0944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _0912_/Q vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _0691_/X vssd1 vssd1 vccd1 vccd1 _0980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ _1101_/CLK _0996_/D vssd1 vssd1 vccd1 vccd1 _0996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 _0676_/X vssd1 vssd1 vccd1 vccd1 _0966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 input65/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0850_ hold104/X hold186/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__mux2_1
X_0781_ hold96/X hold130/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0781_/X sky130_fd_sc_hd__mux2_1
Xinput4 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0979_ _1017_/CLK _0979_/D vssd1 vssd1 vccd1 vccd1 _0979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0902_ _1103_/CLK _0902_/D vssd1 vssd1 vccd1 vccd1 _0902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0833_ hold98/X hold86/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__mux2_1
X_0764_ hold432/X hold436/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0695_ hold237/X hold247/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0695_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0502__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0480_ _0496_/A _0480_/B vssd1 vssd1 vccd1 vccd1 _0480_/X sky130_fd_sc_hd__and2_1
X_1101_ _1101_/CLK _1101_/D vssd1 vssd1 vccd1 vccd1 _1101_/Q sky130_fd_sc_hd__dfxtp_1
X_1032_ _1104_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _1032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0816_ hold497/X hold457/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0816_/X sky130_fd_sc_hd__mux2_1
X_0747_ hold584/X hold101/X _0747_/S vssd1 vssd1 vccd1 vccd1 _0747_/X sky130_fd_sc_hd__mux2_1
Xinput40 input40/A vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput51 hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0678_ hold29/X hold20/X _0682_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold109 _0714_/X vssd1 vssd1 vccd1 vccd1 _1003_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0601_ hold11/X hold5/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0463_ _0462_/X _0461_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0464_/B sky130_fd_sc_hd__mux2_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ _0552_/A _0532_/B vssd1 vssd1 vccd1 vccd1 _0532_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1015_ _1098_/CLK _1015_/D vssd1 vssd1 vccd1 vccd1 _1015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0478__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0464__B _0464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0469__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0515_ _0514_/X _0513_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0446_ _1010_/Q _0978_/Q _0946_/Q _0914_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0446_/X sky130_fd_sc_hd__mux4_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold462 _0817_/X vssd1 vssd1 vccd1 vccd1 _1082_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _0622_/X vssd1 vssd1 vccd1 vccd1 _0913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _1008_/Q vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _0621_/X vssd1 vssd1 vccd1 vccd1 _0912_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _0884_/Q vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _1085_/Q vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1115_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0995_ _1100_/CLK _0995_/D vssd1 vssd1 vccd1 vccd1 _0995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0429_ _0878_/Q _1111_/Q _1079_/Q _1041_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0429_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _0832_/X vssd1 vssd1 vccd1 vccd1 _1097_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _1061_/Q vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _0772_/X vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ hold23/X hold49/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout126_A _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0978_ _1084_/CLK _0978_/D vssd1 vssd1 vccd1 vccd1 _0978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0832_ hold269/X hold267/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0832_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0602__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0901_ _1108_/CLK _0901_/D vssd1 vssd1 vccd1 vccd1 _0901_/Q sky130_fd_sc_hd__dfxtp_1
X_0763_ input1/X _0797_/B _1074_/Q _1073_/Q vssd1 vssd1 vccd1 vccd1 _0787_/S sky130_fd_sc_hd__or4bb_4
X_0694_ hold93/X hold589/X _0698_/S vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1100_ _1100_/CLK _1100_/D vssd1 vssd1 vccd1 vccd1 _1100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1031_ _1104_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0815_ hold348/X hold308/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0815_/X sky130_fd_sc_hd__mux2_1
Xinput30 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _0416_/D sky130_fd_sc_hd__clkbuf_1
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
Xinput41 input41/A vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
X_0746_ hold124/X hold60/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0677_ hold568/X hold2/X _0682_/S vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__mux2_1
XANTENNA__0507__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0600_ hold167/X hold96/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0600_/X sky130_fd_sc_hd__mux2_1
X_0531_ _0530_/X _0529_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0532_/B sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0462_ _1014_/Q _0982_/Q _0950_/Q _0918_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0462_/X sky130_fd_sc_hd__mux4_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1014_ _1092_/CLK _1014_/D vssd1 vssd1 vccd1 vccd1 _1014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0478__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1017_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0729_ hold541/X hold521/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0729_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0469__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0700__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0514_ _1027_/Q _0995_/Q _0963_/Q _0931_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0514_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0610__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ _0882_/Q _1115_/Q _1083_/Q _1045_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0445_/X sky130_fd_sc_hd__mux4_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold430 _0849_/X vssd1 vssd1 vccd1 vccd1 _1114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _1092_/Q vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _0973_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _0858_/Q vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _0590_/X vssd1 vssd1 vccd1 vccd1 _0884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _0820_/X vssd1 vssd1 vccd1 vccd1 _1085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _0720_/X vssd1 vssd1 vccd1 vccd1 _1008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0605__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0994_ _1061_/CLK _0994_/D vssd1 vssd1 vccd1 vccd1 _0994_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0550__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0428_ _0444_/A _0428_/B vssd1 vssd1 vccd1 vccd1 _0428_/X sky130_fd_sc_hd__and2_1
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0515__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0541__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 _0995_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _0860_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 _0785_/X vssd1 vssd1 vccd1 vccd1 _1061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _0930_/Q vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ _1114_/CLK _0977_/D vssd1 vssd1 vccd1 vccd1 _0977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0514__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _1101_/CLK _0900_/D vssd1 vssd1 vccd1 vccd1 _0900_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0505__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0693_ hold394/X hold481/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0762_ _0761_/B _0760_/Y _0761_/Y input1/X vssd1 vssd1 vccd1 vccd1 _0762_/Y sky130_fd_sc_hd__a211oi_1
X_0831_ hold25/X hold5/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0703__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1030_ _1106_/CLK _1030_/D vssd1 vssd1 vccd1 vccd1 _1030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0814_ hold385/X hold375/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0814_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0613__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput31 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _0416_/C sky130_fd_sc_hd__clkbuf_1
Xinput20 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _0412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0745_ hold336/X hold288/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0745_/X sky130_fd_sc_hd__mux2_1
X_0676_ hold279/X hold209/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0676_/X sky130_fd_sc_hd__mux2_1
Xinput42 hold22/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__clkbuf_1
Xinput64 input64/A vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
Xinput53 hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0523__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0530_ hold17/A hold7/A _0967_/Q hold15/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1 vccd1
+ _0530_/X sky130_fd_sc_hd__mux4_1
X_0461_ _0886_/Q _0854_/Q _1087_/Q _1049_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0461_/X sky130_fd_sc_hd__mux4_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0608__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1013_ _1115_/CLK _1013_/D vssd1 vssd1 vccd1 vccd1 _1013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0659_ hold332/X hold291/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0659_/X sky130_fd_sc_hd__mux2_1
X_0728_ hold328/X hold237/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0513_ _0899_/Q _0867_/Q _1100_/Q _1062_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0513_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0444_ _0444_/A _0444_/B vssd1 vssd1 vccd1 vccd1 _0444_/X sky130_fd_sc_hd__and2_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold453 _0562_/X vssd1 vssd1 vccd1 vccd1 _0858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 _0948_/Q vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold420 _0697_/X vssd1 vssd1 vccd1 vccd1 _0986_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold431 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _0859_/Q vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _0827_/X vssd1 vssd1 vccd1 vccd1 _1092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _0684_/X vssd1 vssd1 vccd1 vccd1 _0973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 _1081_/Q vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0711__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0550__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0993_ _1108_/CLK _0993_/D vssd1 vssd1 vccd1 vccd1 _0993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0621__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0427_ _0426_/X _0425_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0428_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0541__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 _0706_/X vssd1 vssd1 vccd1 vccd1 _0995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _1099_/Q vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _0639_/X vssd1 vssd1 vccd1 vccd1 _0930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _0564_/X vssd1 vssd1 vccd1 vccd1 _0860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0531__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 input48/X vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0706__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0976_ _1113_/CLK _0976_/D vssd1 vssd1 vccd1 vccd1 _0976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0514__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0450__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0505__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0830_ hold567/X hold96/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
X_0692_ hold291/X hold301/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0692_/X sky130_fd_sc_hd__mux2_1
X_0761_ _0802_/A _0761_/B vssd1 vssd1 vccd1 vccd1 _0761_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0441__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1105_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _1066_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0813_ hold509/X hold432/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0813_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _0418_/A sky130_fd_sc_hd__clkbuf_1
Xinput32 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _0415_/B sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _0412_/C sky130_fd_sc_hd__clkbuf_1
Xinput43 hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__clkbuf_1
Xinput54 hold19/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0744_ hold571/X hold20/X _0748_/S vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__mux2_1
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
X_0675_ hold126/X hold81/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1089_ _1090_/CLK _1089_/D vssd1 vssd1 vccd1 vccd1 _1089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0714__S _0714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0460_ _0496_/A _0460_/B vssd1 vssd1 vccd1 vccd1 _0460_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ _1012_/CLK _1012_/D vssd1 vssd1 vccd1 vccd1 _1012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0624__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0727_ hold132/X hold93/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0658_ hold442/X hold407/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0658_/X sky130_fd_sc_hd__mux2_1
X_0589_ hold533/X hold512/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0589_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0709__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0443_ _0442_/X _0441_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0444_/B sky130_fd_sc_hd__mux2_1
X_0512_ _0552_/A _0512_/B vssd1 vssd1 vccd1 vccd1 _0512_/X sky130_fd_sc_hd__and2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0619__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 _0563_/X vssd1 vssd1 vccd1 vccd1 _0859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold410 _0558_/X vssd1 vssd1 vccd1 vccd1 _0854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _0950_/Q vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 _1005_/Q vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _1091_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _1047_/Q vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _0658_/X vssd1 vssd1 vccd1 vccd1 _0948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 input35/X vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__clkbuf_2
Xhold498 _0816_/X vssd1 vssd1 vccd1 vccd1 _1081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0439__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _1061_/CLK _0992_/D vssd1 vssd1 vccd1 vccd1 _0992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0426_ _1005_/Q _0973_/Q _0941_/Q _0909_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0426_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold273 _1100_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _0838_/X vssd1 vssd1 vccd1 vccd1 _1103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _1019_/Q vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _0705_/X vssd1 vssd1 vccd1 vccd1 _0994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _0834_/X vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _1089_/Q vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0722__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0632__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0975_ _1112_/CLK _0975_/D vssd1 vssd1 vccd1 vccd1 _0975_/Q sky130_fd_sc_hd__dfxtp_1
X_0409_ input1/X vssd1 vssd1 vccd1 vccd1 _0811_/A sky130_fd_sc_hd__inv_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0450__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0717__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0760_ _0760_/A _0760_/B vssd1 vssd1 vccd1 vccd1 _0760_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0691_ hold407/X hold471/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0691_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0441__S1 _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0627__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0958_ _1098_/CLK _0958_/D vssd1 vssd1 vccd1 vccd1 _0958_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout124_A _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0889_ _1090_/CLK _0889_/D vssd1 vssd1 vccd1 vccd1 _0889_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0447__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput33 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _0415_/A sky130_fd_sc_hd__clkbuf_1
X_0743_ hold17/X hold2/X _0748_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
Xinput44 hold4/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__clkbuf_1
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_1
Xinput11 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _0418_/D sky130_fd_sc_hd__clkbuf_1
Xinput22 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput55 input55/A vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
X_0812_ _1074_/Q _1073_/Q _0812_/C vssd1 vssd1 vccd1 vccd1 _0836_/S sky130_fd_sc_hd__and3_2
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0674_ hold211/X hold176/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1088_ _1115_/CLK _1088_/D vssd1 vssd1 vccd1 vccd1 _1088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0820__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0730__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1113_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1011_ _1017_/CLK _1011_/D vssd1 vssd1 vccd1 vccd1 _1011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0726_ hold501/X hold394/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0726_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0640__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0657_ hold516/X hold512/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0657_/X sky130_fd_sc_hd__mux2_1
X_0588_ hold149/X hold104/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0588_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0815__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0725__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0511_ _0510_/X _0509_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0512_/B sky130_fd_sc_hd__mux2_1
X_0442_ _1009_/Q _0977_/Q _0945_/Q _0913_/Q _0482_/S0 _0546_/S1 vssd1 vssd1 vccd1
+ vccd1 _0442_/X sky130_fd_sc_hd__mux4_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0635__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold411 _1087_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _0845_/X vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _0877_/Q vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
X_0709_ hold209/X hold577/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0709_/X sky130_fd_sc_hd__mux2_1
Xhold488 _0660_/X vssd1 vssd1 vccd1 vccd1 _0950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _0955_/Q vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _0826_/X vssd1 vssd1 vccd1 vccd1 _1091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _0717_/X vssd1 vssd1 vccd1 vccd1 _1005_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _0771_/X vssd1 vssd1 vccd1 vccd1 _1047_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _1113_/Q vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _0718_/X vssd1 vssd1 vccd1 vccd1 _1006_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0455__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0991_ _1066_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0425_ _0877_/Q _1110_/Q _1078_/Q _1040_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0425_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0526__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold285 _0864_/Q vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _0835_/X vssd1 vssd1 vccd1 vccd1 _1100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _0870_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _0987_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _0731_/X vssd1 vssd1 vccd1 vccd1 _1019_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold241 _1101_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _0824_/X vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0517__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput9 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0974_ _1113_/CLK _0974_/D vssd1 vssd1 vccd1 vccd1 _0974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0823__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0690_ hold512/X hold527/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0690_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0733__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0643__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_A _0572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ _1096_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0888_ _1090_/CLK _0888_/D vssd1 vssd1 vccd1 vccd1 _0888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0818__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0728__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0463__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0742_ hold215/X hold209/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0742_/X sky130_fd_sc_hd__mux2_1
X_0673_ hold234/X hold222/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0673_/X sky130_fd_sc_hd__mux2_1
X_0811_ _0811_/A _0811_/B _0811_/C vssd1 vssd1 vccd1 vccd1 _1077_/D sky130_fd_sc_hd__and3_1
Xinput67 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _0804_/B sky130_fd_sc_hd__buf_2
Xinput34 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _0410_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 input45/A vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
Xinput12 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _0418_/C sky130_fd_sc_hd__clkbuf_1
Xinput23 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput56 hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1087_ _1114_/CLK _1087_/D vssd1 vssd1 vccd1 vccd1 _1087_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0638__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1010_ _1084_/CLK _1010_/D vssd1 vssd1 vccd1 vccd1 _1010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0725_ hold360/X hold291/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0656_ hold165/X hold104/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0656_/X sky130_fd_sc_hd__mux2_1
X_0587_ hold446/X hold397/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0831__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold563_A _1077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0510_ _1026_/Q _0994_/Q _0962_/Q _0930_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0510_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0441_ _0881_/Q _1114_/Q _1082_/Q _1044_/Q _0482_/S0 _0546_/S1 vssd1 vssd1 vccd1
+ vccd1 _0441_/X sky130_fd_sc_hd__mux4_1
Xhold1 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0651__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 _1055_/Q vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _1044_/Q vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _0822_/X vssd1 vssd1 vccd1 vccd1 _1087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _0923_/Q vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _1009_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _0665_/X vssd1 vssd1 vccd1 vccd1 _0955_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0639_ hold250/X hold293/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0639_/X sky130_fd_sc_hd__mux2_1
Xhold478 _0848_/X vssd1 vssd1 vccd1 vccd1 _1113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _0916_/Q vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
X_0708_ hold81/X hold570/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
XANTENNA__0826__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0561__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0736__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0990_ _1098_/CLK _0990_/D vssd1 vssd1 vccd1 vccd1 _0990_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0471__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0424_ _0424_/A _0424_/B _0424_/C _0424_/D vssd1 vssd1 vccd1 vccd1 _0444_/A sky130_fd_sc_hd__nor4_2
XANTENNA__0646__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0526__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold231 _0574_/X vssd1 vssd1 vccd1 vccd1 _0870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _0698_/X vssd1 vssd1 vccd1 vccd1 _0987_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold242 _0836_/X vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold220 _0734_/X vssd1 vssd1 vccd1 vccd1 _1022_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 _0568_/X vssd1 vssd1 vccd1 vccd1 _0864_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0462__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 _0866_/Q vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _0898_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _0962_/Q vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0556__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0517__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0453__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0973_ _1110_/CLK _0973_/D vssd1 vssd1 vccd1 vccd1 _0973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0426__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0956_ _1093_/CLK _0956_/D vssd1 vssd1 vccd1 vccd1 _0956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0806__A1 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0887_ _1012_/CLK _0887_/D vssd1 vssd1 vccd1 vccd1 _0887_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput100 _0460_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0834__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0810_ _0809_/B _0809_/C _0809_/A vssd1 vssd1 vccd1 vccd1 _0811_/C sky130_fd_sc_hd__a21o_1
Xinput13 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _0420_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__0744__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0672_ hold297/X hold250/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_we_i vssd1 vssd1 vccd1 vccd1 _0759_/B sky130_fd_sc_hd__clkbuf_4
Xinput46 input46/A vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
Xinput24 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _0420_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0741_ hold90/X hold81/X _0748_/S vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0654__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1086_ _1115_/CLK _1086_/D vssd1 vssd1 vccd1 vccd1 _1086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0939_ _1109_/CLK _0939_/D vssd1 vssd1 vccd1 vccd1 _0939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0829__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0564__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0739__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0655_ hold503/X hold397/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0655_/X sky130_fd_sc_hd__mux2_1
X_0586_ hold491/X hold457/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0586_/X sky130_fd_sc_hd__mux2_1
X_0724_ hold479/X hold407/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0724_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0649__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1069_ _1107_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 _1069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1103_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0559__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0440_ _0444_/A _0440_/B vssd1 vssd1 vccd1 vccd1 _0440_/X sky130_fd_sc_hd__and2_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold413 _0886_/Q vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _0632_/X vssd1 vssd1 vccd1 vccd1 _0923_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _0721_/X vssd1 vssd1 vccd1 vccd1 _1009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold402 _0779_/X vssd1 vssd1 vccd1 vccd1 _1055_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ hold176/X hold575/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0707_/X sky130_fd_sc_hd__mux2_1
Xhold446 _0881_/Q vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _0625_/X vssd1 vssd1 vccd1 vccd1 _0916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold479 _1012_/Q vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_0638_ hold86/X hold142/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0638_/X sky130_fd_sc_hd__mux2_1
Xhold457 input60/X vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__buf_2
X_0569_ hold86/X hold106/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0842__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0423_ _0759_/B input2/X vssd1 vssd1 vccd1 vccd1 _0424_/D sky130_fd_sc_hd__or2_1
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0662__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold243 _1065_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold210 _0709_/X vssd1 vssd1 vccd1 vccd1 _0998_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0462__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold265 _0604_/X vssd1 vssd1 vccd1 vccd1 _0898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _0570_/X vssd1 vssd1 vccd1 vccd1 _0866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _0900_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold254 _0988_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 input49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 input55/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold298 _0672_/X vssd1 vssd1 vccd1 vccd1 _0962_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0837__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0572__S _0572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0453__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0747__S _0747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0972_ _1109_/CLK _0972_/D vssd1 vssd1 vccd1 vccd1 _0972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0657__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0567__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0426__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0886_ _1114_/CLK _0886_/D vssd1 vssd1 vccd1 vccd1 _0886_/Q sky130_fd_sc_hd__dfxtp_1
X_0955_ _1092_/CLK _0955_/D vssd1 vssd1 vccd1 vccd1 _0955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput101 _0464_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0850__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0740_ hold182/X hold176/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__buf_1
Xinput14 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _0413_/B sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _0411_/B sky130_fd_sc_hd__clkbuf_1
X_0671_ hold138/X hold86/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0671_/X sky130_fd_sc_hd__mux2_1
Xinput47 hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__clkbuf_1
Xinput58 input58/A vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1085_ _1111_/CLK _1085_/D vssd1 vssd1 vccd1 vccd1 _1085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0670__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0869_ _1108_/CLK _0869_/D vssd1 vssd1 vccd1 vccd1 _0869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout122_A _1077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0938_ _1105_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0845__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0580__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0723_ hold529/X hold512/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0723_/X sky130_fd_sc_hd__mux2_1
X_0654_ hold493/X hold457/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0654_/X sky130_fd_sc_hd__mux2_1
X_0585_ hold368/X hold308/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0585_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0665__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1068_ _1106_/CLK _1068_/D vssd1 vssd1 vccd1 vccd1 _1068_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0575__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0538__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold414 _0592_/X vssd1 vssd1 vccd1 vccd1 _0886_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 _0587_/X vssd1 vssd1 vccd1 vccd1 _0881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _1040_/Q vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _0941_/Q vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_0706_ hold222/X hold271/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold458 _0687_/X vssd1 vssd1 vccd1 vccd1 _0976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _1018_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
X_0568_ hold267/X hold285/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0568_/X sky130_fd_sc_hd__mux2_1
X_0637_ hold267/X hold338/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0499_ _0498_/X _0497_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0500_/B sky130_fd_sc_hd__mux2_1
XANTENNA__0529__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0424__A _0424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0422_ _0422_/A _0424_/A _0424_/B _0424_/C vssd1 vssd1 vccd1 vccd1 _0422_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold277 _0902_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _0789_/X vssd1 vssd1 vccd1 vccd1 _1065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _0606_/X vssd1 vssd1 vccd1 vccd1 _0900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _0932_/Q vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0699_/X vssd1 vssd1 vccd1 vccd1 _0988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _0964_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 input49/X vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__clkbuf_2
Xhold288 input55/X vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__clkbuf_2
Xhold266 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _1051_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0971_ _1109_/CLK _0971_/D vssd1 vssd1 vccd1 vccd1 _0971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0673__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0848__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0583__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1092_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0954_ _1012_/CLK _0954_/D vssd1 vssd1 vccd1 vccd1 _0954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0885_ _1115_/CLK _0885_/D vssd1 vssd1 vccd1 vccd1 _0885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0668__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0578__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0670_ hold330/X hold267/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0670_/X sky130_fd_sc_hd__mux2_1
Xinput15 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _0413_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 input48/A vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput26 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _0411_/A sky130_fd_sc_hd__clkbuf_1
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1084_ _1084_/CLK _1084_/D vssd1 vssd1 vccd1 vccd1 _1084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0937_ _1106_/CLK _0937_/D vssd1 vssd1 vccd1 vccd1 _0937_/Q sky130_fd_sc_hd__dfxtp_1
X_0868_ _1101_/CLK _0868_/D vssd1 vssd1 vccd1 vccd1 _0868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout115_A _0606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0799_ _0811_/A _0800_/B _0799_/C vssd1 vssd1 vccd1 vccd1 _0799_/X sky130_fd_sc_hd__and3_1
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0771__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0653_ hold350/X hold308/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0653_/X sky130_fd_sc_hd__mux2_1
X_0722_ hold136/X hold104/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0722_/X sky130_fd_sc_hd__mux2_1
X_0584_ hold415/X hold375/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0584_/X sky130_fd_sc_hd__mux2_1
X_1067_ _1105_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0681__S _0681_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0591__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1066_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0538__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0766__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold437 _0764_/X vssd1 vssd1 vccd1 vccd1 _1040_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _0909_/Q vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
X_0705_ hold250/X hold573/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0705_/X sky130_fd_sc_hd__mux2_1
Xhold426 _0730_/X vssd1 vssd1 vccd1 vccd1 _1018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _0878_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _0922_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_0636_ hold5/X hold57/X _0649_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
XANTENNA__0474__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 input39/X vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0676__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0498_ _1023_/Q hold66/A hold51/A hold57/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0498_/X sky130_fd_sc_hd__mux4_1
X_0567_ hold5/X hold47/X _0580_/S vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__mux2_1
XANTENNA__0529__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0465__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold561_A _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0586__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0421_ input1/X _0421_/B _0804_/B vssd1 vssd1 vccd1 vccd1 _0424_/C sky130_fd_sc_hd__or3b_1
Xhold201 _0641_/X vssd1 vssd1 vccd1 vccd1 _0932_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 _0786_/X vssd1 vssd1 vccd1 vccd1 _1062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _0841_/X vssd1 vssd1 vccd1 vccd1 _1106_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _0608_/X vssd1 vssd1 vccd1 vccd1 _0902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _0934_/Q vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _0963_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _0892_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _0674_/X vssd1 vssd1 vccd1 vccd1 _0964_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0619_ hold375/X hold581/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0619_/X sky130_fd_sc_hd__mux2_1
Xhold267 input45/X vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__buf_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0438__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ _1107_/CLK hold65/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0429__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0774__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0884_ _1091_/CLK _0884_/D vssd1 vssd1 vccd1 vccd1 _0884_/Q sky130_fd_sc_hd__dfxtp_1
X_0953_ _1017_/CLK _0953_/D vssd1 vssd1 vccd1 vccd1 _0953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0684__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0594__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _0413_/D sky130_fd_sc_hd__clkbuf_1
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _0420_/B sky130_fd_sc_hd__clkbuf_1
Xinput49 input49/A vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0769__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1083_ _1084_/CLK _1083_/D vssd1 vssd1 vccd1 vccd1 _1083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0936_ _1104_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0867_ _1100_/CLK _0867_/D vssd1 vssd1 vccd1 vccd1 _0867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0679__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout108_A _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0798_ _0615_/B _0759_/B _0804_/B _0615_/A vssd1 vssd1 vccd1 vccd1 _0798_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0589__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0721_ hold423/X hold397/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0721_/X sky130_fd_sc_hd__mux2_1
X_0583_ hold499/X hold432/X _0597_/S vssd1 vssd1 vccd1 vccd1 _0583_/X sky130_fd_sc_hd__mux2_1
X_0652_ hold379/X hold375/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0652_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0499__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_1066_ _1066_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0919_ _1090_/CLK _0919_/D vssd1 vssd1 vccd1 vccd1 _0919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkbuf_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0782__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold438 _1054_/Q vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _0618_/X vssd1 vssd1 vccd1 vccd1 _0909_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 _0890_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _0777_/X vssd1 vssd1 vccd1 vccd1 _1053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _0584_/X vssd1 vssd1 vccd1 vccd1 _0878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0704_ hold86/X hold114/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0704_/X sky130_fd_sc_hd__mux2_1
X_0635_ hold96/X hold144/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0635_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0474__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0566_ hold96/X hold112/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0566_/X sky130_fd_sc_hd__mux2_1
X_0497_ hold11/A hold47/A hold25/A hold41/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0497_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1049_ _1114_/CLK _1049_/D vssd1 vssd1 vccd1 vccd1 _1049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0692__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0465__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0420_ _0420_/A _0420_/B _0420_/C vssd1 vssd1 vccd1 vccd1 _0421_/B sky130_fd_sc_hd__or3_1
XANTENNA__0777__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold224 _0867_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _0673_/X vssd1 vssd1 vccd1 vccd1 _0963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 _0924_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _0901_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold268 _0783_/X vssd1 vssd1 vccd1 vccd1 _1059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _0966_/Q vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _0643_/X vssd1 vssd1 vccd1 vccd1 _0934_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0618_ hold432/X hold448/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0549_ _0908_/Q _0876_/Q _1109_/Q _1071_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0549_/X sky130_fd_sc_hd__mux4_1
Xhold246 _0598_/X vssd1 vssd1 vccd1 vccd1 _0892_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0687__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0438__S1 _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0597__S _0597_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0429__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0790__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0952_ _1115_/CLK _0952_/D vssd1 vssd1 vccd1 vccd1 _0952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0883_ _1017_/CLK _0883_/D vssd1 vssd1 vccd1 vccd1 _0883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0510__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1101_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0501__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
Xinput17 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _0413_/C sky130_fd_sc_hd__clkbuf_1
Xinput28 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _0416_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0785__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1082_ _1114_/CLK _1082_/D vssd1 vssd1 vccd1 vccd1 _1082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0866_ _1101_/CLK _0866_/D vssd1 vssd1 vccd1 vccd1 _0866_/Q sky130_fd_sc_hd__dfxtp_1
X_0935_ _1104_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_0797_ _0811_/A _0797_/B _0797_/C vssd1 vssd1 vccd1 vccd1 _0797_/X sky130_fd_sc_hd__and3_1
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0695__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0720_ hold495/X hold457/X _0731_/S vssd1 vssd1 vccd1 vccd1 _0720_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0651_ hold469/X hold432/X _0665_/S vssd1 vssd1 vccd1 vccd1 _0651_/X sky130_fd_sc_hd__mux2_1
X_0582_ _1073_/Q _0812_/C _1074_/Q vssd1 vssd1 vccd1 vccd1 _0606_/S sky130_fd_sc_hd__and3b_2
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0809__A _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0528__B _0528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1065_ _1103_/CLK _1065_/D vssd1 vssd1 vccd1 vccd1 _1065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0849_ hold397/X hold429/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0849_/X sky130_fd_sc_hd__mux2_1
X_0918_ _1114_/CLK _0918_/D vssd1 vssd1 vccd1 vccd1 _0918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _1049_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
X_0703_ hold267/X hold340/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0703_/X sky130_fd_sc_hd__mux2_1
Xhold406 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input64/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold439 _0778_/X vssd1 vssd1 vccd1 vccd1 _1054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _0596_/X vssd1 vssd1 vccd1 vccd1 _0890_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0634_ hold23/X hold180/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0634_/X sky130_fd_sc_hd__mux2_1
X_0496_ _0496_/A _0496_/B vssd1 vssd1 vccd1 vccd1 _0496_/X sky130_fd_sc_hd__and2_1
X_0565_ hold23/X hold31/X _0580_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1048_ _1115_/CLK _1048_/D vssd1 vssd1 vccd1 vccd1 _1048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0793__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 _0571_/X vssd1 vssd1 vccd1 vccd1 _0867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _1097_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _0607_/X vssd1 vssd1 vccd1 vccd1 _0901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _0633_/X vssd1 vssd1 vccd1 vccd1 _0924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _0984_/Q vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _0856_/Q vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0479_ _0478_/X _0477_/X _1077_/Q vssd1 vssd1 vccd1 vccd1 _0480_/B sky130_fd_sc_hd__mux2_1
X_0548_ _0552_/A _0548_/B vssd1 vssd1 vccd1 vccd1 _0548_/X sky130_fd_sc_hd__and2_1
X_0617_ input1/X _0617_/B vssd1 vssd1 vccd1 vccd1 _0648_/S sky130_fd_sc_hd__or2_4
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0788__S _0795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0698__S _0698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0951_ _1090_/CLK _0951_/D vssd1 vssd1 vccd1 vccd1 _0951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0882_ _1115_/CLK _0882_/D vssd1 vssd1 vccd1 vccd1 _0882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0510__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _0412_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0501__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _0416_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1081_ _1113_/CLK _1081_/D vssd1 vssd1 vccd1 vccd1 _1081_/Q sky130_fd_sc_hd__dfxtp_1
X_0934_ _1103_/CLK _0934_/D vssd1 vssd1 vccd1 vccd1 _0934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0865_ _1025_/CLK _0865_/D vssd1 vssd1 vccd1 vccd1 _0865_/Q sky130_fd_sc_hd__dfxtp_1
X_0796_ _0759_/B _0804_/B _0615_/B vssd1 vssd1 vccd1 vccd1 _0796_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0486__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0581_ _1072_/Q _0759_/B _0804_/B _0811_/A vssd1 vssd1 vccd1 vccd1 _0812_/C sky130_fd_sc_hd__and4b_1
X_0650_ _1074_/Q _1073_/Q _0812_/C vssd1 vssd1 vccd1 vccd1 _0681_/S sky130_fd_sc_hd__and3b_2
X_1064_ _1108_/CLK _1064_/D vssd1 vssd1 vccd1 vccd1 _1064_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0809__B _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1112_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0477__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0779_ hold195/X hold401/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0779_/X sky130_fd_sc_hd__mux2_1
X_0848_ hold457/X hold477/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0848_/X sky130_fd_sc_hd__mux2_1
X_0917_ _1115_/CLK _0917_/D vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout113_A _0681_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold418 _0773_/X vssd1 vssd1 vccd1 vccd1 _1049_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold429 _1114_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0633_ hold195/X hold202/X _0649_/S vssd1 vssd1 vccd1 vccd1 _0633_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 input64/X vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__clkbuf_2
X_0702_ hold5/X hold66/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0564_ hold195/X hold260/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0495_ _0494_/X _0493_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1047_ _1111_/CLK _1047_/D vssd1 vssd1 vccd1 vccd1 _1047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 _1030_/Q vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold226 _1004_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _0956_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 input37/X vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold248 _0695_/X vssd1 vssd1 vccd1 vccd1 _0984_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0616_ _0800_/A _0800_/B vssd1 vssd1 vccd1 vccd1 _0617_/B sky130_fd_sc_hd__or2_1
Xhold259 _0560_/X vssd1 vssd1 vccd1 vccd1 _0856_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0478_ _1018_/Q _0986_/Q _0954_/Q _0922_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0478_/X sky130_fd_sc_hd__mux4_1
X_0547_ _0546_/X _0545_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold590 _1046_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0881_ _1114_/CLK _0881_/D vssd1 vssd1 vccd1 vccd1 _0881_/Q sky130_fd_sc_hd__dfxtp_1
X_0950_ _1091_/CLK _0950_/D vssd1 vssd1 vccd1 vccd1 _0950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _0412_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1090_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1080_ _1112_/CLK _1080_/D vssd1 vssd1 vccd1 vccd1 _1080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0864_ _1100_/CLK _0864_/D vssd1 vssd1 vccd1 vccd1 _0864_/Q sky130_fd_sc_hd__dfxtp_1
X_0795_ hold147/X hold592/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0795_/X sky130_fd_sc_hd__mux2_1
X_0933_ _1105_/CLK _0933_/D vssd1 vssd1 vccd1 vccd1 _0933_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout130 _1075_/Q vssd1 vssd1 vccd1 vccd1 _0542_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0486__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0580_ hold147/X hold161/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1063_ _1101_/CLK _1063_/D vssd1 vssd1 vccd1 vccd1 _1063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0477__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0916_ _1111_/CLK _0916_/D vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0778_ hold198/X hold438/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0778_/X sky130_fd_sc_hd__mux2_1
X_0847_ hold308/X hold326/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0847_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout106_A _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_0563_ hold198/X hold475/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0563_/X sky130_fd_sc_hd__mux2_1
X_0632_ hold198/X hold434/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0632_/X sky130_fd_sc_hd__mux2_1
Xhold408 _0556_/X vssd1 vssd1 vccd1 vccd1 _0852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _0986_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_0701_ hold96/X hold151/X _0715_/S vssd1 vssd1 vccd1 vccd1 _0701_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0494_ _1022_/Q _0990_/Q _0958_/Q _0926_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0494_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0600__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1046_ _1084_/CLK _1046_/D vssd1 vssd1 vccd1 vccd1 _1046_/Q sky130_fd_sc_hd__dfxtp_1
X_1115_ _1115_/CLK _1115_/D vssd1 vssd1 vccd1 vccd1 _1115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold216 _0742_/X vssd1 vssd1 vccd1 vccd1 _1030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _0715_/X vssd1 vssd1 vccd1 vccd1 _1004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _0666_/X vssd1 vssd1 vccd1 vccd1 _0956_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0546_ _1035_/Q _1003_/Q _0971_/Q _0939_/Q _1075_/Q _0546_/S1 vssd1 vssd1 vccd1 vccd1
+ _0546_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold249 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input48/A sky130_fd_sc_hd__dlygate4sd3_1
X_0615_ _0615_/A _0615_/B _0759_/B _0804_/B vssd1 vssd1 vccd1 vccd1 _0800_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold238 _0629_/X vssd1 vssd1 vccd1 vccd1 _0920_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0477_ _0890_/Q _0858_/Q _1091_/Q _1053_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0477_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1029_ _1107_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0522__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ hold53/A hold9/A hold13/A hold55/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1 vccd1
+ _0529_/X sky130_fd_sc_hd__mux4_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0513__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 _1069_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _0978_/Q vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0880_ _1113_/CLK _0880_/D vssd1 vssd1 vccd1 vccd1 _0880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ _1101_/CLK _0932_/D vssd1 vssd1 vccd1 vccd1 _0932_/Q sky130_fd_sc_hd__dfxtp_1
X_0794_ hold101/X hold188/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0794_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0863_ _1066_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0603__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout131 _1075_/Q vssd1 vssd1 vccd1 vccd1 _0550_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_14_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1062_ _1100_/CLK _1062_/D vssd1 vssd1 vccd1 vccd1 _1062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0915_ _1084_/CLK _0915_/D vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0777_ hold404/X hold579/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0777_/X sky130_fd_sc_hd__mux2_1
X_0846_ hold375/X hold387/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ hold23/X hold45/X _0715_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
Xhold409 _0854_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
X_0562_ hold404/X hold452/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0562_/X sky130_fd_sc_hd__mux2_1
X_0631_ hold404/X hold459/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0631_/X sky130_fd_sc_hd__mux2_1
X_1114_ _1114_/CLK _1114_/D vssd1 vssd1 vccd1 vccd1 _1114_/Q sky130_fd_sc_hd__dfxtp_1
X_0493_ _0894_/Q _0862_/Q _1095_/Q _1057_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0493_/X sky130_fd_sc_hd__mux4_1
X_1045_ _1112_/CLK _1045_/D vssd1 vssd1 vccd1 vccd1 _1045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0829_ hold569/X hold23/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0701__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 _1093_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 _1108_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 _1103_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0611__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold228 _0931_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_0614_ hold171/X hold147/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0614_/X sky130_fd_sc_hd__mux2_1
X_0545_ _0907_/Q _0875_/Q _1108_/Q _1070_/Q _1075_/Q _0546_/S1 vssd1 vssd1 vccd1 vccd1
+ _0545_/X sky130_fd_sc_hd__mux4_1
X_0476_ _0496_/A _0476_/B vssd1 vssd1 vccd1 vccd1 _0476_/X sky130_fd_sc_hd__and2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1028_ _1101_/CLK _1028_/D vssd1 vssd1 vccd1 vccd1 _1028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1107_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0431__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0606__S _0606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0522__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0459_ _0458_/X _0457_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0460_/B sky130_fd_sc_hd__mux2_1
X_0528_ _0552_/A _0528_/B vssd1 vssd1 vccd1 vccd1 _0528_/X sky130_fd_sc_hd__and2_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0513__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 _1071_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _0910_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _0997_/Q vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput90 _0540_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout129_A _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0498__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0931_ _1100_/CLK _0931_/D vssd1 vssd1 vccd1 vccd1 _0931_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0489__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0862_ _1098_/CLK _0862_/D vssd1 vssd1 vccd1 vccd1 _0862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0793_ hold60/X hold580/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout121 hold563/X vssd1 vssd1 vccd1 vccd1 _0809_/A sky130_fd_sc_hd__buf_8
Xfanout110 _0698_/S vssd1 vssd1 vccd1 vccd1 _0715_/S sky130_fd_sc_hd__buf_6
XANTENNA__0484__B _0484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0704__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1061_ _1061_/CLK _1061_/D vssd1 vssd1 vccd1 vccd1 _1061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0845_ hold432/X hold585/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0845_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0614__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0914_ _1084_/CLK _0914_/D vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dfxtp_1
X_0776_ hold521/X hold574/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0776_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0492_ _0496_/A _0492_/B vssd1 vssd1 vccd1 vccd1 _0492_/X sky130_fd_sc_hd__and2_1
X_0630_ hold521/X hold531/X _0632_/S vssd1 vssd1 vccd1 vccd1 _0630_/X sky130_fd_sc_hd__mux2_1
Xmax_cap118 _0496_/A vssd1 vssd1 vccd1 vccd1 _0552_/A sky130_fd_sc_hd__clkbuf_4
X_0561_ hold521/X hold535/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0561_/X sky130_fd_sc_hd__mux2_1
X_1044_ _1110_/CLK _1044_/D vssd1 vssd1 vccd1 vccd1 _1044_/Q sky130_fd_sc_hd__dfxtp_1
X_1113_ _1113_/CLK _1113_/D vssd1 vssd1 vccd1 vccd1 _1113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0609__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0828_ hold206/X hold195/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0828_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout111_A _0714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0759_ _0802_/A _0759_/B vssd1 vssd1 vccd1 vccd1 _0760_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0519__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold229 _0640_/X vssd1 vssd1 vccd1 vccd1 _0931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold207 _0828_/X vssd1 vssd1 vccd1 vccd1 _1093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 _0843_/X vssd1 vssd1 vccd1 vccd1 _1108_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0613_ hold184/X hold101/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0613_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0475_ _0474_/X _0473_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0476_/B sky130_fd_sc_hd__mux2_1
X_0544_ _0552_/A _0544_/B vssd1 vssd1 vccd1 vccd1 _0544_/X sky130_fd_sc_hd__and2_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ _1103_/CLK _1027_/D vssd1 vssd1 vccd1 vccd1 _1027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0712__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0622__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0527_ _0526_/X _0525_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0528_/B sky130_fd_sc_hd__mux2_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0458_ _1013_/Q _0981_/Q _0949_/Q _0917_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0458_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold582 _0977_/Q vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _0852_/Q vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _1032_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold560 _0799_/X vssd1 vssd1 vccd1 vccd1 _1073_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0707__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 _0504_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput91 _0544_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1111_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0527__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0498__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold390 _0557_/X vssd1 vssd1 vccd1 vccd1 _0853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0792_ hold288/X hold346/X _0795_/S vssd1 vssd1 vccd1 vccd1 _0792_/X sky130_fd_sc_hd__mux2_1
X_0930_ _1093_/CLK _0930_/D vssd1 vssd1 vccd1 vccd1 _0930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0489__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0861_ _1096_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout111 _0714_/S vssd1 vssd1 vccd1 vccd1 _0698_/S sky130_fd_sc_hd__buf_8
Xfanout122 _1077_/Q vssd1 vssd1 vccd1 vccd1 _0547_/S sky130_fd_sc_hd__buf_8
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0720__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1060_ _1098_/CLK hold87/X vssd1 vssd1 vccd1 vccd1 _1060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0913_ _1114_/CLK _0913_/D vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dfxtp_1
X_0844_ hold155/X hold147/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0844_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0630__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0775_ hold237/X hold299/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0715__S _0715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap119 _0444_/A vssd1 vssd1 vccd1 vccd1 _0496_/A sky130_fd_sc_hd__clkbuf_4
X_0491_ _0490_/X _0489_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0492_/B sky130_fd_sc_hd__mux2_1
X_0560_ hold237/X hold258/X _0850_/S vssd1 vssd1 vccd1 vccd1 _0560_/X sky130_fd_sc_hd__mux2_1
X_1043_ _1111_/CLK _1043_/D vssd1 vssd1 vccd1 vccd1 _1043_/Q sky130_fd_sc_hd__dfxtp_1
X_1112_ _1112_/CLK _1112_/D vssd1 vssd1 vccd1 vccd1 _1112_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0625__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0827_ hold485/X hold198/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout104_A _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0758_ _0802_/C _0755_/C _0755_/B vssd1 vssd1 vccd1 vccd1 _0760_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0689_ hold104/X hold591/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0689_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0535__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0534__S0 _0542_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0612_ hold72/X hold60/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__mux2_1
Xhold219 _1022_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold208 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0474_ _1017_/Q _0985_/Q _0953_/Q _0921_/Q _0804_/D _0482_/S1 vssd1 vssd1 vccd1 vccd1
+ _0474_/X sky130_fd_sc_hd__mux4_1
X_0543_ _0542_/X _0541_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0544_/B sky130_fd_sc_hd__mux2_1
XANTENNA__0525__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1026_ _1093_/CLK _1026_/D vssd1 vssd1 vccd1 vccd1 _1026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
X_0526_ _1030_/Q _0998_/Q _0966_/Q _0934_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0526_/X sky130_fd_sc_hd__mux4_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0457_ _0885_/Q _0853_/Q _1086_/Q _1048_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0457_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1009_ _1114_/CLK _1009_/D vssd1 vssd1 vccd1 vccd1 _1009_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0813__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold583 _1062_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _0891_/Q vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _1059_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _1075_/Q vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _1037_/Q vssd1 vssd1 vccd1 vccd1 _0802_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0723__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput70 _0428_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput81 _0432_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput92 _0436_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0633__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0509_ _0898_/Q _0866_/Q _1099_/Q _1061_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0509_/X sky130_fd_sc_hd__mux4_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0543__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold380 _0652_/X vssd1 vssd1 vccd1 vccd1 _0942_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0718__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 _0887_/Q vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0860_ _1093_/CLK _0860_/D vssd1 vssd1 vccd1 vccd1 _0860_/Q sky130_fd_sc_hd__dfxtp_1
X_0791_ hold20/X hold78/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0628__S _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0989_ _1096_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout112 _0665_/S vssd1 vssd1 vccd1 vccd1 _0682_/S sky130_fd_sc_hd__buf_8
Xfanout123 _0482_/S1 vssd1 vssd1 vccd1 vccd1 _0809_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ _1113_/CLK _0912_/D vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0843_ hold217/X hold101/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0843_/X sky130_fd_sc_hd__mux2_1
X_0774_ hold93/X hold310/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0774_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0821__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0731__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0490_ hold27/A hold45/A hold43/A _0925_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0490_/X sky130_fd_sc_hd__mux4_1
X_1111_ _1111_/CLK _1111_/D vssd1 vssd1 vccd1 vccd1 _1111_/Q sky130_fd_sc_hd__dfxtp_1
X_1042_ _1112_/CLK _1042_/D vssd1 vssd1 vccd1 vccd1 _1042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0641__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0688_ hold397/X hold582/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0688_/X sky130_fd_sc_hd__mux2_1
X_0826_ hold421/X hold404/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0826_/X sky130_fd_sc_hd__mux2_1
X_0757_ _0802_/B _0761_/B _0756_/Y _0811_/A vssd1 vssd1 vccd1 vccd1 _0757_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0816__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0551__S _1077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0726__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0534__S1 _0542_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0611_ hold316/X hold288/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0611_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 input52/X vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0542_ _1034_/Q hold76/A hold64/A hold83/A _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0542_/X sky130_fd_sc_hd__mux4_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0473_ _0889_/Q _0857_/Q _1090_/Q _1052_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0473_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0470__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0525__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1025_ _1025_/CLK _1025_/D vssd1 vssd1 vccd1 vccd1 _1025_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0636__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0809_ _0809_/A _0809_/B _0809_/C vssd1 vssd1 vccd1 vccd1 _0811_/B sky130_fd_sc_hd__nand3_1
XANTENNA__0461__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__clkbuf_2
X_0525_ _0902_/Q _0870_/Q _1103_/Q _1065_/Q _0550_/S0 _0550_/S1 vssd1 vssd1 vccd1
+ vccd1 _0525_/X sky130_fd_sc_hd__mux4_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0456_ _0496_/A _0456_/B vssd1 vssd1 vccd1 vccd1 _0456_/X sky130_fd_sc_hd__and2_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1113_/CLK _1008_/D vssd1 vssd1 vccd1 vccd1 _1008_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold540 _0696_/X vssd1 vssd1 vccd1 vccd1 _0985_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _0806_/X vssd1 vssd1 vccd1 vccd1 _1075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _0750_/Y vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _0994_/Q vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _1035_/Q vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0434__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold595 _1060_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0425__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 _0468_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput82 _0508_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput93 _0548_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0439_ _0438_/X _0437_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0440_/B sky130_fd_sc_hd__mux2_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0508_ _0552_/A _0508_/B vssd1 vssd1 vccd1 vccd1 _0508_/X sky130_fd_sc_hd__and2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_8_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0824__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold381 _0974_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _0593_/X vssd1 vssd1 vccd1 vccd1 _0887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _1007_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1100_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0734__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0790_ hold2/X hold55/X _0795_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0988_ _1025_/CLK _0988_/D vssd1 vssd1 vccd1 vccd1 _0988_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0644__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 _0632_/S vssd1 vssd1 vccd1 vccd1 _0649_/S sky130_fd_sc_hd__buf_8
Xfanout113 _0681_/S vssd1 vssd1 vccd1 vccd1 _0665_/S sky130_fd_sc_hd__buf_8
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout124 _0546_/S1 vssd1 vssd1 vccd1 vccd1 _0482_/S1 sky130_fd_sc_hd__buf_6
XANTENNA__0819__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0729__S _0731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0911_ _1112_/CLK _0911_/D vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dfxtp_1
X_0842_ hold74/X hold60/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0773_ hold394/X hold417/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0773_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0639__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1110_/CLK _1110_/D vssd1 vssd1 vccd1 vccd1 _1110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0459__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1041_ _1111_/CLK _1041_/D vssd1 vssd1 vccd1 vccd1 _1041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0825_ hold525/X hold521/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0687_ hold457/X hold576/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0687_/X sky130_fd_sc_hd__mux2_1
X_0756_ _0754_/Y _0755_/X _0761_/B vssd1 vssd1 vccd1 vccd1 _0756_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0832__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0742__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0541_ hold72/A hold70/A hold74/A _1069_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0541_/X sky130_fd_sc_hd__mux4_1
X_0472_ _0496_/A _0472_/B vssd1 vssd1 vccd1 vccd1 _0472_/X sky130_fd_sc_hd__and2_1
X_0610_ hold39/X hold20/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__mux2_1
XANTENNA__0470__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ _1061_/CLK _1024_/D vssd1 vssd1 vccd1 vccd1 _1024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0652__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0808_ _0809_/B _0809_/C _0807_/Y vssd1 vssd1 vccd1 vccd1 _1076_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0461__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0739_ hold354/X hold222/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0827__S _0827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0562__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0737__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__clkbuf_2
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__clkbuf_2
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0455_ _0454_/X _0453_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0456_/B sky130_fd_sc_hd__mux2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0552_/A _0524_/B vssd1 vssd1 vccd1 vccd1 _0524_/X sky130_fd_sc_hd__and2_1
X_1007_ _1112_/CLK _1007_/D vssd1 vssd1 vccd1 vccd1 _1007_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0647__S _0649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold585 _1110_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0434__S1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 _0723_/X vssd1 vssd1 vccd1 vccd1 _1011_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _1077_/Q vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _1017_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _0751_/X vssd1 vssd1 vccd1 vccd1 _1037_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _1052_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0557__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0425__S1 _0482_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput94 _0552_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
Xoutput72 _0472_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput83 _0512_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0467__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0438_ _1008_/Q _0976_/Q _0944_/Q _0912_/Q _0482_/S0 _0546_/S1 vssd1 vssd1 vccd1
+ vccd1 _0438_/X sky130_fd_sc_hd__mux4_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ _0506_/X _0505_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0508_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0840__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 _0685_/X vssd1 vssd1 vccd1 vccd1 _0974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _0719_/X vssd1 vssd1 vccd1 vccd1 _1007_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _1013_/Q vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0987_ _1061_/CLK _0987_/D vssd1 vssd1 vccd1 vccd1 _0987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0660__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 _0648_/S vssd1 vssd1 vccd1 vccd1 _0632_/S sky130_fd_sc_hd__buf_8
Xfanout125 _0546_/S1 vssd1 vssd1 vccd1 vccd1 _0542_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout114 _0597_/S vssd1 vssd1 vccd1 vccd1 _0614_/S sky130_fd_sc_hd__buf_8
XANTENNA__0835__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0570__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 _1063_/Q vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0745__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ hold565/X hold288/X _0844_/S vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__mux2_1
X_0910_ _1113_/CLK _0910_/D vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ hold291/X hold587/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0772_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0655__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0546__S0 _1075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0565__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1040_ _1114_/CLK _1040_/D vssd1 vssd1 vccd1 vccd1 _1040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0537__S0 _0550_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0475__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0755_ _1037_/Q _0755_/B _0755_/C vssd1 vssd1 vccd1 vccd1 _0755_/X sky130_fd_sc_hd__and3_1
X_0824_ hold295/X hold237/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0824_/X sky130_fd_sc_hd__mux2_1
X_0686_ hold308/X hold578/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0686_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire120 _0422_/Y vssd1 vssd1 vccd1 vccd1 wire120/X sky130_fd_sc_hd__buf_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ _0552_/A _0540_/B vssd1 vssd1 vccd1 vccd1 _0540_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0471_ _0470_/X _0469_/X _0809_/A vssd1 vssd1 vccd1 vccd1 _0472_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1023_ _1104_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _1023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_8_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1114_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0738_ hold356/X hold250/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0738_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout102_A _0632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0807_ _0809_/B _0809_/C input1/X vssd1 vssd1 vccd1 vccd1 _0807_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0669_ hold51/X hold5/X _0682_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0843__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0454_ _1012_/Q _0980_/Q _0948_/Q _0916_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0454_/X sky130_fd_sc_hd__mux4_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ _0522_/X _0521_/X _0547_/S vssd1 vssd1 vccd1 vccd1 _0524_/B sky130_fd_sc_hd__mux2_1
X_1006_ _1113_/CLK _1006_/D vssd1 vssd1 vccd1 vccd1 _1006_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0663__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold586 _0918_/Q vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _0996_/Q vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _1020_/Q vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _0921_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold520 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _0729_/X vssd1 vssd1 vccd1 vccd1 _1017_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _1039_/Q vssd1 vssd1 vccd1 vccd1 _0802_/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0838__S _0844_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0573__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0748__S _0748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 _0516_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput95 _0440_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
Xoutput73 _0476_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0483__S _0809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0506_ _1025_/Q _0993_/Q _0961_/Q _0929_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0506_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0437_ _0880_/Q _1113_/Q _1081_/Q _1043_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0437_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0658__S _0665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0568__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold372 _1086_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _0855_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 input66/X vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__clkbuf_2
Xhold361 _0725_/X vssd1 vssd1 vccd1 vccd1 _1013_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 _0943_/Q vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1104_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0986_ _1091_/CLK _0986_/D vssd1 vssd1 vccd1 vccd1 _0986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout126 _0546_/S1 vssd1 vssd1 vccd1 vccd1 _0550_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout104 _0827_/S vssd1 vssd1 vccd1 vccd1 _0844_/S sky130_fd_sc_hd__buf_8
Xfanout115 _0606_/S vssd1 vssd1 vccd1 vccd1 _0597_/S sky130_fd_sc_hd__buf_8
XFILLER_0_64_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 _0925_/Q vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold191 _0787_/X vssd1 vssd1 vccd1 vccd1 _1063_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0771_ hold407/X hold454/X _0778_/S vssd1 vssd1 vccd1 vccd1 _0771_/X sky130_fd_sc_hd__mux2_1
X_0840_ hold68/X hold20/X _0844_/S vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0671__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0969_ _1106_/CLK _0969_/D vssd1 vssd1 vccd1 vccd1 _0969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0846__S _0850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0546__S1 _0546_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0482__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0537__S1 _0550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0491__S _0547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0685_ hold375/X hold381/X _0698_/S vssd1 vssd1 vccd1 vccd1 _0685_/X sky130_fd_sc_hd__mux2_1
X_0823_ hold324/X hold93/X _0827_/S vssd1 vssd1 vccd1 vccd1 _0823_/X sky130_fd_sc_hd__mux2_1
X_0754_ _0755_/B _0755_/C _1037_/Q vssd1 vssd1 vccd1 vccd1 _0754_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__0473__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1099_ _1101_/CLK _1099_/D vssd1 vssd1 vccd1 vccd1 _1099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0666__S _0682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0576__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0470_ _1016_/Q _0984_/Q _0952_/Q _0920_/Q _0804_/D _0809_/B vssd1 vssd1 vccd1 vccd1
+ _0470_/X sky130_fd_sc_hd__mux4_1
X_1022_ _1025_/CLK _1022_/D vssd1 vssd1 vccd1 vccd1 _1022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0737_ hold192/X hold86/X _0748_/S vssd1 vssd1 vccd1 vccd1 _0737_/X sky130_fd_sc_hd__mux2_1
X_0668_ hold110/X hold96/X _0682_/S vssd1 vssd1 vccd1 vccd1 _0668_/X sky130_fd_sc_hd__mux2_1
X_0806_ _0804_/D _0803_/X _0805_/Y vssd1 vssd1 vccd1 vccd1 _0806_/X sky130_fd_sc_hd__o21a_1
XANTENNA__0446__S0 _0804_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0599_ hold37/X hold23/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0437__S0 _0482_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0522_ hold90/A _0997_/Q _0965_/Q _0933_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0522_/X sky130_fd_sc_hd__mux4_1
X_0453_ _0884_/Q _0852_/Q _1085_/Q _1047_/Q _0482_/S0 _0482_/S1 vssd1 vssd1 vccd1
+ vccd1 _0453_/X sky130_fd_sc_hd__mux4_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _1110_/CLK _1005_/D vssd1 vssd1 vccd1 vccd1 _1005_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0808__A1 _0809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 _0813_/X vssd1 vssd1 vccd1 vccd1 _1078_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold565 _1106_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _0976_/Q vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _1048_/Q vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 input38/X vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__clkbuf_2
Xhold543 _0953_/Q vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _0630_/X vssd1 vssd1 vccd1 vccd1 _0921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _0762_/Y vssd1 vssd1 vccd1 vccd1 _1039_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput85 _0520_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput96 _0444_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
Xoutput74 _0480_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0764__S _0778_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0436_ _0444_/A _0436_/B vssd1 vssd1 vccd1 vccd1 _0436_/X sky130_fd_sc_hd__and2_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0505_ hold88/A _0865_/Q hold98/A _1060_/Q _0542_/S0 _0542_/S1 vssd1 vssd1 vccd1
+ vccd1 _0505_/X sky130_fd_sc_hd__mux4_1
.ends

