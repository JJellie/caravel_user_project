magic
tech sky130A
magscale 1 2
timestamp 1726655002
<< viali >>
rect 37013 21505 37047 21539
rect 5641 21437 5675 21471
rect 9505 21437 9539 21471
rect 12173 21437 12207 21471
rect 12909 21437 12943 21471
rect 15393 21437 15427 21471
rect 18613 21437 18647 21471
rect 27813 21437 27847 21471
rect 28641 21437 28675 21471
rect 30757 21437 30791 21471
rect 33425 21437 33459 21471
rect 37841 21437 37875 21471
rect 38669 21437 38703 21471
rect 40509 21437 40543 21471
rect 43269 21437 43303 21471
rect 44005 21437 44039 21471
rect 44189 21437 44223 21471
rect 46121 21437 46155 21471
rect 48237 21437 48271 21471
rect 49157 21437 49191 21471
rect 53389 21437 53423 21471
rect 56609 21437 56643 21471
rect 36369 21369 36403 21403
rect 37289 21369 37323 21403
rect 47133 21369 47167 21403
rect 52009 21369 52043 21403
rect 4997 21301 5031 21335
rect 5917 21301 5951 21335
rect 8677 21301 8711 21335
rect 8953 21301 8987 21335
rect 11529 21301 11563 21335
rect 12265 21301 12299 21335
rect 14841 21301 14875 21335
rect 18061 21301 18095 21335
rect 22109 21301 22143 21335
rect 24869 21301 24903 21335
rect 27261 21301 27295 21335
rect 28089 21301 28123 21335
rect 30297 21301 30331 21335
rect 31401 21301 31435 21335
rect 32413 21301 32447 21335
rect 33977 21301 34011 21335
rect 34437 21301 34471 21335
rect 38025 21301 38059 21335
rect 39037 21301 39071 21335
rect 39957 21301 39991 21335
rect 42717 21301 42751 21335
rect 43453 21301 43487 21335
rect 44833 21301 44867 21335
rect 45845 21301 45879 21335
rect 46765 21301 46799 21335
rect 47593 21301 47627 21335
rect 48513 21301 48547 21335
rect 52837 21301 52871 21335
rect 53849 21301 53883 21335
rect 55965 21301 55999 21335
rect 56057 21301 56091 21335
rect 5825 21097 5859 21131
rect 12173 21097 12207 21131
rect 18797 21097 18831 21131
rect 27077 21097 27111 21131
rect 27261 21097 27295 21131
rect 35633 21097 35667 21131
rect 39865 21097 39899 21131
rect 45937 21097 45971 21131
rect 49341 21097 49375 21131
rect 56057 21097 56091 21131
rect 10701 21029 10735 21063
rect 15301 21029 15335 21063
rect 24409 21029 24443 21063
rect 30389 21029 30423 21063
rect 36553 21029 36587 21063
rect 43729 21029 43763 21063
rect 4905 20961 4939 20995
rect 5181 20961 5215 20995
rect 8217 20961 8251 20995
rect 8401 20961 8435 20995
rect 14657 20961 14691 20995
rect 15393 20961 15427 20995
rect 17693 20961 17727 20995
rect 18337 20961 18371 20995
rect 24225 20961 24259 20995
rect 24961 20961 24995 20995
rect 27813 20961 27847 20995
rect 30297 20961 30331 20995
rect 31033 20961 31067 20995
rect 36461 20961 36495 20995
rect 37105 20961 37139 20995
rect 37473 20961 37507 20995
rect 37657 20961 37691 20995
rect 39221 20961 39255 20995
rect 46489 20961 46523 20995
rect 46949 20961 46983 20995
rect 48789 20961 48823 20995
rect 49617 20961 49651 20995
rect 52285 20961 52319 20995
rect 52469 20961 52503 20995
rect 54401 20961 54435 20995
rect 55413 20961 55447 20995
rect 56701 20961 56735 20995
rect 4629 20893 4663 20927
rect 6561 20893 6595 20927
rect 6929 20893 6963 20927
rect 9137 20893 9171 20927
rect 10149 20893 10183 20927
rect 10793 20893 10827 20927
rect 12817 20893 12851 20927
rect 13553 20893 13587 20927
rect 14933 20893 14967 20927
rect 19809 20893 19843 20927
rect 20085 20893 20119 20927
rect 22109 20893 22143 20927
rect 22845 20893 22879 20927
rect 23489 20893 23523 20927
rect 25237 20893 25271 20927
rect 25881 20893 25915 20927
rect 27629 20893 27663 20927
rect 28641 20893 28675 20927
rect 31861 20893 31895 20927
rect 34253 20893 34287 20927
rect 35265 20893 35299 20927
rect 36921 20893 36955 20927
rect 41245 20893 41279 20927
rect 41889 20893 41923 20927
rect 42349 20893 42383 20927
rect 42616 20893 42650 20927
rect 44373 20893 44407 20927
rect 46305 20893 46339 20927
rect 46397 20893 46431 20927
rect 47133 20893 47167 20927
rect 48145 20893 48179 20927
rect 50721 20893 50755 20927
rect 51457 20893 51491 20927
rect 53573 20893 53607 20927
rect 55597 20893 55631 20927
rect 56977 20893 57011 20927
rect 57529 20893 57563 20927
rect 5365 20825 5399 20859
rect 5917 20825 5951 20859
rect 11060 20825 11094 20859
rect 13001 20825 13035 20859
rect 18153 20825 18187 20859
rect 20352 20825 20386 20859
rect 22293 20825 22327 20859
rect 24777 20825 24811 20859
rect 27721 20825 27755 20859
rect 30757 20825 30791 20859
rect 32597 20825 32631 20859
rect 34008 20825 34042 20859
rect 38945 20825 38979 20859
rect 41000 20825 41034 20859
rect 41337 20825 41371 20859
rect 47041 20825 47075 20859
rect 47593 20825 47627 20859
rect 48881 20825 48915 20859
rect 50169 20825 50203 20859
rect 56517 20825 56551 20859
rect 4261 20757 4295 20791
rect 4721 20757 4755 20791
rect 5457 20757 5491 20791
rect 7757 20757 7791 20791
rect 8125 20757 8159 20791
rect 9781 20757 9815 20791
rect 12265 20757 12299 20791
rect 14381 20757 14415 20791
rect 14841 20757 14875 20791
rect 16037 20757 16071 20791
rect 17785 20757 17819 20791
rect 18245 20757 18279 20791
rect 19257 20757 19291 20791
rect 21465 20757 21499 20791
rect 21557 20757 21591 20791
rect 23581 20757 23615 20791
rect 24869 20757 24903 20791
rect 28089 20757 28123 20791
rect 29009 20757 29043 20791
rect 29653 20757 29687 20791
rect 30849 20757 30883 20791
rect 31217 20757 31251 20791
rect 32137 20757 32171 20791
rect 32873 20757 32907 20791
rect 34713 20757 34747 20791
rect 35817 20757 35851 20791
rect 37013 20757 37047 20791
rect 37749 20757 37783 20791
rect 38117 20757 38151 20791
rect 38485 20757 38519 20791
rect 38577 20757 38611 20791
rect 39037 20757 39071 20791
rect 39681 20757 39715 20791
rect 43821 20757 43855 20791
rect 44833 20757 44867 20791
rect 45201 20757 45235 20791
rect 45753 20757 45787 20791
rect 47501 20757 47535 20791
rect 48973 20757 49007 20791
rect 50905 20757 50939 20791
rect 51917 20757 51951 20791
rect 52561 20757 52595 20791
rect 52929 20757 52963 20791
rect 53021 20757 53055 20791
rect 53757 20757 53791 20791
rect 55045 20757 55079 20791
rect 55689 20757 55723 20791
rect 56149 20757 56183 20791
rect 56609 20757 56643 20791
rect 6929 20553 6963 20587
rect 8861 20553 8895 20587
rect 10977 20553 11011 20587
rect 11805 20553 11839 20587
rect 14657 20553 14691 20587
rect 18613 20553 18647 20587
rect 18981 20553 19015 20587
rect 21833 20553 21867 20587
rect 24869 20553 24903 20587
rect 28365 20553 28399 20587
rect 28457 20553 28491 20587
rect 29745 20553 29779 20587
rect 31585 20553 31619 20587
rect 31953 20553 31987 20587
rect 37105 20553 37139 20587
rect 39957 20553 39991 20587
rect 40049 20553 40083 20587
rect 40417 20553 40451 20587
rect 43821 20553 43855 20587
rect 47317 20553 47351 20587
rect 57161 20553 57195 20587
rect 4804 20485 4838 20519
rect 15792 20485 15826 20519
rect 17408 20485 17442 20519
rect 27252 20485 27286 20519
rect 28825 20485 28859 20519
rect 30880 20485 30914 20519
rect 37473 20485 37507 20519
rect 42708 20485 42742 20519
rect 46204 20485 46238 20519
rect 50660 20485 50694 20519
rect 51448 20485 51482 20519
rect 53113 20485 53147 20519
rect 56048 20485 56082 20519
rect 8585 20417 8619 20451
rect 9985 20417 10019 20451
rect 10241 20417 10275 20451
rect 11897 20417 11931 20451
rect 13507 20417 13541 20451
rect 14381 20417 14415 20451
rect 16037 20417 16071 20451
rect 17141 20417 17175 20451
rect 20520 20417 20554 20451
rect 21557 20417 21591 20451
rect 22201 20417 22235 20451
rect 22661 20417 22695 20451
rect 23745 20417 23779 20451
rect 25605 20417 25639 20451
rect 25881 20417 25915 20451
rect 26617 20417 26651 20451
rect 26801 20417 26835 20451
rect 29653 20417 29687 20451
rect 31125 20417 31159 20451
rect 31493 20417 31527 20451
rect 32965 20417 32999 20451
rect 33977 20417 34011 20451
rect 34161 20417 34195 20451
rect 34621 20417 34655 20451
rect 35725 20417 35759 20451
rect 35992 20417 36026 20451
rect 38393 20417 38427 20451
rect 39405 20417 39439 20451
rect 45845 20417 45879 20451
rect 48375 20417 48409 20451
rect 49433 20417 49467 20451
rect 54652 20417 54686 20451
rect 55781 20417 55815 20451
rect 3893 20349 3927 20383
rect 4537 20349 4571 20383
rect 7573 20349 7607 20383
rect 7711 20349 7745 20383
rect 7849 20349 7883 20383
rect 8769 20349 8803 20383
rect 10793 20349 10827 20383
rect 10885 20349 10919 20383
rect 11621 20349 11655 20383
rect 13369 20349 13403 20383
rect 13645 20349 13679 20383
rect 14565 20349 14599 20383
rect 19073 20349 19107 20383
rect 19165 20349 19199 20383
rect 20363 20349 20397 20383
rect 20637 20349 20671 20383
rect 21373 20349 21407 20383
rect 22293 20349 22327 20383
rect 22385 20349 22419 20383
rect 23213 20349 23247 20383
rect 23489 20349 23523 20383
rect 25764 20349 25798 20383
rect 26985 20349 27019 20383
rect 28917 20349 28951 20383
rect 29009 20349 29043 20383
rect 31401 20349 31435 20383
rect 33103 20349 33137 20383
rect 33241 20349 33275 20383
rect 33517 20349 33551 20383
rect 34437 20349 34471 20383
rect 34529 20349 34563 20383
rect 38531 20349 38565 20383
rect 38669 20349 38703 20383
rect 38945 20349 38979 20383
rect 39589 20349 39623 20383
rect 39773 20349 39807 20383
rect 42441 20349 42475 20383
rect 45937 20349 45971 20383
rect 48237 20349 48271 20383
rect 48513 20349 48547 20383
rect 49249 20349 49283 20383
rect 50905 20349 50939 20383
rect 51181 20349 51215 20383
rect 52837 20349 52871 20383
rect 53021 20349 53055 20383
rect 54493 20349 54527 20383
rect 54769 20349 54803 20383
rect 55505 20349 55539 20383
rect 55689 20349 55723 20383
rect 5917 20281 5951 20315
rect 8125 20281 8159 20315
rect 11345 20281 11379 20315
rect 13921 20281 13955 20315
rect 18521 20281 18555 20315
rect 20913 20281 20947 20315
rect 26157 20281 26191 20315
rect 35265 20281 35299 20315
rect 48789 20281 48823 20315
rect 52561 20281 52595 20315
rect 53481 20281 53515 20315
rect 55045 20281 55079 20315
rect 4445 20213 4479 20247
rect 12265 20213 12299 20247
rect 12633 20213 12667 20247
rect 12725 20213 12759 20247
rect 19717 20213 19751 20247
rect 24961 20213 24995 20247
rect 32321 20213 32355 20247
rect 34989 20213 35023 20247
rect 37749 20213 37783 20247
rect 41429 20213 41463 20247
rect 44557 20213 44591 20247
rect 47593 20213 47627 20247
rect 49525 20213 49559 20247
rect 53849 20213 53883 20247
rect 5641 20009 5675 20043
rect 8677 20009 8711 20043
rect 10517 20009 10551 20043
rect 12265 20009 12299 20043
rect 14105 20009 14139 20043
rect 19257 20009 19291 20043
rect 21741 20009 21775 20043
rect 23581 20009 23615 20043
rect 25237 20009 25271 20043
rect 27721 20009 27755 20043
rect 29009 20009 29043 20043
rect 31217 20009 31251 20043
rect 33977 20009 34011 20043
rect 34713 20009 34747 20043
rect 37473 20009 37507 20043
rect 39865 20009 39899 20043
rect 42717 20009 42751 20043
rect 43913 20009 43947 20043
rect 46765 20009 46799 20043
rect 49525 20009 49559 20043
rect 51457 20009 51491 20043
rect 53941 20009 53975 20043
rect 56701 20009 56735 20043
rect 56793 20009 56827 20043
rect 5549 19941 5583 19975
rect 9689 19941 9723 19975
rect 13001 19941 13035 19975
rect 18521 19941 18555 19975
rect 31125 19941 31159 19975
rect 39405 19941 39439 19975
rect 42165 19941 42199 19975
rect 43729 19941 43763 19975
rect 7297 19873 7331 19907
rect 9137 19873 9171 19907
rect 9873 19873 9907 19907
rect 17141 19873 17175 19907
rect 20361 19873 20395 19907
rect 21925 19873 21959 19907
rect 24961 19873 24995 19907
rect 28365 19873 28399 19907
rect 31769 19873 31803 19907
rect 36093 19873 36127 19907
rect 40417 19873 40451 19907
rect 41797 19873 41831 19907
rect 43361 19873 43395 19907
rect 44557 19873 44591 19907
rect 47501 19873 47535 19907
rect 50721 19873 50755 19907
rect 51549 19873 51583 19907
rect 53573 19873 53607 19907
rect 57345 19873 57379 19907
rect 4169 19805 4203 19839
rect 6285 19805 6319 19839
rect 9321 19805 9355 19839
rect 10885 19805 10919 19839
rect 15485 19805 15519 19839
rect 16129 19805 16163 19839
rect 19901 19805 19935 19839
rect 20628 19805 20662 19839
rect 23489 19805 23523 19839
rect 24225 19805 24259 19839
rect 25789 19805 25823 19839
rect 26341 19805 26375 19839
rect 26608 19805 26642 19839
rect 29745 19805 29779 19839
rect 32597 19805 32631 19839
rect 35265 19805 35299 19839
rect 37749 19805 37783 19839
rect 38025 19805 38059 19839
rect 42533 19805 42567 19839
rect 43177 19805 43211 19839
rect 44281 19805 44315 19839
rect 45293 19805 45327 19839
rect 45385 19805 45419 19839
rect 48145 19805 48179 19839
rect 49801 19805 49835 19839
rect 55137 19805 55171 19839
rect 55321 19805 55355 19839
rect 4436 19737 4470 19771
rect 7564 19737 7598 19771
rect 11152 19737 11186 19771
rect 15240 19737 15274 19771
rect 17408 19737 17442 19771
rect 19073 19737 19107 19771
rect 24869 19737 24903 19771
rect 29990 19737 30024 19771
rect 32864 19737 32898 19771
rect 36360 19737 36394 19771
rect 38292 19737 38326 19771
rect 45652 19737 45686 19771
rect 48412 19737 48446 19771
rect 51816 19737 51850 19771
rect 53021 19737 53055 19771
rect 55588 19737 55622 19771
rect 9229 19669 9263 19703
rect 12541 19669 12575 19703
rect 15577 19669 15611 19703
rect 20177 19669 20211 19703
rect 22569 19669 22603 19703
rect 24409 19669 24443 19703
rect 24777 19669 24811 19703
rect 32137 19669 32171 19703
rect 34345 19669 34379 19703
rect 35633 19669 35667 19703
rect 43085 19669 43119 19703
rect 44373 19669 44407 19703
rect 46857 19669 46891 19703
rect 47869 19669 47903 19703
rect 50169 19669 50203 19703
rect 52929 19669 52963 19703
rect 54309 19669 54343 19703
rect 7665 19465 7699 19499
rect 9873 19465 9907 19499
rect 14565 19465 14599 19499
rect 15761 19465 15795 19499
rect 17601 19465 17635 19499
rect 22109 19465 22143 19499
rect 24869 19465 24903 19499
rect 33701 19465 33735 19499
rect 34069 19465 34103 19499
rect 37289 19465 37323 19499
rect 38761 19465 38795 19499
rect 39681 19465 39715 19499
rect 48973 19465 49007 19499
rect 49525 19465 49559 19499
rect 55597 19465 55631 19499
rect 55873 19465 55907 19499
rect 22201 19397 22235 19431
rect 34161 19397 34195 19431
rect 49433 19397 49467 19431
rect 7021 19329 7055 19363
rect 9505 19329 9539 19363
rect 12541 19329 12575 19363
rect 14657 19329 14691 19363
rect 21189 19329 21223 19363
rect 23745 19329 23779 19363
rect 34805 19329 34839 19363
rect 44097 19329 44131 19363
rect 44281 19329 44315 19363
rect 45477 19329 45511 19363
rect 4169 19261 4203 19295
rect 4629 19261 4663 19295
rect 6469 19261 6503 19295
rect 8309 19261 8343 19295
rect 8861 19261 8895 19295
rect 11253 19261 11287 19295
rect 12081 19261 12115 19295
rect 14473 19261 14507 19295
rect 15117 19261 15151 19295
rect 18153 19261 18187 19295
rect 19349 19261 19383 19295
rect 22017 19261 22051 19295
rect 23489 19261 23523 19295
rect 25237 19261 25271 19295
rect 27997 19261 28031 19295
rect 28825 19261 28859 19295
rect 31125 19261 31159 19295
rect 32781 19261 32815 19295
rect 33517 19261 33551 19295
rect 33609 19261 33643 19295
rect 37933 19261 37967 19295
rect 38669 19261 38703 19295
rect 39313 19261 39347 19295
rect 42257 19261 42291 19295
rect 43085 19261 43119 19295
rect 43244 19261 43278 19295
rect 43361 19261 43395 19295
rect 46029 19261 46063 19295
rect 47317 19261 47351 19295
rect 49249 19261 49283 19295
rect 53481 19261 53515 19295
rect 56425 19261 56459 19295
rect 15025 19193 15059 19227
rect 19717 19193 19751 19227
rect 22569 19193 22603 19227
rect 41521 19193 41555 19227
rect 43637 19193 43671 19227
rect 49893 19193 49927 19227
rect 3525 19125 3559 19159
rect 5273 19125 5307 19159
rect 8677 19125 8711 19159
rect 10701 19125 10735 19159
rect 11529 19125 11563 19159
rect 12909 19125 12943 19159
rect 13645 19125 13679 19159
rect 13921 19125 13955 19159
rect 21465 19125 21499 19159
rect 22937 19125 22971 19159
rect 27261 19125 27295 19159
rect 27445 19125 27479 19159
rect 28273 19125 28307 19159
rect 30573 19125 30607 19159
rect 31585 19125 31619 19159
rect 32137 19125 32171 19159
rect 33149 19125 33183 19159
rect 35081 19125 35115 19159
rect 36921 19125 36955 19159
rect 38025 19125 38059 19159
rect 41613 19125 41647 19159
rect 42441 19125 42475 19159
rect 44557 19125 44591 19159
rect 46857 19125 46891 19159
rect 47777 19125 47811 19159
rect 48237 19125 48271 19159
rect 48605 19125 48639 19159
rect 50169 19125 50203 19159
rect 52193 19125 52227 19159
rect 52929 19125 52963 19159
rect 4537 18921 4571 18955
rect 6469 18921 6503 18955
rect 8493 18921 8527 18955
rect 11161 18921 11195 18955
rect 27445 18921 27479 18955
rect 30757 18921 30791 18955
rect 40969 18921 41003 18955
rect 42625 18921 42659 18955
rect 45569 18921 45603 18955
rect 4813 18853 4847 18887
rect 9689 18853 9723 18887
rect 17601 18853 17635 18887
rect 21373 18853 21407 18887
rect 22201 18853 22235 18887
rect 24409 18853 24443 18887
rect 35449 18853 35483 18887
rect 37749 18853 37783 18887
rect 42533 18853 42567 18887
rect 52285 18853 52319 18887
rect 56149 18853 56183 18887
rect 3985 18785 4019 18819
rect 7021 18785 7055 18819
rect 9137 18785 9171 18819
rect 10057 18785 10091 18819
rect 11621 18785 11655 18819
rect 11805 18785 11839 18819
rect 13737 18785 13771 18819
rect 14197 18785 14231 18819
rect 17509 18785 17543 18819
rect 18245 18785 18279 18819
rect 19993 18785 20027 18819
rect 21557 18785 21591 18819
rect 22845 18785 22879 18819
rect 24225 18785 24259 18819
rect 25053 18785 25087 18819
rect 26525 18785 26559 18819
rect 27169 18785 27203 18819
rect 27997 18785 28031 18819
rect 31309 18785 31343 18819
rect 32229 18785 32263 18819
rect 33057 18785 33091 18819
rect 34897 18785 34931 18819
rect 36093 18785 36127 18819
rect 37105 18785 37139 18819
rect 37289 18785 37323 18819
rect 38393 18785 38427 18819
rect 41153 18785 41187 18819
rect 43177 18785 43211 18819
rect 44741 18785 44775 18819
rect 45477 18785 45511 18819
rect 46213 18785 46247 18819
rect 48421 18785 48455 18819
rect 48789 18785 48823 18819
rect 52193 18785 52227 18819
rect 52837 18785 52871 18819
rect 55137 18785 55171 18819
rect 55505 18785 55539 18819
rect 4169 18717 4203 18751
rect 5641 18717 5675 18751
rect 7849 18717 7883 18751
rect 9321 18717 9355 18751
rect 11069 18717 11103 18751
rect 11529 18717 11563 18751
rect 12541 18717 12575 18751
rect 14473 18717 14507 18751
rect 14933 18717 14967 18751
rect 17969 18717 18003 18751
rect 19073 18717 19107 18751
rect 19809 18717 19843 18751
rect 23489 18717 23523 18751
rect 25881 18717 25915 18751
rect 26985 18717 27019 18751
rect 27813 18717 27847 18751
rect 28825 18717 28859 18751
rect 30113 18717 30147 18751
rect 31125 18717 31159 18751
rect 32045 18717 32079 18751
rect 33241 18717 33275 18751
rect 34253 18717 34287 18751
rect 34989 18717 35023 18751
rect 36829 18717 36863 18751
rect 38577 18717 38611 18751
rect 43453 18717 43487 18751
rect 44005 18717 44039 18751
rect 45937 18717 45971 18751
rect 47041 18717 47075 18751
rect 47685 18717 47719 18751
rect 48237 18717 48271 18751
rect 49065 18717 49099 18751
rect 50353 18717 50387 18751
rect 53665 18717 53699 18751
rect 55781 18717 55815 18751
rect 56793 18717 56827 18751
rect 57529 18717 57563 18751
rect 4077 18649 4111 18683
rect 4997 18649 5031 18683
rect 6837 18649 6871 18683
rect 20260 18649 20294 18683
rect 27905 18649 27939 18683
rect 31217 18649 31251 18683
rect 33149 18649 33183 18683
rect 33701 18649 33735 18683
rect 35081 18649 35115 18683
rect 36277 18649 36311 18683
rect 41420 18649 41454 18683
rect 43085 18649 43119 18683
rect 44189 18649 44223 18683
rect 48329 18649 48363 18683
rect 52653 18649 52687 18683
rect 6377 18581 6411 18615
rect 6929 18581 6963 18615
rect 7297 18581 7331 18615
rect 9229 18581 9263 18615
rect 10425 18581 10459 18615
rect 11989 18581 12023 18615
rect 13001 18581 13035 18615
rect 13185 18581 13219 18615
rect 13553 18581 13587 18615
rect 13645 18581 13679 18615
rect 14381 18581 14415 18615
rect 14841 18581 14875 18615
rect 15577 18581 15611 18615
rect 18061 18581 18095 18615
rect 18429 18581 18463 18615
rect 19257 18581 19291 18615
rect 21741 18581 21775 18615
rect 21833 18581 21867 18615
rect 22293 18581 22327 18615
rect 23581 18581 23615 18615
rect 24777 18581 24811 18615
rect 24869 18581 24903 18615
rect 25237 18581 25271 18615
rect 26617 18581 26651 18615
rect 27077 18581 27111 18615
rect 28273 18581 28307 18615
rect 29561 18581 29595 18615
rect 30665 18581 30699 18615
rect 31585 18581 31619 18615
rect 31953 18581 31987 18615
rect 32689 18581 32723 18615
rect 33609 18581 33643 18615
rect 35541 18581 35575 18615
rect 37381 18581 37415 18615
rect 37841 18581 37875 18615
rect 39221 18581 39255 18615
rect 39589 18581 39623 18615
rect 42993 18581 43027 18615
rect 46029 18581 46063 18615
rect 46397 18581 46431 18615
rect 47133 18581 47167 18615
rect 47869 18581 47903 18615
rect 48973 18581 49007 18615
rect 49433 18581 49467 18615
rect 50997 18581 51031 18615
rect 51549 18581 51583 18615
rect 52745 18581 52779 18615
rect 53113 18581 53147 18615
rect 54125 18581 54159 18615
rect 55689 18581 55723 18615
rect 56241 18581 56275 18615
rect 56977 18581 57011 18615
rect 8217 18377 8251 18411
rect 11529 18377 11563 18411
rect 11897 18377 11931 18411
rect 11989 18377 12023 18411
rect 12633 18377 12667 18411
rect 18337 18377 18371 18411
rect 18797 18377 18831 18411
rect 19165 18377 19199 18411
rect 22661 18377 22695 18411
rect 24961 18377 24995 18411
rect 28549 18377 28583 18411
rect 28641 18377 28675 18411
rect 29101 18377 29135 18411
rect 32413 18377 32447 18411
rect 34437 18377 34471 18411
rect 38669 18377 38703 18411
rect 39037 18377 39071 18411
rect 43177 18377 43211 18411
rect 44741 18377 44775 18411
rect 46213 18377 46247 18411
rect 46673 18377 46707 18411
rect 47041 18377 47075 18411
rect 47593 18377 47627 18411
rect 52561 18377 52595 18411
rect 53113 18377 53147 18411
rect 53481 18377 53515 18411
rect 53941 18377 53975 18411
rect 57253 18377 57287 18411
rect 4712 18309 4746 18343
rect 10232 18309 10266 18343
rect 15770 18309 15804 18343
rect 17224 18309 17258 18343
rect 18705 18309 18739 18343
rect 23734 18309 23768 18343
rect 27436 18309 27470 18343
rect 29009 18309 29043 18343
rect 30380 18309 30414 18343
rect 37556 18309 37590 18343
rect 46581 18309 46615 18343
rect 50660 18309 50694 18343
rect 51448 18309 51482 18343
rect 53021 18309 53055 18343
rect 56140 18309 56174 18343
rect 2973 18241 3007 18275
rect 3240 18241 3274 18275
rect 4445 18241 4479 18275
rect 6377 18241 6411 18275
rect 9433 18241 9467 18275
rect 13277 18241 13311 18275
rect 16037 18241 16071 18275
rect 16957 18241 16991 18275
rect 20407 18241 20441 18275
rect 22201 18241 22235 18275
rect 23213 18241 23247 18275
rect 26617 18241 26651 18275
rect 30113 18241 30147 18275
rect 33149 18241 33183 18275
rect 34161 18241 34195 18275
rect 35550 18241 35584 18275
rect 35817 18241 35851 18275
rect 37013 18241 37047 18275
rect 37289 18241 37323 18275
rect 39129 18241 39163 18275
rect 40877 18241 40911 18275
rect 41144 18241 41178 18275
rect 42717 18241 42751 18275
rect 42809 18241 42843 18275
rect 43269 18241 43303 18275
rect 44833 18241 44867 18275
rect 45100 18241 45134 18275
rect 48375 18241 48409 18275
rect 54585 18241 54619 18275
rect 55597 18241 55631 18275
rect 55781 18241 55815 18275
rect 6561 18173 6595 18207
rect 7297 18173 7331 18207
rect 7414 18173 7448 18207
rect 7573 18173 7607 18207
rect 9689 18173 9723 18207
rect 9965 18173 9999 18207
rect 12173 18173 12207 18207
rect 13415 18173 13449 18207
rect 13553 18173 13587 18207
rect 14289 18173 14323 18207
rect 14473 18173 14507 18207
rect 18521 18173 18555 18207
rect 19533 18173 19567 18207
rect 20269 18173 20303 18207
rect 20545 18173 20579 18207
rect 21281 18173 21315 18207
rect 21465 18173 21499 18207
rect 22293 18173 22327 18207
rect 22385 18173 22419 18207
rect 23489 18173 23523 18207
rect 25605 18173 25639 18207
rect 25764 18173 25798 18207
rect 25881 18173 25915 18207
rect 26157 18173 26191 18207
rect 26801 18173 26835 18207
rect 27169 18173 27203 18207
rect 29193 18173 29227 18207
rect 33287 18173 33321 18207
rect 33425 18173 33459 18207
rect 34345 18173 34379 18207
rect 38945 18173 38979 18207
rect 40141 18173 40175 18207
rect 42533 18173 42567 18207
rect 43821 18173 43855 18207
rect 46489 18173 46523 18207
rect 48239 18173 48273 18207
rect 48513 18173 48547 18207
rect 48789 18173 48823 18207
rect 49249 18173 49283 18207
rect 49433 18173 49467 18207
rect 50905 18173 50939 18207
rect 51181 18173 51215 18207
rect 52837 18173 52871 18207
rect 54723 18173 54757 18207
rect 54861 18173 54895 18207
rect 55873 18173 55907 18207
rect 58449 18173 58483 18207
rect 5825 18105 5859 18139
rect 7021 18105 7055 18139
rect 8309 18105 8343 18139
rect 13829 18105 13863 18139
rect 19625 18105 19659 18139
rect 20821 18105 20855 18139
rect 24869 18105 24903 18139
rect 31493 18105 31527 18139
rect 33701 18105 33735 18139
rect 39497 18105 39531 18139
rect 42257 18105 42291 18139
rect 53757 18105 53791 18139
rect 55137 18105 55171 18139
rect 4353 18037 4387 18071
rect 11345 18037 11379 18071
rect 14657 18037 14691 18071
rect 21833 18037 21867 18071
rect 31861 18037 31895 18071
rect 32505 18037 32539 18071
rect 39589 18037 39623 18071
rect 47317 18037 47351 18071
rect 49525 18037 49559 18071
rect 57897 18037 57931 18071
rect 3801 17833 3835 17867
rect 5917 17833 5951 17867
rect 8677 17833 8711 17867
rect 9689 17833 9723 17867
rect 9781 17833 9815 17867
rect 14105 17833 14139 17867
rect 14841 17833 14875 17867
rect 18429 17833 18463 17867
rect 20177 17833 20211 17867
rect 24225 17833 24259 17867
rect 25789 17833 25823 17867
rect 28457 17833 28491 17867
rect 33701 17833 33735 17867
rect 44833 17833 44867 17867
rect 46489 17833 46523 17867
rect 48697 17833 48731 17867
rect 49893 17833 49927 17867
rect 53113 17833 53147 17867
rect 54125 17833 54159 17867
rect 56057 17833 56091 17867
rect 57713 17833 57747 17867
rect 13921 17765 13955 17799
rect 18337 17765 18371 17799
rect 37197 17765 37231 17799
rect 38117 17765 38151 17799
rect 42717 17765 42751 17799
rect 46397 17765 46431 17799
rect 53021 17765 53055 17799
rect 4353 17697 4387 17731
rect 5273 17697 5307 17731
rect 7297 17697 7331 17731
rect 9137 17697 9171 17731
rect 10517 17697 10551 17731
rect 12541 17697 12575 17731
rect 14657 17697 14691 17731
rect 15393 17697 15427 17731
rect 16221 17697 16255 17731
rect 16957 17697 16991 17731
rect 19073 17697 19107 17731
rect 24409 17697 24443 17731
rect 27077 17697 27111 17731
rect 30205 17697 30239 17731
rect 34437 17697 34471 17731
rect 34805 17697 34839 17731
rect 37473 17697 37507 17731
rect 38393 17697 38427 17731
rect 38669 17697 38703 17731
rect 47133 17697 47167 17731
rect 49249 17697 49283 17731
rect 50721 17697 50755 17731
rect 53757 17697 53791 17731
rect 55413 17697 55447 17731
rect 55597 17697 55631 17731
rect 3525 17629 3559 17663
rect 4261 17629 4295 17663
rect 7030 17629 7064 17663
rect 9321 17629 9355 17663
rect 10333 17629 10367 17663
rect 10773 17629 10807 17663
rect 12449 17629 12483 17663
rect 15301 17629 15335 17663
rect 19625 17629 19659 17663
rect 21649 17629 21683 17663
rect 22293 17629 22327 17663
rect 26433 17629 26467 17663
rect 27344 17629 27378 17663
rect 32321 17629 32355 17663
rect 34989 17629 35023 17663
rect 37657 17629 37691 17663
rect 38510 17629 38544 17663
rect 45017 17629 45051 17663
rect 45284 17629 45318 17663
rect 47317 17629 47351 17663
rect 51181 17629 51215 17663
rect 51641 17629 51675 17663
rect 56333 17629 56367 17663
rect 58357 17629 58391 17663
rect 4169 17561 4203 17595
rect 4629 17561 4663 17595
rect 5641 17561 5675 17595
rect 12808 17561 12842 17595
rect 15209 17561 15243 17595
rect 15669 17561 15703 17595
rect 17224 17561 17258 17595
rect 21404 17561 21438 17595
rect 24676 17561 24710 17595
rect 30472 17561 30506 17595
rect 31861 17561 31895 17595
rect 32588 17561 32622 17595
rect 35081 17561 35115 17595
rect 36737 17561 36771 17595
rect 47584 17561 47618 17595
rect 49525 17561 49559 17595
rect 50169 17561 50203 17595
rect 51908 17561 51942 17595
rect 56600 17561 56634 17595
rect 57805 17561 57839 17595
rect 2973 17493 3007 17527
rect 8309 17493 8343 17527
rect 9229 17493 9263 17527
rect 11897 17493 11931 17527
rect 20269 17493 20303 17527
rect 21741 17493 21775 17527
rect 23857 17493 23891 17527
rect 25881 17493 25915 17527
rect 28733 17493 28767 17527
rect 31585 17493 31619 17527
rect 33977 17493 34011 17527
rect 35449 17493 35483 17527
rect 39313 17493 39347 17527
rect 42349 17493 42383 17527
rect 43269 17493 43303 17527
rect 48973 17493 49007 17527
rect 49433 17493 49467 17527
rect 55045 17493 55079 17527
rect 55689 17493 55723 17527
rect 3341 17289 3375 17323
rect 6837 17289 6871 17323
rect 9229 17289 9263 17323
rect 13001 17289 13035 17323
rect 14749 17289 14783 17323
rect 17417 17289 17451 17323
rect 20545 17289 20579 17323
rect 21005 17289 21039 17323
rect 22109 17289 22143 17323
rect 25053 17289 25087 17323
rect 26065 17289 26099 17323
rect 31033 17289 31067 17323
rect 32137 17289 32171 17323
rect 32873 17289 32907 17323
rect 37841 17289 37875 17323
rect 39773 17289 39807 17323
rect 43729 17289 43763 17323
rect 47225 17289 47259 17323
rect 47777 17289 47811 17323
rect 48513 17289 48547 17323
rect 57069 17289 57103 17323
rect 57437 17289 57471 17323
rect 3709 17221 3743 17255
rect 9873 17221 9907 17255
rect 24593 17221 24627 17255
rect 38976 17221 39010 17255
rect 3801 17153 3835 17187
rect 4169 17153 4203 17187
rect 8125 17153 8159 17187
rect 13553 17153 13587 17187
rect 17969 17153 18003 17187
rect 20913 17153 20947 17187
rect 31585 17153 31619 17187
rect 32781 17153 32815 17187
rect 33517 17153 33551 17187
rect 39681 17153 39715 17187
rect 48421 17153 48455 17187
rect 49157 17153 49191 17187
rect 3249 17085 3283 17119
rect 3985 17085 4019 17119
rect 4721 17085 4755 17119
rect 6193 17085 6227 17119
rect 8769 17085 8803 17119
rect 21097 17085 21131 17119
rect 24317 17085 24351 17119
rect 24501 17085 24535 17119
rect 25605 17085 25639 17119
rect 39221 17085 39255 17119
rect 39865 17085 39899 17119
rect 42993 17085 43027 17119
rect 43453 17085 43487 17119
rect 43637 17085 43671 17119
rect 44281 17085 44315 17119
rect 45569 17085 45603 17119
rect 56609 17085 56643 17119
rect 56885 17085 56919 17119
rect 56977 17085 57011 17119
rect 58449 17085 58483 17119
rect 24961 17017 24995 17051
rect 44925 17017 44959 17051
rect 2605 16949 2639 16983
rect 5181 16949 5215 16983
rect 8217 16949 8251 16983
rect 12449 16949 12483 16983
rect 18337 16949 18371 16983
rect 19349 16949 19383 16983
rect 20361 16949 20395 16983
rect 24133 16949 24167 16983
rect 34345 16949 34379 16983
rect 35541 16949 35575 16983
rect 37013 16949 37047 16983
rect 37473 16949 37507 16983
rect 39313 16949 39347 16983
rect 41613 16949 41647 16983
rect 42441 16949 42475 16983
rect 44097 16949 44131 16983
rect 44833 16949 44867 16983
rect 53205 16949 53239 16983
rect 53573 16949 53607 16983
rect 55781 16949 55815 16983
rect 56149 16949 56183 16983
rect 57897 16949 57931 16983
rect 4537 16745 4571 16779
rect 6469 16745 6503 16779
rect 23489 16745 23523 16779
rect 31677 16745 31711 16779
rect 33793 16745 33827 16779
rect 39129 16745 39163 16779
rect 44557 16745 44591 16779
rect 51089 16745 51123 16779
rect 5733 16677 5767 16711
rect 13185 16677 13219 16711
rect 32045 16677 32079 16711
rect 41705 16677 41739 16711
rect 44281 16677 44315 16711
rect 57345 16677 57379 16711
rect 5340 16609 5374 16643
rect 6193 16609 6227 16643
rect 6377 16609 6411 16643
rect 8585 16609 8619 16643
rect 9505 16609 9539 16643
rect 17693 16609 17727 16643
rect 18797 16609 18831 16643
rect 23673 16609 23707 16643
rect 25605 16609 25639 16643
rect 36001 16609 36035 16643
rect 37841 16609 37875 16643
rect 42257 16609 42291 16643
rect 42349 16609 42383 16643
rect 42901 16609 42935 16643
rect 45569 16609 45603 16643
rect 56517 16609 56551 16643
rect 56793 16609 56827 16643
rect 57989 16609 58023 16643
rect 2237 16541 2271 16575
rect 2504 16541 2538 16575
rect 4353 16541 4387 16575
rect 5181 16541 5215 16575
rect 5457 16541 5491 16575
rect 7849 16541 7883 16575
rect 11529 16541 11563 16575
rect 12357 16541 12391 16575
rect 13829 16541 13863 16575
rect 14105 16541 14139 16575
rect 15393 16541 15427 16575
rect 18337 16541 18371 16575
rect 21373 16541 21407 16575
rect 25053 16541 25087 16575
rect 26341 16541 26375 16575
rect 30849 16541 30883 16575
rect 35265 16541 35299 16575
rect 37013 16541 37047 16575
rect 37933 16541 37967 16575
rect 40141 16541 40175 16575
rect 40325 16541 40359 16575
rect 43168 16541 43202 16575
rect 45385 16541 45419 16575
rect 47777 16541 47811 16575
rect 49157 16541 49191 16575
rect 50721 16541 50755 16575
rect 53849 16541 53883 16575
rect 56977 16541 57011 16575
rect 7604 16473 7638 16507
rect 34253 16473 34287 16507
rect 40592 16473 40626 16507
rect 3617 16405 3651 16439
rect 3801 16405 3835 16439
rect 7941 16405 7975 16439
rect 8309 16405 8343 16439
rect 8401 16405 8435 16439
rect 8953 16405 8987 16439
rect 10885 16405 10919 16439
rect 11713 16405 11747 16439
rect 12725 16405 12759 16439
rect 13277 16405 13311 16439
rect 14749 16405 14783 16439
rect 14841 16405 14875 16439
rect 17049 16405 17083 16439
rect 17785 16405 17819 16439
rect 20821 16405 20855 16439
rect 24225 16405 24259 16439
rect 24409 16405 24443 16439
rect 25789 16405 25823 16439
rect 30297 16405 30331 16439
rect 31217 16405 31251 16439
rect 34713 16405 34747 16439
rect 35449 16405 35483 16439
rect 36461 16405 36495 16439
rect 37197 16405 37231 16439
rect 38577 16405 38611 16439
rect 41797 16405 41831 16439
rect 42165 16405 42199 16439
rect 45017 16405 45051 16439
rect 45477 16405 45511 16439
rect 48421 16405 48455 16439
rect 48605 16405 48639 16439
rect 50169 16405 50203 16439
rect 53205 16405 53239 16439
rect 56885 16405 56919 16439
rect 57437 16405 57471 16439
rect 3525 16201 3559 16235
rect 3893 16201 3927 16235
rect 3985 16201 4019 16235
rect 6193 16201 6227 16235
rect 7297 16201 7331 16235
rect 8769 16201 8803 16235
rect 11529 16201 11563 16235
rect 11897 16201 11931 16235
rect 13185 16201 13219 16235
rect 13645 16201 13679 16235
rect 14105 16201 14139 16235
rect 19717 16201 19751 16235
rect 24041 16201 24075 16235
rect 24869 16201 24903 16235
rect 25881 16201 25915 16235
rect 30481 16201 30515 16235
rect 33977 16201 34011 16235
rect 37105 16201 37139 16235
rect 41245 16201 41279 16235
rect 42441 16201 42475 16235
rect 47593 16201 47627 16235
rect 48053 16201 48087 16235
rect 51733 16201 51767 16235
rect 53021 16201 53055 16235
rect 53297 16201 53331 16235
rect 55781 16201 55815 16235
rect 57713 16201 57747 16235
rect 2320 16133 2354 16167
rect 7634 16133 7668 16167
rect 16948 16133 16982 16167
rect 33885 16133 33919 16167
rect 35112 16133 35146 16167
rect 35992 16133 36026 16167
rect 38424 16133 38458 16167
rect 49516 16133 49550 16167
rect 56600 16133 56634 16167
rect 2053 16065 2087 16099
rect 7389 16065 7423 16099
rect 9413 16065 9447 16099
rect 11989 16065 12023 16099
rect 13277 16065 13311 16099
rect 14013 16065 14047 16099
rect 19349 16065 19383 16099
rect 20933 16065 20967 16099
rect 21189 16065 21223 16099
rect 23949 16065 23983 16099
rect 26249 16065 26283 16099
rect 26341 16065 26375 16099
rect 26985 16065 27019 16099
rect 30849 16065 30883 16099
rect 30941 16065 30975 16099
rect 31309 16065 31343 16099
rect 35357 16065 35391 16099
rect 35725 16065 35759 16099
rect 38669 16065 38703 16099
rect 41797 16065 41831 16099
rect 43361 16065 43395 16099
rect 44097 16065 44131 16099
rect 47961 16065 47995 16099
rect 49249 16065 49283 16099
rect 53665 16065 53699 16099
rect 54861 16065 54895 16099
rect 58449 16065 58483 16099
rect 4169 15997 4203 16031
rect 6745 15997 6779 16031
rect 11345 15997 11379 16031
rect 12173 15997 12207 16031
rect 13001 15997 13035 16031
rect 13921 15997 13955 16031
rect 14933 15997 14967 16031
rect 16681 15997 16715 16031
rect 18981 15997 19015 16031
rect 22937 15997 22971 16031
rect 24133 15997 24167 16031
rect 25513 15997 25547 16031
rect 26525 15997 26559 16031
rect 27537 15997 27571 16031
rect 28365 15997 28399 16031
rect 30389 15997 30423 16031
rect 31033 15997 31067 16031
rect 31861 15997 31895 16031
rect 39313 15997 39347 16031
rect 43085 15997 43119 16031
rect 43244 15997 43278 16031
rect 43637 15997 43671 16031
rect 44281 15997 44315 16031
rect 44925 15997 44959 16031
rect 48145 15997 48179 16031
rect 49065 15997 49099 16031
rect 51273 15997 51307 16031
rect 53757 15997 53791 16031
rect 53849 15997 53883 16031
rect 54677 15997 54711 16031
rect 55413 15997 55447 16031
rect 56333 15997 56367 16031
rect 3433 15929 3467 15963
rect 12817 15929 12851 15963
rect 14473 15929 14507 15963
rect 18061 15929 18095 15963
rect 23581 15929 23615 15963
rect 42165 15929 42199 15963
rect 47317 15929 47351 15963
rect 4629 15861 4663 15895
rect 8861 15861 8895 15895
rect 10701 15861 10735 15895
rect 15577 15861 15611 15895
rect 18337 15861 18371 15895
rect 19809 15861 19843 15895
rect 21557 15861 21591 15895
rect 23489 15861 23523 15895
rect 24961 15861 24995 15895
rect 27813 15861 27847 15895
rect 32597 15861 32631 15895
rect 37289 15861 37323 15895
rect 38761 15861 38795 15895
rect 41061 15861 41095 15895
rect 44373 15861 44407 15895
rect 45293 15861 45327 15895
rect 47041 15861 47075 15895
rect 48421 15861 48455 15895
rect 50629 15861 50663 15895
rect 50721 15861 50755 15895
rect 52561 15861 52595 15895
rect 54125 15861 54159 15895
rect 56149 15861 56183 15895
rect 57897 15861 57931 15895
rect 7757 15657 7791 15691
rect 9229 15657 9263 15691
rect 11529 15657 11563 15691
rect 14105 15657 14139 15691
rect 18061 15657 18095 15691
rect 21189 15657 21223 15691
rect 22753 15657 22787 15691
rect 25145 15657 25179 15691
rect 27629 15657 27663 15691
rect 36829 15657 36863 15691
rect 37657 15657 37691 15691
rect 40141 15657 40175 15691
rect 49065 15657 49099 15691
rect 49985 15657 50019 15691
rect 54217 15657 54251 15691
rect 54309 15657 54343 15691
rect 20453 15589 20487 15623
rect 26893 15589 26927 15623
rect 31217 15589 31251 15623
rect 33517 15589 33551 15623
rect 35449 15589 35483 15623
rect 41705 15589 41739 15623
rect 44097 15589 44131 15623
rect 8401 15521 8435 15555
rect 12863 15521 12897 15555
rect 13001 15521 13035 15555
rect 13277 15521 13311 15555
rect 13737 15521 13771 15555
rect 13921 15521 13955 15555
rect 18521 15521 18555 15555
rect 18705 15521 18739 15555
rect 20039 15521 20073 15555
rect 20177 15521 20211 15555
rect 21833 15521 21867 15555
rect 24593 15521 24627 15555
rect 24685 15521 24719 15555
rect 25513 15521 25547 15555
rect 26341 15521 26375 15555
rect 26500 15521 26534 15555
rect 27353 15521 27387 15555
rect 31401 15521 31435 15555
rect 32965 15521 32999 15555
rect 33241 15521 33275 15555
rect 33977 15521 34011 15555
rect 34897 15521 34931 15555
rect 36093 15521 36127 15555
rect 37381 15521 37415 15555
rect 38209 15521 38243 15555
rect 40325 15521 40359 15555
rect 42349 15521 42383 15555
rect 43177 15521 43211 15555
rect 43545 15521 43579 15555
rect 43637 15521 43671 15555
rect 44741 15521 44775 15555
rect 49433 15521 49467 15555
rect 50353 15521 50387 15555
rect 54861 15521 54895 15555
rect 56103 15521 56137 15555
rect 56517 15521 56551 15555
rect 57161 15521 57195 15555
rect 57437 15521 57471 15555
rect 57529 15521 57563 15555
rect 3249 15453 3283 15487
rect 4353 15453 4387 15487
rect 5917 15453 5951 15487
rect 6653 15453 6687 15487
rect 8125 15453 8159 15487
rect 10149 15453 10183 15487
rect 10416 15453 10450 15487
rect 12725 15453 12759 15487
rect 15229 15453 15263 15487
rect 15485 15453 15519 15487
rect 16589 15453 16623 15487
rect 16856 15453 16890 15487
rect 19901 15453 19935 15487
rect 20913 15453 20947 15487
rect 21097 15453 21131 15487
rect 22569 15453 22603 15487
rect 23866 15453 23900 15487
rect 24133 15453 24167 15487
rect 26617 15453 26651 15487
rect 27537 15453 27571 15487
rect 29009 15453 29043 15487
rect 29837 15453 29871 15487
rect 33124 15453 33158 15487
rect 34161 15453 34195 15487
rect 36461 15453 36495 15487
rect 37197 15453 37231 15487
rect 38025 15453 38059 15487
rect 42257 15453 42291 15487
rect 43729 15453 43763 15487
rect 46213 15453 46247 15487
rect 47685 15453 47719 15487
rect 47952 15453 47986 15487
rect 50629 15453 50663 15487
rect 52377 15453 52411 15487
rect 52745 15453 52779 15487
rect 52837 15453 52871 15487
rect 54677 15453 54711 15487
rect 55965 15453 55999 15487
rect 56241 15453 56275 15487
rect 56977 15453 57011 15487
rect 7021 15385 7055 15419
rect 24777 15385 24811 15419
rect 28764 15385 28798 15419
rect 30104 15385 30138 15419
rect 40592 15385 40626 15419
rect 42165 15385 42199 15419
rect 42625 15385 42659 15419
rect 46480 15385 46514 15419
rect 49525 15385 49559 15419
rect 53104 15385 53138 15419
rect 58265 15385 58299 15419
rect 2697 15317 2731 15351
rect 3801 15317 3835 15351
rect 5273 15317 5307 15351
rect 6101 15317 6135 15351
rect 8217 15317 8251 15351
rect 11989 15317 12023 15351
rect 12081 15317 12115 15351
rect 15761 15317 15795 15351
rect 16405 15317 16439 15351
rect 17969 15317 18003 15351
rect 18429 15317 18463 15351
rect 19257 15317 19291 15351
rect 21557 15317 21591 15351
rect 21649 15317 21683 15351
rect 22017 15317 22051 15351
rect 25697 15317 25731 15351
rect 29377 15317 29411 15351
rect 31585 15317 31619 15351
rect 31677 15317 31711 15351
rect 32045 15317 32079 15351
rect 32321 15317 32355 15351
rect 34529 15317 34563 15351
rect 34989 15317 35023 15351
rect 35081 15317 35115 15351
rect 35541 15317 35575 15351
rect 37289 15317 37323 15351
rect 38117 15317 38151 15351
rect 41797 15317 41831 15351
rect 44189 15317 44223 15351
rect 47593 15317 47627 15351
rect 49617 15317 49651 15351
rect 54769 15317 54803 15351
rect 55321 15317 55355 15351
rect 57621 15317 57655 15351
rect 57989 15317 58023 15351
rect 2973 15113 3007 15147
rect 3341 15113 3375 15147
rect 5733 15113 5767 15147
rect 6193 15113 6227 15147
rect 6745 15113 6779 15147
rect 7481 15113 7515 15147
rect 11529 15113 11563 15147
rect 11897 15113 11931 15147
rect 13185 15113 13219 15147
rect 17877 15113 17911 15147
rect 19165 15113 19199 15147
rect 21465 15113 21499 15147
rect 23489 15113 23523 15147
rect 24961 15113 24995 15147
rect 26709 15113 26743 15147
rect 27905 15113 27939 15147
rect 29193 15113 29227 15147
rect 31309 15113 31343 15147
rect 32137 15113 32171 15147
rect 34805 15113 34839 15147
rect 35265 15113 35299 15147
rect 37841 15113 37875 15147
rect 41245 15113 41279 15147
rect 42901 15113 42935 15147
rect 44741 15113 44775 15147
rect 46765 15113 46799 15147
rect 47961 15113 47995 15147
rect 54585 15113 54619 15147
rect 57529 15113 57563 15147
rect 3433 15045 3467 15079
rect 10232 15045 10266 15079
rect 14320 15045 14354 15079
rect 17049 15045 17083 15079
rect 20352 15045 20386 15079
rect 21833 15045 21867 15079
rect 23848 15045 23882 15079
rect 30104 15045 30138 15079
rect 33232 15045 33266 15079
rect 48697 15045 48731 15079
rect 52469 15045 52503 15079
rect 5825 14977 5859 15011
rect 11989 14977 12023 15011
rect 12357 14977 12391 15011
rect 13001 14977 13035 15011
rect 17509 14977 17543 15011
rect 17969 14977 18003 15011
rect 18613 14977 18647 15011
rect 20085 14977 20119 15011
rect 25329 14977 25363 15011
rect 25596 14977 25630 15011
rect 27813 14977 27847 15011
rect 31953 14977 31987 15011
rect 37473 14977 37507 15011
rect 41797 14977 41831 15011
rect 44117 14977 44151 15011
rect 44373 14977 44407 15011
rect 49433 14977 49467 15011
rect 49571 14977 49605 15011
rect 49709 14977 49743 15011
rect 50629 14977 50663 15011
rect 51845 14977 51879 15011
rect 52101 14977 52135 15011
rect 52929 14977 52963 15011
rect 53196 14977 53230 15011
rect 55229 14977 55263 15011
rect 56416 14977 56450 15011
rect 57897 14977 57931 15011
rect 58449 14977 58483 15011
rect 2881 14909 2915 14943
rect 3617 14909 3651 14943
rect 4353 14909 4387 14943
rect 5641 14909 5675 14943
rect 6469 14909 6503 14943
rect 6653 14909 6687 14943
rect 8585 14909 8619 14943
rect 9965 14909 9999 14943
rect 12081 14909 12115 14943
rect 14565 14909 14599 14943
rect 17233 14909 17267 14943
rect 17417 14909 17451 14943
rect 19441 14909 19475 14943
rect 22385 14909 22419 14943
rect 23581 14909 23615 14943
rect 27629 14909 27663 14943
rect 28549 14909 28583 14943
rect 29837 14909 29871 14943
rect 32689 14909 32723 14943
rect 32965 14909 32999 14943
rect 34621 14909 34655 14943
rect 34713 14909 34747 14943
rect 35817 14909 35851 14943
rect 38669 14909 38703 14943
rect 47409 14909 47443 14943
rect 48053 14909 48087 14943
rect 48145 14909 48179 14943
rect 49985 14909 50019 14943
rect 50445 14909 50479 14943
rect 56149 14909 56183 14943
rect 11345 14841 11379 14875
rect 16497 14841 16531 14875
rect 28273 14841 28307 14875
rect 31217 14841 31251 14875
rect 35173 14841 35207 14875
rect 39773 14841 39807 14875
rect 47593 14841 47627 14875
rect 50721 14841 50755 14875
rect 54309 14841 54343 14875
rect 2237 14773 2271 14807
rect 3801 14773 3835 14807
rect 7113 14773 7147 14807
rect 8033 14773 8067 14807
rect 14933 14773 14967 14807
rect 19993 14773 20027 14807
rect 27353 14773 27387 14807
rect 34345 14773 34379 14807
rect 36645 14773 36679 14807
rect 39313 14773 39347 14807
rect 42165 14773 42199 14807
rect 42993 14773 43027 14807
rect 46581 14773 46615 14807
rect 48789 14773 48823 14807
rect 55505 14773 55539 14807
rect 56057 14773 56091 14807
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 7021 14569 7055 14603
rect 11805 14569 11839 14603
rect 13921 14569 13955 14603
rect 21005 14569 21039 14603
rect 31401 14569 31435 14603
rect 38209 14569 38243 14603
rect 52285 14569 52319 14603
rect 54217 14569 54251 14603
rect 3525 14501 3559 14535
rect 5641 14501 5675 14535
rect 31953 14501 31987 14535
rect 48513 14501 48547 14535
rect 50537 14501 50571 14535
rect 51457 14501 51491 14535
rect 57253 14501 57287 14535
rect 5227 14433 5261 14467
rect 5365 14433 5399 14467
rect 6285 14433 6319 14467
rect 8585 14433 8619 14467
rect 12357 14433 12391 14467
rect 20453 14433 20487 14467
rect 39589 14433 39623 14467
rect 50813 14433 50847 14467
rect 52101 14433 52135 14467
rect 52837 14433 52871 14467
rect 56609 14433 56643 14467
rect 57897 14433 57931 14467
rect 2145 14365 2179 14399
rect 2412 14365 2446 14399
rect 5089 14365 5123 14399
rect 6101 14365 6135 14399
rect 8318 14365 8352 14399
rect 9505 14365 9539 14399
rect 10609 14365 10643 14399
rect 14197 14365 14231 14399
rect 17509 14365 17543 14399
rect 18337 14365 18371 14399
rect 20177 14365 20211 14399
rect 20637 14365 20671 14399
rect 21649 14365 21683 14399
rect 25421 14365 25455 14399
rect 26249 14365 26283 14399
rect 30849 14365 30883 14399
rect 34345 14365 34379 14399
rect 35265 14365 35299 14399
rect 38117 14365 38151 14399
rect 40417 14365 40451 14399
rect 43085 14365 43119 14399
rect 44097 14365 44131 14399
rect 49157 14365 49191 14399
rect 53665 14365 53699 14399
rect 16865 14297 16899 14331
rect 24685 14297 24719 14331
rect 37105 14297 37139 14331
rect 39344 14297 39378 14331
rect 39865 14297 39899 14331
rect 48605 14297 48639 14331
rect 49617 14297 49651 14331
rect 51089 14297 51123 14331
rect 51549 14297 51583 14331
rect 56333 14297 56367 14331
rect 56885 14297 56919 14331
rect 6561 14229 6595 14263
rect 7205 14229 7239 14263
rect 8953 14229 8987 14263
rect 10057 14229 10091 14263
rect 14841 14229 14875 14263
rect 16957 14229 16991 14263
rect 17785 14229 17819 14263
rect 20545 14229 20579 14263
rect 21097 14229 21131 14263
rect 24869 14229 24903 14263
rect 25605 14229 25639 14263
rect 26893 14229 26927 14263
rect 30297 14229 30331 14263
rect 32229 14229 32263 14263
rect 32873 14229 32907 14263
rect 33149 14229 33183 14263
rect 33793 14229 33827 14263
rect 34713 14229 34747 14263
rect 37473 14229 37507 14263
rect 42533 14229 42567 14263
rect 43453 14229 43487 14263
rect 44557 14229 44591 14263
rect 47409 14229 47443 14263
rect 50997 14229 51031 14263
rect 53113 14229 53147 14263
rect 56793 14229 56827 14263
rect 57345 14229 57379 14263
rect 3617 14025 3651 14059
rect 4077 14025 4111 14059
rect 4721 14025 4755 14059
rect 6193 14025 6227 14059
rect 8033 14025 8067 14059
rect 10241 14025 10275 14059
rect 12541 14025 12575 14059
rect 13001 14025 13035 14059
rect 16957 14025 16991 14059
rect 17325 14025 17359 14059
rect 20085 14025 20119 14059
rect 20269 14025 20303 14059
rect 25329 14025 25363 14059
rect 25421 14025 25455 14059
rect 25881 14025 25915 14059
rect 27721 14025 27755 14059
rect 28089 14025 28123 14059
rect 30021 14025 30055 14059
rect 30481 14025 30515 14059
rect 30941 14025 30975 14059
rect 34437 14025 34471 14059
rect 37657 14025 37691 14059
rect 39037 14025 39071 14059
rect 39497 14025 39531 14059
rect 47961 14025 47995 14059
rect 48329 14025 48363 14059
rect 49433 14025 49467 14059
rect 53021 14025 53055 14059
rect 53205 14025 53239 14059
rect 57897 14025 57931 14059
rect 5080 13957 5114 13991
rect 8769 13957 8803 13991
rect 14136 13957 14170 13991
rect 14565 13957 14599 13991
rect 24216 13957 24250 13991
rect 34805 13957 34839 13991
rect 56600 13957 56634 13991
rect 2145 13889 2179 13923
rect 2401 13889 2435 13923
rect 3985 13889 4019 13923
rect 4813 13889 4847 13923
rect 7941 13889 7975 13923
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 11529 13889 11563 13923
rect 15485 13889 15519 13923
rect 17417 13889 17451 13923
rect 21393 13889 21427 13923
rect 21833 13889 21867 13923
rect 23949 13889 23983 13923
rect 25789 13889 25823 13923
rect 30849 13889 30883 13923
rect 31309 13889 31343 13923
rect 33232 13889 33266 13923
rect 35817 13889 35851 13923
rect 37749 13889 37783 13923
rect 39129 13889 39163 13923
rect 40509 13889 40543 13923
rect 43260 13889 43294 13923
rect 44465 13889 44499 13923
rect 48973 13889 49007 13923
rect 50557 13889 50591 13923
rect 50813 13889 50847 13923
rect 52193 13889 52227 13923
rect 53573 13889 53607 13923
rect 54033 13889 54067 13923
rect 4261 13821 4295 13855
rect 7849 13821 7883 13855
rect 10149 13821 10183 13855
rect 10885 13821 10919 13855
rect 12081 13821 12115 13855
rect 14381 13821 14415 13855
rect 15209 13821 15243 13855
rect 16497 13821 16531 13855
rect 17601 13821 17635 13855
rect 18613 13821 18647 13855
rect 19349 13821 19383 13855
rect 21649 13821 21683 13855
rect 22385 13821 22419 13855
rect 25973 13821 26007 13855
rect 27169 13821 27203 13855
rect 27445 13821 27479 13855
rect 27629 13821 27663 13855
rect 28733 13821 28767 13855
rect 31125 13821 31159 13855
rect 31861 13821 31895 13855
rect 32689 13821 32723 13855
rect 32965 13821 32999 13855
rect 34897 13821 34931 13855
rect 35035 13821 35069 13855
rect 37105 13821 37139 13855
rect 37841 13821 37875 13855
rect 38853 13821 38887 13855
rect 39589 13821 39623 13855
rect 42993 13821 43027 13855
rect 45017 13821 45051 13855
rect 47409 13821 47443 13855
rect 47777 13821 47811 13855
rect 47869 13821 47903 13855
rect 50905 13821 50939 13855
rect 51457 13821 51491 13855
rect 53665 13821 53699 13855
rect 53757 13821 53791 13855
rect 54677 13821 54711 13855
rect 55321 13821 55355 13855
rect 56333 13821 56367 13855
rect 58449 13821 58483 13855
rect 3525 13753 3559 13787
rect 8401 13753 8435 13787
rect 26525 13753 26559 13787
rect 34345 13753 34379 13787
rect 37289 13753 37323 13787
rect 38393 13753 38427 13787
rect 57713 13753 57747 13787
rect 11345 13685 11379 13719
rect 17969 13685 18003 13719
rect 18705 13685 18739 13719
rect 28181 13685 28215 13719
rect 29285 13685 29319 13719
rect 30389 13685 30423 13719
rect 32137 13685 32171 13719
rect 35265 13685 35299 13719
rect 36461 13685 36495 13719
rect 40233 13685 40267 13719
rect 42257 13685 42291 13719
rect 44373 13685 44407 13719
rect 46765 13685 46799 13719
rect 48421 13685 48455 13719
rect 51641 13685 51675 13719
rect 54769 13685 54803 13719
rect 56149 13685 56183 13719
rect 14933 13481 14967 13515
rect 16129 13481 16163 13515
rect 17693 13481 17727 13515
rect 19073 13481 19107 13515
rect 21465 13481 21499 13515
rect 25513 13481 25547 13515
rect 27813 13481 27847 13515
rect 31217 13481 31251 13515
rect 34713 13481 34747 13515
rect 37473 13481 37507 13515
rect 43361 13481 43395 13515
rect 44281 13481 44315 13515
rect 49249 13481 49283 13515
rect 50905 13481 50939 13515
rect 10885 13413 10919 13447
rect 18521 13413 18555 13447
rect 24409 13413 24443 13447
rect 27077 13413 27111 13447
rect 33425 13413 33459 13447
rect 34345 13413 34379 13447
rect 35817 13413 35851 13447
rect 51733 13413 51767 13447
rect 54125 13413 54159 13447
rect 58265 13413 58299 13447
rect 11621 13345 11655 13379
rect 12679 13345 12713 13379
rect 12817 13345 12851 13379
rect 13093 13345 13127 13379
rect 13553 13345 13587 13379
rect 14197 13345 14231 13379
rect 15393 13345 15427 13379
rect 15577 13345 15611 13379
rect 16313 13345 16347 13379
rect 17877 13345 17911 13379
rect 18061 13345 18095 13379
rect 19533 13345 19567 13379
rect 20269 13345 20303 13379
rect 20913 13345 20947 13379
rect 24225 13345 24259 13379
rect 24961 13345 24995 13379
rect 25881 13345 25915 13379
rect 27721 13345 27755 13379
rect 31401 13345 31435 13379
rect 31585 13345 31619 13379
rect 32873 13345 32907 13379
rect 33011 13345 33045 13379
rect 33149 13345 33183 13379
rect 33885 13345 33919 13379
rect 35357 13345 35391 13379
rect 38025 13345 38059 13379
rect 38485 13345 38519 13379
rect 40049 13345 40083 13379
rect 42809 13345 42843 13379
rect 42993 13345 43027 13379
rect 43637 13345 43671 13379
rect 43821 13345 43855 13379
rect 46397 13345 46431 13379
rect 50353 13345 50387 13379
rect 51089 13345 51123 13379
rect 54309 13345 54343 13379
rect 54493 13345 54527 13379
rect 56103 13345 56137 13379
rect 56241 13345 56275 13379
rect 56517 13345 56551 13379
rect 56977 13345 57011 13379
rect 57805 13345 57839 13379
rect 6469 13277 6503 13311
rect 9505 13277 9539 13311
rect 11437 13277 11471 13311
rect 12541 13277 12575 13311
rect 13737 13277 13771 13311
rect 14381 13277 14415 13311
rect 15301 13277 15335 13311
rect 16580 13277 16614 13311
rect 19993 13277 20027 13311
rect 21005 13277 21039 13311
rect 21097 13277 21131 13311
rect 24869 13277 24903 13311
rect 26525 13277 26559 13311
rect 26663 13277 26697 13311
rect 26801 13277 26835 13311
rect 27537 13277 27571 13311
rect 29193 13277 29227 13311
rect 29837 13277 29871 13311
rect 31677 13277 31711 13311
rect 34069 13277 34103 13311
rect 36093 13277 36127 13311
rect 37841 13277 37875 13311
rect 38761 13277 38795 13311
rect 38878 13277 38912 13311
rect 39037 13277 39071 13311
rect 40233 13277 40267 13311
rect 40877 13277 40911 13311
rect 45753 13277 45787 13311
rect 47869 13277 47903 13311
rect 49893 13277 49927 13311
rect 50445 13277 50479 13311
rect 52101 13277 52135 13311
rect 52745 13277 52779 13311
rect 53012 13277 53046 13311
rect 55965 13277 55999 13311
rect 57161 13277 57195 13311
rect 57621 13277 57655 13311
rect 9772 13209 9806 13243
rect 20085 13209 20119 13243
rect 23489 13209 23523 13243
rect 28948 13209 28982 13243
rect 30104 13209 30138 13243
rect 36360 13209 36394 13243
rect 41144 13209 41178 13243
rect 46664 13209 46698 13243
rect 48136 13209 48170 13243
rect 51365 13209 51399 13243
rect 54585 13209 54619 13243
rect 57713 13209 57747 13243
rect 7113 13141 7147 13175
rect 10977 13141 11011 13175
rect 11345 13141 11379 13175
rect 11897 13141 11931 13175
rect 14473 13141 14507 13175
rect 14841 13141 14875 13175
rect 18153 13141 18187 13175
rect 19625 13141 19659 13175
rect 23581 13141 23615 13175
rect 24777 13141 24811 13175
rect 32045 13141 32079 13175
rect 32229 13141 32263 13175
rect 35081 13141 35115 13175
rect 35173 13141 35207 13175
rect 39681 13141 39715 13175
rect 40141 13141 40175 13175
rect 40601 13141 40635 13175
rect 42257 13141 42291 13175
rect 42349 13141 42383 13175
rect 42717 13141 42751 13175
rect 43913 13141 43947 13175
rect 44833 13141 44867 13175
rect 45201 13141 45235 13175
rect 47777 13141 47811 13175
rect 49341 13141 49375 13175
rect 50537 13141 50571 13175
rect 51273 13141 51307 13175
rect 52469 13141 52503 13175
rect 54953 13141 54987 13175
rect 55321 13141 55355 13175
rect 57253 13141 57287 13175
rect 6377 12937 6411 12971
rect 10977 12937 11011 12971
rect 12817 12937 12851 12971
rect 18061 12937 18095 12971
rect 24869 12937 24903 12971
rect 26341 12937 26375 12971
rect 26801 12937 26835 12971
rect 27813 12937 27847 12971
rect 29285 12937 29319 12971
rect 32321 12937 32355 12971
rect 34253 12937 34287 12971
rect 34621 12937 34655 12971
rect 37105 12937 37139 12971
rect 38761 12937 38795 12971
rect 41613 12937 41647 12971
rect 45017 12937 45051 12971
rect 47593 12937 47627 12971
rect 47961 12937 47995 12971
rect 48605 12937 48639 12971
rect 50997 12937 51031 12971
rect 52469 12937 52503 12971
rect 57529 12937 57563 12971
rect 8125 12869 8159 12903
rect 12449 12869 12483 12903
rect 16948 12869 16982 12903
rect 20269 12869 20303 12903
rect 30104 12869 30138 12903
rect 31309 12869 31343 12903
rect 33916 12869 33950 12903
rect 35992 12869 36026 12903
rect 37657 12869 37691 12903
rect 39896 12869 39930 12903
rect 40233 12869 40267 12903
rect 46152 12869 46186 12903
rect 46489 12869 46523 12903
rect 48053 12869 48087 12903
rect 1593 12801 1627 12835
rect 1860 12801 1894 12835
rect 5089 12801 5123 12835
rect 5273 12801 5307 12835
rect 6193 12801 6227 12835
rect 7490 12801 7524 12835
rect 7757 12801 7791 12835
rect 9597 12801 9631 12835
rect 9864 12801 9898 12835
rect 11529 12801 11563 12835
rect 12081 12801 12115 12835
rect 14217 12801 14251 12835
rect 14473 12801 14507 12835
rect 15117 12801 15151 12835
rect 16681 12801 16715 12835
rect 18337 12801 18371 12835
rect 19119 12801 19153 12835
rect 19257 12801 19291 12835
rect 19993 12801 20027 12835
rect 23653 12801 23687 12835
rect 25513 12801 25547 12835
rect 26433 12801 26467 12835
rect 27905 12801 27939 12835
rect 29837 12801 29871 12835
rect 31953 12801 31987 12835
rect 35725 12801 35759 12835
rect 42257 12801 42291 12835
rect 43888 12801 43922 12835
rect 44005 12801 44039 12835
rect 44741 12801 44775 12835
rect 46397 12801 46431 12835
rect 49433 12801 49467 12835
rect 49571 12801 49605 12835
rect 49709 12801 49743 12835
rect 50629 12801 50663 12835
rect 51089 12801 51123 12835
rect 51549 12801 51583 12835
rect 53104 12801 53138 12835
rect 54309 12801 54343 12835
rect 54953 12801 54987 12835
rect 55689 12801 55723 12835
rect 56057 12801 56091 12835
rect 56149 12801 56183 12835
rect 56416 12801 56450 12835
rect 58449 12801 58483 12835
rect 3065 12733 3099 12767
rect 5549 12733 5583 12767
rect 14565 12733 14599 12767
rect 18981 12733 19015 12767
rect 19533 12733 19567 12767
rect 20177 12733 20211 12767
rect 20821 12733 20855 12767
rect 23397 12733 23431 12767
rect 25881 12733 25915 12767
rect 26157 12733 26191 12767
rect 27629 12733 27663 12767
rect 28641 12733 28675 12767
rect 34161 12733 34195 12767
rect 34713 12733 34747 12767
rect 34897 12733 34931 12767
rect 35357 12733 35391 12767
rect 37749 12733 37783 12767
rect 37933 12733 37967 12767
rect 40141 12733 40175 12767
rect 40785 12733 40819 12767
rect 42625 12733 42659 12767
rect 43729 12733 43763 12767
rect 44925 12733 44959 12767
rect 47041 12733 47075 12767
rect 48145 12733 48179 12767
rect 48789 12733 48823 12767
rect 49985 12733 50019 12767
rect 50445 12733 50479 12767
rect 50905 12733 50939 12767
rect 52101 12733 52135 12767
rect 52837 12733 52871 12767
rect 2973 12665 3007 12699
rect 15577 12665 15611 12699
rect 24777 12665 24811 12699
rect 28273 12665 28307 12699
rect 31217 12665 31251 12699
rect 44281 12665 44315 12699
rect 54217 12665 54251 12699
rect 3709 12597 3743 12631
rect 5181 12597 5215 12631
rect 11253 12597 11287 12631
rect 13093 12597 13127 12631
rect 16129 12597 16163 12631
rect 16405 12597 16439 12631
rect 21189 12597 21223 12631
rect 23213 12597 23247 12631
rect 27445 12597 27479 12631
rect 32781 12597 32815 12631
rect 37289 12597 37323 12631
rect 38301 12597 38335 12631
rect 43085 12597 43119 12631
rect 51457 12597 51491 12631
rect 55229 12597 55263 12631
rect 57897 12597 57931 12631
rect 2237 12393 2271 12427
rect 5457 12393 5491 12427
rect 10425 12393 10459 12427
rect 15025 12393 15059 12427
rect 19993 12393 20027 12427
rect 27721 12393 27755 12427
rect 31677 12393 31711 12427
rect 34345 12393 34379 12427
rect 35357 12393 35391 12427
rect 36829 12393 36863 12427
rect 37657 12393 37691 12427
rect 38577 12393 38611 12427
rect 46857 12393 46891 12427
rect 48513 12393 48547 12427
rect 49341 12393 49375 12427
rect 52561 12393 52595 12427
rect 52929 12393 52963 12427
rect 54125 12393 54159 12427
rect 57253 12393 57287 12427
rect 12909 12325 12943 12359
rect 14749 12325 14783 12359
rect 27629 12325 27663 12359
rect 42625 12325 42659 12359
rect 45753 12325 45787 12359
rect 50169 12325 50203 12359
rect 57161 12325 57195 12359
rect 11069 12257 11103 12291
rect 13369 12257 13403 12291
rect 13461 12257 13495 12291
rect 14105 12257 14139 12291
rect 19349 12257 19383 12291
rect 21649 12257 21683 12291
rect 22385 12257 22419 12291
rect 28273 12257 28307 12291
rect 34713 12257 34747 12291
rect 37473 12257 37507 12291
rect 38301 12257 38335 12291
rect 43269 12257 43303 12291
rect 44189 12257 44223 12291
rect 45109 12257 45143 12291
rect 46121 12257 46155 12291
rect 51549 12257 51583 12291
rect 52193 12257 52227 12291
rect 56517 12257 56551 12291
rect 57805 12257 57839 12291
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 4353 12189 4387 12223
rect 4609 12189 4643 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5089 12189 5123 12223
rect 5273 12189 5307 12223
rect 5733 12189 5767 12223
rect 6377 12189 6411 12223
rect 8033 12189 8067 12223
rect 10149 12189 10183 12223
rect 11161 12189 11195 12223
rect 11713 12189 11747 12223
rect 13277 12189 13311 12223
rect 16497 12189 16531 12223
rect 19533 12189 19567 12223
rect 20085 12189 20119 12223
rect 20637 12189 20671 12223
rect 24041 12189 24075 12223
rect 24961 12189 24995 12223
rect 26249 12189 26283 12223
rect 36277 12189 36311 12223
rect 41245 12189 41279 12223
rect 45385 12189 45419 12223
rect 47409 12189 47443 12223
rect 56701 12189 56735 12223
rect 5181 12121 5215 12155
rect 6285 12121 6319 12155
rect 6622 12121 6656 12155
rect 9597 12121 9631 12155
rect 12817 12121 12851 12155
rect 17141 12121 17175 12155
rect 18889 12121 18923 12155
rect 21097 12121 21131 12155
rect 22201 12121 22235 12155
rect 25605 12121 25639 12155
rect 26516 12121 26550 12155
rect 29561 12121 29595 12155
rect 33149 12121 33183 12155
rect 40417 12121 40451 12155
rect 41512 12121 41546 12155
rect 43085 12121 43119 12155
rect 43545 12121 43579 12155
rect 44557 12121 44591 12155
rect 46397 12121 46431 12155
rect 51304 12121 51338 12155
rect 4445 12053 4479 12087
rect 7757 12053 7791 12087
rect 9229 12053 9263 12087
rect 12081 12053 12115 12087
rect 17049 12053 17083 12087
rect 19625 12053 19659 12087
rect 21833 12053 21867 12087
rect 22293 12053 22327 12087
rect 23489 12053 23523 12087
rect 24409 12053 24443 12087
rect 25881 12053 25915 12087
rect 30849 12053 30883 12087
rect 32045 12053 32079 12087
rect 35725 12053 35759 12087
rect 36645 12053 36679 12087
rect 40141 12053 40175 12087
rect 42717 12053 42751 12087
rect 43177 12053 43211 12087
rect 45293 12053 45327 12087
rect 48789 12053 48823 12087
rect 51641 12053 51675 12087
rect 56241 12053 56275 12087
rect 56793 12053 56827 12087
rect 3985 11849 4019 11883
rect 4537 11849 4571 11883
rect 5181 11849 5215 11883
rect 6101 11849 6135 11883
rect 11161 11849 11195 11883
rect 16865 11849 16899 11883
rect 18153 11849 18187 11883
rect 19993 11849 20027 11883
rect 24041 11849 24075 11883
rect 24501 11849 24535 11883
rect 26985 11849 27019 11883
rect 31125 11849 31159 11883
rect 32781 11849 32815 11883
rect 35909 11849 35943 11883
rect 36369 11849 36403 11883
rect 37105 11849 37139 11883
rect 38209 11849 38243 11883
rect 39129 11849 39163 11883
rect 39681 11849 39715 11883
rect 42441 11849 42475 11883
rect 46949 11849 46983 11883
rect 51641 11849 51675 11883
rect 54585 11849 54619 11883
rect 4169 11781 4203 11815
rect 5733 11781 5767 11815
rect 5825 11781 5859 11815
rect 6837 11781 6871 11815
rect 18512 11781 18546 11815
rect 22836 11781 22870 11815
rect 42165 11781 42199 11815
rect 43269 11781 43303 11815
rect 3901 11713 3935 11747
rect 4077 11713 4111 11747
rect 4353 11713 4387 11747
rect 4997 11713 5031 11747
rect 5549 11713 5583 11747
rect 5917 11713 5951 11747
rect 7481 11713 7515 11747
rect 7573 11713 7607 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 9597 11713 9631 11747
rect 17233 11713 17267 11747
rect 18245 11713 18279 11747
rect 21649 11713 21683 11747
rect 24409 11713 24443 11747
rect 27629 11713 27663 11747
rect 28917 11713 28951 11747
rect 35725 11713 35759 11747
rect 36277 11713 36311 11747
rect 42993 11713 43027 11747
rect 54125 11713 54159 11747
rect 4721 11645 4755 11679
rect 4813 11645 4847 11679
rect 4905 11645 4939 11679
rect 7665 11645 7699 11679
rect 9873 11645 9907 11679
rect 15025 11645 15059 11679
rect 17325 11645 17359 11679
rect 17417 11645 17451 11679
rect 20821 11645 20855 11679
rect 21833 11645 21867 11679
rect 22477 11645 22511 11679
rect 22569 11645 22603 11679
rect 24593 11645 24627 11679
rect 25513 11645 25547 11679
rect 29285 11645 29319 11679
rect 30665 11645 30699 11679
rect 33149 11645 33183 11679
rect 34437 11645 34471 11679
rect 36461 11645 36495 11679
rect 37841 11645 37875 11679
rect 39405 11645 39439 11679
rect 39589 11645 39623 11679
rect 45109 11645 45143 11679
rect 45661 11645 45695 11679
rect 48421 11645 48455 11679
rect 51273 11645 51307 11679
rect 57161 11645 57195 11679
rect 19625 11577 19659 11611
rect 23949 11577 23983 11611
rect 28365 11577 28399 11611
rect 32413 11577 32447 11611
rect 37289 11577 37323 11611
rect 44557 11577 44591 11611
rect 7573 11509 7607 11543
rect 7941 11509 7975 11543
rect 8861 11509 8895 11543
rect 9045 11509 9079 11543
rect 9321 11509 9355 11543
rect 14473 11509 14507 11543
rect 16405 11509 16439 11543
rect 20269 11509 20303 11543
rect 21005 11509 21039 11543
rect 26157 11509 26191 11543
rect 26525 11509 26559 11543
rect 28825 11509 28859 11543
rect 30021 11509 30055 11543
rect 33793 11509 33827 11543
rect 33885 11509 33919 11543
rect 40049 11509 40083 11543
rect 47777 11509 47811 11543
rect 50261 11509 50295 11543
rect 50537 11509 50571 11543
rect 50721 11509 50755 11543
rect 56609 11509 56643 11543
rect 3433 11305 3467 11339
rect 3617 11305 3651 11339
rect 3985 11305 4019 11339
rect 4169 11305 4203 11339
rect 5549 11305 5583 11339
rect 11529 11305 11563 11339
rect 12173 11305 12207 11339
rect 13737 11305 13771 11339
rect 18429 11305 18463 11339
rect 19441 11305 19475 11339
rect 23305 11305 23339 11339
rect 25237 11305 25271 11339
rect 30941 11305 30975 11339
rect 37473 11305 37507 11339
rect 43729 11305 43763 11339
rect 50905 11305 50939 11339
rect 52929 11305 52963 11339
rect 10609 11237 10643 11271
rect 13553 11237 13587 11271
rect 15485 11237 15519 11271
rect 22569 11237 22603 11271
rect 36277 11237 36311 11271
rect 37565 11237 37599 11271
rect 38761 11237 38795 11271
rect 42625 11237 42659 11271
rect 44741 11237 44775 11271
rect 47869 11237 47903 11271
rect 50997 11237 51031 11271
rect 54401 11237 54435 11271
rect 4537 11169 4571 11203
rect 5641 11169 5675 11203
rect 16129 11169 16163 11203
rect 18337 11169 18371 11203
rect 21189 11169 21223 11203
rect 23857 11169 23891 11203
rect 26617 11169 26651 11203
rect 27261 11169 27295 11203
rect 28825 11169 28859 11203
rect 28917 11169 28951 11203
rect 34897 11169 34931 11203
rect 36921 11169 36955 11203
rect 38209 11169 38243 11203
rect 38368 11169 38402 11203
rect 39221 11169 39255 11203
rect 40417 11169 40451 11203
rect 41981 11169 42015 11203
rect 43177 11169 43211 11203
rect 44189 11169 44223 11203
rect 44281 11169 44315 11203
rect 46305 11169 46339 11203
rect 47225 11169 47259 11203
rect 49985 11169 50019 11203
rect 50353 11169 50387 11203
rect 50445 11169 50479 11203
rect 51549 11169 51583 11203
rect 51825 11169 51859 11203
rect 3341 11101 3375 11135
rect 4069 11103 4103 11137
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 4905 11101 4939 11135
rect 5273 11101 5307 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9413 11101 9447 11135
rect 10149 11101 10183 11135
rect 10517 11101 10551 11135
rect 11437 11101 11471 11135
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 14105 11101 14139 11135
rect 16865 11101 16899 11135
rect 18981 11101 19015 11135
rect 19717 11101 19751 11135
rect 21445 11101 21479 11135
rect 22937 11101 22971 11135
rect 25145 11101 25179 11135
rect 28549 11101 28583 11135
rect 29561 11101 29595 11135
rect 31217 11101 31251 11135
rect 32413 11101 32447 11135
rect 33333 11101 33367 11135
rect 38485 11101 38519 11135
rect 39405 11101 39439 11135
rect 41797 11101 41831 11135
rect 43085 11101 43119 11135
rect 45569 11101 45603 11135
rect 47409 11101 47443 11135
rect 48513 11101 48547 11135
rect 51365 11101 51399 11135
rect 53021 11101 53055 11135
rect 54493 11101 54527 11135
rect 55045 11101 55079 11135
rect 56241 11101 56275 11135
rect 56333 11101 56367 11135
rect 56600 11101 56634 11135
rect 58357 11101 58391 11135
rect 3249 11033 3283 11067
rect 3617 11033 3651 11067
rect 8033 11033 8067 11067
rect 8769 11033 8803 11067
rect 10793 11033 10827 11067
rect 11161 11033 11195 11067
rect 13829 11033 13863 11067
rect 14361 11033 14395 11067
rect 15577 11033 15611 11067
rect 18070 11033 18104 11067
rect 19984 11033 20018 11067
rect 26350 11033 26384 11067
rect 29828 11033 29862 11067
rect 31953 11033 31987 11067
rect 33057 11033 33091 11067
rect 34161 11033 34195 11067
rect 35164 11033 35198 11067
rect 36737 11033 36771 11067
rect 45017 11033 45051 11067
rect 47501 11033 47535 11067
rect 50537 11033 50571 11067
rect 51457 11033 51491 11067
rect 53288 11033 53322 11067
rect 57805 11033 57839 11067
rect 5365 10965 5399 10999
rect 5457 10965 5491 10999
rect 9045 10965 9079 10999
rect 11713 10965 11747 10999
rect 16957 10965 16991 10999
rect 21097 10965 21131 10999
rect 26709 10965 26743 10999
rect 27721 10965 27755 10999
rect 27905 10965 27939 10999
rect 29009 10965 29043 10999
rect 29377 10965 29411 10999
rect 36369 10965 36403 10999
rect 36829 10965 36863 10999
rect 39865 10965 39899 10999
rect 42533 10965 42567 10999
rect 42993 10965 43027 10999
rect 44373 10965 44407 10999
rect 45753 10965 45787 10999
rect 46673 10965 46707 10999
rect 47961 10965 47995 10999
rect 48881 10965 48915 10999
rect 52469 10965 52503 10999
rect 57713 10965 57747 10999
rect 5641 10761 5675 10795
rect 11345 10761 11379 10795
rect 14565 10761 14599 10795
rect 15025 10761 15059 10795
rect 18061 10761 18095 10795
rect 20453 10761 20487 10795
rect 20913 10761 20947 10795
rect 22845 10761 22879 10795
rect 25421 10761 25455 10795
rect 25789 10761 25823 10795
rect 30021 10761 30055 10795
rect 40509 10761 40543 10795
rect 41337 10761 41371 10795
rect 42165 10761 42199 10795
rect 45293 10761 45327 10795
rect 47869 10761 47903 10795
rect 48329 10761 48363 10795
rect 50813 10761 50847 10795
rect 4169 10693 4203 10727
rect 9873 10693 9907 10727
rect 16948 10693 16982 10727
rect 21557 10693 21591 10727
rect 28150 10693 28184 10727
rect 33272 10693 33306 10727
rect 34069 10693 34103 10727
rect 35440 10693 35474 10727
rect 36921 10693 36955 10727
rect 39037 10693 39071 10727
rect 44180 10693 44214 10727
rect 46296 10693 46330 10727
rect 51948 10693 51982 10727
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 3433 10625 3467 10659
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 8861 10625 8895 10659
rect 10221 10625 10255 10659
rect 13360 10625 13394 10659
rect 14933 10625 14967 10659
rect 19993 10625 20027 10659
rect 20821 10625 20855 10659
rect 21833 10625 21867 10659
rect 23673 10625 23707 10659
rect 23949 10625 23983 10659
rect 24685 10625 24719 10659
rect 24869 10625 24903 10659
rect 29377 10625 29411 10659
rect 30916 10625 30950 10659
rect 31033 10625 31067 10659
rect 33517 10625 33551 10659
rect 33977 10625 34011 10659
rect 35173 10625 35207 10659
rect 37565 10625 37599 10659
rect 37821 10625 37855 10659
rect 42441 10625 42475 10659
rect 42697 10625 42731 10659
rect 43913 10625 43947 10659
rect 47961 10625 47995 10659
rect 49525 10625 49559 10659
rect 49801 10625 49835 10659
rect 50721 10625 50755 10659
rect 52193 10625 52227 10659
rect 52561 10625 52595 10659
rect 52929 10625 52963 10659
rect 53196 10625 53230 10659
rect 55137 10625 55171 10659
rect 55413 10625 55447 10659
rect 56149 10625 56183 10659
rect 56793 10625 56827 10659
rect 3525 10557 3559 10591
rect 8493 10557 8527 10591
rect 9045 10557 9079 10591
rect 9965 10557 9999 10591
rect 13093 10557 13127 10591
rect 15117 10557 15151 10591
rect 15945 10557 15979 10591
rect 16681 10557 16715 10591
rect 20361 10557 20395 10591
rect 21097 10557 21131 10591
rect 22477 10557 22511 10591
rect 23811 10557 23845 10591
rect 24225 10557 24259 10591
rect 25881 10557 25915 10591
rect 25973 10557 26007 10591
rect 27905 10557 27939 10591
rect 30757 10557 30791 10591
rect 31309 10557 31343 10591
rect 31769 10557 31803 10591
rect 31953 10557 31987 10591
rect 34253 10557 34287 10591
rect 45661 10557 45695 10591
rect 46029 10557 46063 10591
rect 47685 10557 47719 10591
rect 49663 10557 49697 10591
rect 50077 10557 50111 10591
rect 50537 10557 50571 10591
rect 55275 10557 55309 10591
rect 56333 10557 56367 10591
rect 56517 10557 56551 10591
rect 56701 10557 56735 10591
rect 58449 10557 58483 10591
rect 2881 10489 2915 10523
rect 3801 10489 3835 10523
rect 4353 10489 4387 10523
rect 13001 10489 13035 10523
rect 14473 10489 14507 10523
rect 33609 10489 33643 10523
rect 36553 10489 36587 10523
rect 38945 10489 38979 10523
rect 47409 10489 47443 10523
rect 54309 10489 54343 10523
rect 55689 10489 55723 10523
rect 57161 10489 57195 10523
rect 6653 10421 6687 10455
rect 15393 10421 15427 10455
rect 18705 10421 18739 10455
rect 23029 10421 23063 10455
rect 25329 10421 25363 10455
rect 29285 10421 29319 10455
rect 30113 10421 30147 10455
rect 32137 10421 32171 10455
rect 34713 10421 34747 10455
rect 43821 10421 43855 10455
rect 48605 10421 48639 10455
rect 48881 10421 48915 10455
rect 54493 10421 54527 10455
rect 57437 10421 57471 10455
rect 57897 10421 57931 10455
rect 3157 10217 3191 10251
rect 6745 10217 6779 10251
rect 7757 10217 7791 10251
rect 9321 10217 9355 10251
rect 9689 10217 9723 10251
rect 13277 10217 13311 10251
rect 19625 10217 19659 10251
rect 20545 10217 20579 10251
rect 26525 10217 26559 10251
rect 28549 10217 28583 10251
rect 35817 10217 35851 10251
rect 36553 10217 36587 10251
rect 37473 10217 37507 10251
rect 39405 10217 39439 10251
rect 46213 10217 46247 10251
rect 51641 10217 51675 10251
rect 53297 10217 53331 10251
rect 54861 10217 54895 10251
rect 57713 10217 57747 10251
rect 6101 10149 6135 10183
rect 7941 10149 7975 10183
rect 9597 10149 9631 10183
rect 14105 10149 14139 10183
rect 20361 10149 20395 10183
rect 21557 10149 21591 10183
rect 25329 10149 25363 10183
rect 37657 10149 37691 10183
rect 38393 10149 38427 10183
rect 39865 10149 39899 10183
rect 42717 10149 42751 10183
rect 47869 10149 47903 10183
rect 52837 10149 52871 10183
rect 2881 10081 2915 10115
rect 4077 10081 4111 10115
rect 13921 10081 13955 10115
rect 14565 10081 14599 10115
rect 14749 10081 14783 10115
rect 16359 10081 16393 10115
rect 16497 10081 16531 10115
rect 16773 10081 16807 10115
rect 17233 10081 17267 10115
rect 18061 10081 18095 10115
rect 21005 10081 21039 10115
rect 21097 10081 21131 10115
rect 22937 10081 22971 10115
rect 23949 10081 23983 10115
rect 24777 10081 24811 10115
rect 25605 10081 25639 10115
rect 29101 10081 29135 10115
rect 30113 10081 30147 10115
rect 36369 10081 36403 10115
rect 37105 10081 37139 10115
rect 38301 10081 38335 10115
rect 38945 10081 38979 10115
rect 41245 10081 41279 10115
rect 41337 10081 41371 10115
rect 43775 10081 43809 10115
rect 43913 10081 43947 10115
rect 44189 10081 44223 10115
rect 44833 10081 44867 10115
rect 48973 10081 49007 10115
rect 51549 10081 51583 10115
rect 53849 10081 53883 10115
rect 54309 10081 54343 10115
rect 55873 10081 55907 10115
rect 2513 10013 2547 10047
rect 2667 10013 2701 10047
rect 3248 10013 3282 10047
rect 3341 10013 3375 10047
rect 6345 10013 6379 10047
rect 6469 10013 6503 10047
rect 6836 10013 6870 10047
rect 6929 10013 6963 10047
rect 8125 10013 8159 10047
rect 8953 10013 8987 10047
rect 9123 10013 9157 10047
rect 9689 10013 9723 10047
rect 12817 10013 12851 10047
rect 14473 10013 14507 10047
rect 16221 10013 16255 10047
rect 17417 10013 17451 10047
rect 18889 10013 18923 10047
rect 22293 10013 22327 10047
rect 24961 10013 24995 10047
rect 26709 10013 26743 10047
rect 33333 10013 33367 10047
rect 33977 10013 34011 10047
rect 38761 10013 38795 10047
rect 43637 10013 43671 10047
rect 44649 10013 44683 10047
rect 45937 10013 45971 10047
rect 46489 10013 46523 10047
rect 48513 10013 48547 10047
rect 49617 10013 49651 10047
rect 52193 10013 52227 10047
rect 57365 10013 57399 10047
rect 57621 10013 57655 10047
rect 58265 10013 58299 10047
rect 7573 9945 7607 9979
rect 7789 9945 7823 9979
rect 8677 9945 8711 9979
rect 9413 9945 9447 9979
rect 10333 9945 10367 9979
rect 15393 9945 15427 9979
rect 17877 9945 17911 9979
rect 18337 9945 18371 9979
rect 20637 9945 20671 9979
rect 21189 9945 21223 9979
rect 21649 9945 21683 9979
rect 23673 9945 23707 9979
rect 28917 9945 28951 9979
rect 29561 9945 29595 9979
rect 33088 9945 33122 9979
rect 41000 9945 41034 9979
rect 41604 9945 41638 9979
rect 45109 9945 45143 9979
rect 46756 9945 46790 9979
rect 47961 9945 47995 9979
rect 49433 9945 49467 9979
rect 51304 9945 51338 9979
rect 53665 9945 53699 9979
rect 54401 9945 54435 9979
rect 55321 9945 55355 9979
rect 7481 9877 7515 9911
rect 9965 9877 9999 9911
rect 12265 9877 12299 9911
rect 15577 9877 15611 9911
rect 17509 9877 17543 9911
rect 17969 9877 18003 9911
rect 22385 9877 22419 9911
rect 23305 9877 23339 9911
rect 23765 9877 23799 9911
rect 24869 9877 24903 9911
rect 27997 9877 28031 9911
rect 29009 9877 29043 9911
rect 30481 9877 30515 9911
rect 31401 9877 31435 9911
rect 31861 9877 31895 9911
rect 31953 9877 31987 9911
rect 33425 9877 33459 9911
rect 38853 9877 38887 9911
rect 42993 9877 43027 9911
rect 49985 9877 50019 9911
rect 50169 9877 50203 9911
rect 53113 9877 53147 9911
rect 53757 9877 53791 9911
rect 54493 9877 54527 9911
rect 56241 9877 56275 9911
rect 3065 9673 3099 9707
rect 12265 9673 12299 9707
rect 19625 9673 19659 9707
rect 32965 9673 32999 9707
rect 41153 9673 41187 9707
rect 41613 9673 41647 9707
rect 43453 9673 43487 9707
rect 45477 9673 45511 9707
rect 49065 9673 49099 9707
rect 50629 9673 50663 9707
rect 51825 9673 51859 9707
rect 53297 9673 53331 9707
rect 4629 9605 4663 9639
rect 6745 9605 6779 9639
rect 7849 9605 7883 9639
rect 8217 9605 8251 9639
rect 9229 9605 9263 9639
rect 12633 9605 12667 9639
rect 14197 9605 14231 9639
rect 18153 9605 18187 9639
rect 18521 9605 18555 9639
rect 20444 9605 20478 9639
rect 22201 9605 22235 9639
rect 28549 9605 28583 9639
rect 31309 9605 31343 9639
rect 32505 9605 32539 9639
rect 36369 9605 36403 9639
rect 39313 9605 39347 9639
rect 44373 9605 44407 9639
rect 45385 9605 45419 9639
rect 47777 9605 47811 9639
rect 56885 9605 56919 9639
rect 58265 9605 58299 9639
rect 3801 9537 3835 9571
rect 3985 9537 4019 9571
rect 4353 9537 4387 9571
rect 4997 9537 5031 9571
rect 5365 9537 5399 9571
rect 6561 9537 6595 9571
rect 7941 9537 7975 9571
rect 8033 9537 8067 9571
rect 8585 9537 8619 9571
rect 10618 9537 10652 9571
rect 13093 9537 13127 9571
rect 17049 9537 17083 9571
rect 17509 9537 17543 9571
rect 20177 9537 20211 9571
rect 23489 9537 23523 9571
rect 24501 9537 24535 9571
rect 26074 9537 26108 9571
rect 28641 9537 28675 9571
rect 29009 9537 29043 9571
rect 29653 9537 29687 9571
rect 30573 9537 30607 9571
rect 30757 9537 30791 9571
rect 32597 9537 32631 9571
rect 33057 9537 33091 9571
rect 33609 9537 33643 9571
rect 34069 9537 34103 9571
rect 36553 9537 36587 9571
rect 38853 9537 38887 9571
rect 40325 9537 40359 9571
rect 42809 9537 42843 9571
rect 42901 9537 42935 9571
rect 44005 9537 44039 9571
rect 48421 9537 48455 9571
rect 51181 9537 51215 9571
rect 53849 9537 53883 9571
rect 54033 9537 54067 9571
rect 54585 9537 54619 9571
rect 57529 9537 57563 9571
rect 58081 9537 58115 9571
rect 58449 9537 58483 9571
rect 8861 9469 8895 9503
rect 10885 9469 10919 9503
rect 12725 9469 12759 9503
rect 12817 9469 12851 9503
rect 13461 9469 13495 9503
rect 14749 9469 14783 9503
rect 15301 9469 15335 9503
rect 16773 9469 16807 9503
rect 16957 9469 16991 9503
rect 21925 9469 21959 9503
rect 22109 9469 22143 9503
rect 23627 9469 23661 9503
rect 23765 9469 23799 9503
rect 24041 9469 24075 9503
rect 24685 9469 24719 9503
rect 26341 9469 26375 9503
rect 27445 9469 27479 9503
rect 28089 9469 28123 9503
rect 28733 9469 28767 9503
rect 32413 9469 32447 9503
rect 35357 9469 35391 9503
rect 39037 9469 39071 9503
rect 39221 9469 39255 9503
rect 39773 9469 39807 9503
rect 40509 9469 40543 9503
rect 42257 9469 42291 9503
rect 42993 9469 43027 9503
rect 45569 9469 45603 9503
rect 46949 9469 46983 9503
rect 55597 9469 55631 9503
rect 55873 9469 55907 9503
rect 56977 9469 57011 9503
rect 57069 9469 57103 9503
rect 6101 9401 6135 9435
rect 8217 9401 8251 9435
rect 8677 9401 8711 9435
rect 9505 9401 9539 9435
rect 11805 9401 11839 9435
rect 21557 9401 21591 9435
rect 26709 9401 26743 9435
rect 28181 9401 28215 9435
rect 38669 9401 38703 9435
rect 39681 9401 39715 9435
rect 42441 9401 42475 9435
rect 7021 9333 7055 9367
rect 8769 9333 8803 9367
rect 12081 9333 12115 9367
rect 15577 9333 15611 9367
rect 16037 9333 16071 9367
rect 16405 9333 16439 9367
rect 17417 9333 17451 9367
rect 20085 9333 20119 9367
rect 22569 9333 22603 9367
rect 22845 9333 22879 9367
rect 24961 9333 24995 9367
rect 29929 9333 29963 9367
rect 31861 9333 31895 9367
rect 34345 9333 34379 9367
rect 35909 9333 35943 9367
rect 37841 9333 37875 9367
rect 38209 9333 38243 9367
rect 45017 9333 45051 9367
rect 46029 9333 46063 9367
rect 46397 9333 46431 9367
rect 47317 9333 47351 9367
rect 48697 9333 48731 9367
rect 49985 9333 50019 9367
rect 53021 9333 53055 9367
rect 55137 9333 55171 9367
rect 56425 9333 56459 9367
rect 56517 9333 56551 9367
rect 4813 9129 4847 9163
rect 5549 9129 5583 9163
rect 8401 9129 8435 9163
rect 13369 9129 13403 9163
rect 18797 9129 18831 9163
rect 22017 9129 22051 9163
rect 24409 9129 24443 9163
rect 28825 9129 28859 9163
rect 37565 9129 37599 9163
rect 42809 9129 42843 9163
rect 43729 9129 43763 9163
rect 44557 9129 44591 9163
rect 46581 9129 46615 9163
rect 51457 9129 51491 9163
rect 53849 9129 53883 9163
rect 56517 9129 56551 9163
rect 3341 9061 3375 9095
rect 4905 9061 4939 9095
rect 13829 9061 13863 9095
rect 21741 9061 21775 9095
rect 24133 9061 24167 9095
rect 29285 9061 29319 9095
rect 45569 9061 45603 9095
rect 49709 9061 49743 9095
rect 53021 9061 53055 9095
rect 56333 9061 56367 9095
rect 58357 9061 58391 9095
rect 4353 8993 4387 9027
rect 7481 8993 7515 9027
rect 9045 8993 9079 9027
rect 15531 8993 15565 9027
rect 15669 8993 15703 9027
rect 15945 8993 15979 9027
rect 18429 8993 18463 9027
rect 22661 8993 22695 9027
rect 24961 8993 24995 9027
rect 25697 8993 25731 9027
rect 25881 8993 25915 9027
rect 26617 8993 26651 9027
rect 31125 8993 31159 9027
rect 31217 8993 31251 9027
rect 39037 8993 39071 9027
rect 43453 8993 43487 9027
rect 45201 8993 45235 9027
rect 47133 8993 47167 9027
rect 49249 8993 49283 9027
rect 50261 8993 50295 9027
rect 52377 8993 52411 9027
rect 53573 8993 53607 9027
rect 54401 8993 54435 9027
rect 54861 8993 54895 9027
rect 57069 8993 57103 9027
rect 57529 8993 57563 9027
rect 1961 8925 1995 8959
rect 5273 8925 5307 8959
rect 9505 8925 9539 8959
rect 9873 8925 9907 8959
rect 11621 8925 11655 8959
rect 11989 8925 12023 8959
rect 12256 8925 12290 8959
rect 15393 8925 15427 8959
rect 16405 8925 16439 8959
rect 16589 8925 16623 8959
rect 20361 8925 20395 8959
rect 22753 8925 22787 8959
rect 27445 8925 27479 8959
rect 27712 8925 27746 8959
rect 29561 8925 29595 8959
rect 31769 8925 31803 8959
rect 32873 8925 32907 8959
rect 33425 8925 33459 8959
rect 34713 8925 34747 8959
rect 36737 8925 36771 8959
rect 38945 8925 38979 8959
rect 40417 8925 40451 8959
rect 48053 8925 48087 8959
rect 54309 8925 54343 8959
rect 55873 8925 55907 8959
rect 2228 8857 2262 8891
rect 9137 8857 9171 8891
rect 9597 8857 9631 8891
rect 18162 8857 18196 8891
rect 20628 8857 20662 8891
rect 23020 8857 23054 8891
rect 25605 8857 25639 8891
rect 26065 8857 26099 8891
rect 30389 8857 30423 8891
rect 32597 8857 32631 8891
rect 34980 8857 35014 8891
rect 36185 8857 36219 8891
rect 38700 8857 38734 8891
rect 39865 8857 39899 8891
rect 44465 8857 44499 8891
rect 46949 8857 46983 8891
rect 49065 8857 49099 8891
rect 50445 8857 50479 8891
rect 50537 8857 50571 8891
rect 51549 8857 51583 8891
rect 53389 8857 53423 8891
rect 55321 8857 55355 8891
rect 56977 8857 57011 8891
rect 3801 8789 3835 8823
rect 6929 8789 6963 8823
rect 14289 8789 14323 8823
rect 14749 8789 14783 8823
rect 17049 8789 17083 8823
rect 25237 8789 25271 8823
rect 31309 8789 31343 8823
rect 31677 8789 31711 8823
rect 33793 8789 33827 8823
rect 34437 8789 34471 8823
rect 36093 8789 36127 8823
rect 39681 8789 39715 8823
rect 40785 8789 40819 8823
rect 41153 8789 41187 8823
rect 42349 8789 42383 8823
rect 44281 8789 44315 8823
rect 45937 8789 45971 8823
rect 46305 8789 46339 8823
rect 47041 8789 47075 8823
rect 47409 8789 47443 8823
rect 48329 8789 48363 8823
rect 48697 8789 48731 8823
rect 49157 8789 49191 8823
rect 50905 8789 50939 8823
rect 52929 8789 52963 8823
rect 53481 8789 53515 8823
rect 54217 8789 54251 8823
rect 56885 8789 56919 8823
rect 57621 8789 57655 8823
rect 57713 8789 57747 8823
rect 58081 8789 58115 8823
rect 2421 8585 2455 8619
rect 3985 8585 4019 8619
rect 5733 8585 5767 8619
rect 7757 8585 7791 8619
rect 9873 8585 9907 8619
rect 10057 8585 10091 8619
rect 13277 8585 13311 8619
rect 16037 8585 16071 8619
rect 17785 8585 17819 8619
rect 21833 8585 21867 8619
rect 23213 8585 23247 8619
rect 25881 8585 25915 8619
rect 29929 8585 29963 8619
rect 32137 8585 32171 8619
rect 36001 8585 36035 8619
rect 36461 8585 36495 8619
rect 39129 8585 39163 8619
rect 39773 8585 39807 8619
rect 44833 8585 44867 8619
rect 47225 8585 47259 8619
rect 48421 8585 48455 8619
rect 50629 8585 50663 8619
rect 51181 8585 51215 8619
rect 54217 8585 54251 8619
rect 57621 8585 57655 8619
rect 57897 8585 57931 8619
rect 2237 8517 2271 8551
rect 4169 8517 4203 8551
rect 5549 8517 5583 8551
rect 9689 8517 9723 8551
rect 27721 8517 27755 8551
rect 28058 8517 28092 8551
rect 40509 8517 40543 8551
rect 46112 8517 46146 8551
rect 47869 8517 47903 8551
rect 50721 8517 50755 8551
rect 2053 8449 2087 8483
rect 2329 8449 2363 8483
rect 3249 8449 3283 8483
rect 4353 8449 4387 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 8309 8449 8343 8483
rect 8769 8449 8803 8483
rect 8953 8449 8987 8483
rect 9597 8449 9631 8483
rect 11904 8449 11938 8483
rect 12164 8449 12198 8483
rect 13369 8449 13403 8483
rect 14657 8449 14691 8483
rect 14924 8449 14958 8483
rect 17693 8449 17727 8483
rect 18153 8449 18187 8483
rect 18705 8449 18739 8483
rect 22477 8449 22511 8483
rect 23765 8449 23799 8483
rect 25237 8449 25271 8483
rect 27169 8449 27203 8483
rect 30573 8449 30607 8483
rect 30849 8449 30883 8483
rect 31585 8449 31619 8483
rect 33261 8449 33295 8483
rect 33517 8449 33551 8483
rect 34253 8449 34287 8483
rect 34520 8449 34554 8483
rect 36093 8449 36127 8483
rect 36737 8449 36771 8483
rect 38402 8449 38436 8483
rect 38669 8449 38703 8483
rect 39681 8449 39715 8483
rect 43453 8449 43487 8483
rect 43720 8449 43754 8483
rect 44925 8449 44959 8483
rect 47961 8449 47995 8483
rect 49065 8449 49099 8483
rect 49341 8449 49375 8483
rect 52469 8449 52503 8483
rect 52745 8449 52779 8483
rect 53001 8449 53035 8483
rect 54861 8449 54895 8483
rect 56057 8449 56091 8483
rect 56497 8449 56531 8483
rect 58449 8449 58483 8483
rect 2973 8381 3007 8415
rect 3893 8381 3927 8415
rect 6377 8381 6411 8415
rect 6653 8381 6687 8415
rect 13737 8381 13771 8415
rect 17877 8381 17911 8415
rect 19441 8381 19475 8415
rect 22845 8381 22879 8415
rect 25145 8381 25179 8415
rect 27813 8381 27847 8415
rect 30711 8381 30745 8415
rect 31769 8381 31803 8415
rect 35909 8381 35943 8415
rect 38945 8381 38979 8415
rect 39037 8381 39071 8415
rect 40233 8381 40267 8415
rect 41429 8381 41463 8415
rect 42257 8381 42291 8415
rect 42993 8381 43027 8415
rect 45569 8381 45603 8415
rect 45845 8381 45879 8415
rect 47777 8381 47811 8415
rect 49224 8381 49258 8415
rect 49617 8381 49651 8415
rect 50077 8381 50111 8415
rect 50261 8381 50295 8415
rect 50445 8381 50479 8415
rect 51733 8381 51767 8415
rect 54999 8381 55033 8415
rect 55137 8381 55171 8415
rect 55413 8381 55447 8415
rect 55873 8381 55907 8415
rect 56241 8381 56275 8415
rect 2053 8313 2087 8347
rect 5181 8313 5215 8347
rect 10425 8313 10459 8347
rect 11345 8313 11379 8347
rect 17141 8313 17175 8347
rect 26709 8313 26743 8347
rect 29193 8313 29227 8347
rect 29561 8313 29595 8347
rect 31125 8313 31159 8347
rect 33793 8313 33827 8347
rect 39497 8313 39531 8347
rect 42441 8313 42475 8347
rect 51089 8313 51123 8347
rect 54125 8313 54159 8347
rect 5549 8245 5583 8279
rect 5917 8245 5951 8279
rect 9873 8245 9907 8279
rect 11805 8245 11839 8279
rect 17325 8245 17359 8279
rect 20085 8245 20119 8279
rect 21649 8245 21683 8279
rect 24225 8245 24259 8279
rect 35633 8245 35667 8279
rect 37289 8245 37323 8279
rect 40877 8245 40911 8279
rect 41613 8245 41647 8279
rect 48329 8245 48363 8279
rect 51917 8245 51951 8279
rect 3893 8041 3927 8075
rect 4445 8041 4479 8075
rect 5549 8041 5583 8075
rect 10149 8041 10183 8075
rect 10885 8041 10919 8075
rect 11897 8041 11931 8075
rect 13645 8041 13679 8075
rect 17969 8041 18003 8075
rect 33609 8041 33643 8075
rect 41797 8041 41831 8075
rect 44741 8041 44775 8075
rect 47961 8041 47995 8075
rect 49525 8041 49559 8075
rect 53941 8041 53975 8075
rect 4629 7973 4663 8007
rect 8309 7973 8343 8007
rect 12633 7973 12667 8007
rect 18705 7973 18739 8007
rect 22569 7973 22603 8007
rect 25789 7973 25823 8007
rect 32781 7973 32815 8007
rect 50169 7973 50203 8007
rect 54953 7973 54987 8007
rect 7849 7905 7883 7939
rect 8401 7905 8435 7939
rect 8769 7905 8803 7939
rect 12541 7905 12575 7939
rect 13185 7905 13219 7939
rect 14749 7905 14783 7939
rect 15209 7905 15243 7939
rect 16589 7905 16623 7939
rect 17325 7905 17359 7939
rect 18981 7905 19015 7939
rect 29377 7905 29411 7939
rect 31769 7905 31803 7939
rect 32229 7905 32263 7939
rect 32321 7905 32355 7939
rect 34161 7905 34195 7939
rect 35541 7905 35575 7939
rect 36921 7905 36955 7939
rect 37197 7905 37231 7939
rect 37657 7905 37691 7939
rect 37841 7905 37875 7939
rect 38485 7905 38519 7939
rect 44189 7905 44223 7939
rect 45569 7905 45603 7939
rect 47225 7905 47259 7939
rect 51549 7905 51583 7939
rect 52561 7905 52595 7939
rect 54585 7905 54619 7939
rect 55781 7905 55815 7939
rect 55873 7905 55907 7939
rect 57713 7905 57747 7939
rect 58357 7905 58391 7939
rect 2789 7837 2823 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 5181 7837 5215 7871
rect 7941 7837 7975 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 11621 7837 11655 7871
rect 13001 7837 13035 7871
rect 15485 7837 15519 7871
rect 20637 7837 20671 7871
rect 21281 7837 21315 7871
rect 23581 7837 23615 7871
rect 26525 7837 26559 7871
rect 26893 7837 26927 7871
rect 30021 7837 30055 7871
rect 32413 7837 32447 7871
rect 33425 7837 33459 7871
rect 35357 7837 35391 7871
rect 36645 7837 36679 7871
rect 36783 7837 36817 7871
rect 39313 7837 39347 7871
rect 40417 7837 40451 7871
rect 41889 7837 41923 7871
rect 42156 7837 42190 7871
rect 47409 7837 47443 7871
rect 48145 7837 48179 7871
rect 52469 7837 52503 7871
rect 55689 7837 55723 7871
rect 3433 7769 3467 7803
rect 4261 7769 4295 7803
rect 5365 7769 5399 7803
rect 9137 7769 9171 7803
rect 9597 7769 9631 7803
rect 13093 7769 13127 7803
rect 14105 7769 14139 7803
rect 15393 7769 15427 7803
rect 15945 7769 15979 7803
rect 18521 7769 18555 7803
rect 20392 7769 20426 7803
rect 20729 7769 20763 7803
rect 30288 7769 30322 7803
rect 38301 7769 38335 7803
rect 40049 7769 40083 7803
rect 40684 7769 40718 7803
rect 44373 7769 44407 7803
rect 45017 7769 45051 7803
rect 46980 7769 47014 7803
rect 48412 7769 48446 7803
rect 51304 7769 51338 7803
rect 52828 7769 52862 7803
rect 54033 7769 54067 7803
rect 57468 7769 57502 7803
rect 57805 7769 57839 7803
rect 4471 7701 4505 7735
rect 7297 7701 7331 7735
rect 7573 7701 7607 7735
rect 10517 7701 10551 7735
rect 11069 7701 11103 7735
rect 15853 7701 15887 7735
rect 19257 7701 19291 7735
rect 23029 7701 23063 7735
rect 24041 7701 24075 7735
rect 25973 7701 26007 7735
rect 28181 7701 28215 7735
rect 28733 7701 28767 7735
rect 29837 7701 29871 7735
rect 31401 7701 31435 7735
rect 32873 7701 32907 7735
rect 34897 7701 34931 7735
rect 35265 7701 35299 7735
rect 36001 7701 36035 7735
rect 37933 7701 37967 7735
rect 38393 7701 38427 7735
rect 38761 7701 38795 7735
rect 43269 7701 43303 7735
rect 43637 7701 43671 7735
rect 44281 7701 44315 7735
rect 45845 7701 45879 7735
rect 49893 7701 49927 7735
rect 52009 7701 52043 7735
rect 55321 7701 55355 7735
rect 56333 7701 56367 7735
rect 5825 7497 5859 7531
rect 6193 7497 6227 7531
rect 12817 7497 12851 7531
rect 15025 7497 15059 7531
rect 28457 7497 28491 7531
rect 28825 7497 28859 7531
rect 29745 7497 29779 7531
rect 31861 7497 31895 7531
rect 32413 7497 32447 7531
rect 34253 7497 34287 7531
rect 34713 7497 34747 7531
rect 35541 7497 35575 7531
rect 36829 7497 36863 7531
rect 38393 7497 38427 7531
rect 40877 7497 40911 7531
rect 41061 7497 41095 7531
rect 41521 7497 41555 7531
rect 42441 7497 42475 7531
rect 44925 7497 44959 7531
rect 46765 7497 46799 7531
rect 47593 7497 47627 7531
rect 48605 7497 48639 7531
rect 49341 7497 49375 7531
rect 53481 7497 53515 7531
rect 54125 7497 54159 7531
rect 57253 7497 57287 7531
rect 57621 7497 57655 7531
rect 57897 7497 57931 7531
rect 2605 7429 2639 7463
rect 4537 7429 4571 7463
rect 5273 7429 5307 7463
rect 10609 7429 10643 7463
rect 11529 7429 11563 7463
rect 20821 7429 20855 7463
rect 24685 7429 24719 7463
rect 25504 7429 25538 7463
rect 42165 7429 42199 7463
rect 53849 7429 53883 7463
rect 55873 7429 55907 7463
rect 2237 7361 2271 7395
rect 3525 7361 3559 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 6653 7361 6687 7395
rect 8861 7361 8895 7395
rect 9091 7361 9125 7395
rect 9597 7361 9631 7395
rect 9965 7361 9999 7395
rect 13737 7361 13771 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 15669 7361 15703 7395
rect 17417 7361 17451 7395
rect 17601 7361 17635 7395
rect 19441 7361 19475 7395
rect 19533 7361 19567 7395
rect 22201 7361 22235 7395
rect 22468 7361 22502 7395
rect 25237 7361 25271 7395
rect 28917 7361 28951 7395
rect 29837 7361 29871 7395
rect 30941 7361 30975 7395
rect 32689 7361 32723 7395
rect 33977 7361 34011 7395
rect 34345 7361 34379 7395
rect 35265 7361 35299 7395
rect 37841 7361 37875 7395
rect 39681 7361 39715 7395
rect 41429 7361 41463 7395
rect 42809 7361 42843 7395
rect 42901 7361 42935 7395
rect 43269 7361 43303 7395
rect 44189 7361 44223 7395
rect 46029 7361 46063 7395
rect 48237 7361 48271 7395
rect 49157 7361 49191 7395
rect 49985 7361 50019 7395
rect 51733 7361 51767 7395
rect 54769 7361 54803 7395
rect 56333 7361 56367 7395
rect 57529 7361 57563 7395
rect 4997 7293 5031 7327
rect 5089 7293 5123 7327
rect 7205 7293 7239 7327
rect 8125 7293 8159 7327
rect 8217 7293 8251 7327
rect 9229 7293 9263 7327
rect 10793 7293 10827 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 18889 7293 18923 7327
rect 19257 7293 19291 7327
rect 24317 7293 24351 7327
rect 27537 7293 27571 7327
rect 28365 7293 28399 7327
rect 29009 7293 29043 7327
rect 31033 7293 31067 7327
rect 31125 7293 31159 7327
rect 33425 7293 33459 7327
rect 36093 7293 36127 7327
rect 37565 7293 37599 7327
rect 40141 7293 40175 7327
rect 40509 7293 40543 7327
rect 41613 7293 41647 7327
rect 42993 7293 43027 7327
rect 43821 7293 43855 7327
rect 55229 7293 55263 7327
rect 58449 7293 58483 7327
rect 2881 7225 2915 7259
rect 4537 7225 4571 7259
rect 8401 7225 8435 7259
rect 8769 7225 8803 7259
rect 13369 7225 13403 7259
rect 23581 7225 23615 7259
rect 26617 7225 26651 7259
rect 56977 7225 57011 7259
rect 2605 7157 2639 7191
rect 2789 7157 2823 7191
rect 7021 7157 7055 7191
rect 7757 7157 7791 7191
rect 8309 7157 8343 7191
rect 8999 7157 9033 7191
rect 11345 7157 11379 7191
rect 14933 7157 14967 7191
rect 16865 7157 16899 7191
rect 18153 7157 18187 7191
rect 18337 7157 18371 7191
rect 19901 7157 19935 7191
rect 21557 7157 21591 7191
rect 22017 7157 22051 7191
rect 23765 7157 23799 7191
rect 26985 7157 27019 7191
rect 27905 7157 27939 7191
rect 29561 7157 29595 7191
rect 30389 7157 30423 7191
rect 30573 7157 30607 7191
rect 36461 7157 36495 7191
rect 38669 7157 38703 7191
rect 39037 7157 39071 7191
rect 44649 7157 44683 7191
rect 45293 7157 45327 7191
rect 45661 7157 45695 7191
rect 46489 7157 46523 7191
rect 52009 7157 52043 7191
rect 52561 7157 52595 7191
rect 52929 7157 52963 7191
rect 55505 7157 55539 7191
rect 4537 6953 4571 6987
rect 14105 6953 14139 6987
rect 23489 6953 23523 6987
rect 26341 6953 26375 6987
rect 45477 6953 45511 6987
rect 55597 6953 55631 6987
rect 5457 6885 5491 6919
rect 21373 6885 21407 6919
rect 34989 6885 35023 6919
rect 36921 6885 36955 6919
rect 44005 6885 44039 6919
rect 44373 6885 44407 6919
rect 45293 6885 45327 6919
rect 53481 6885 53515 6919
rect 3341 6817 3375 6851
rect 4353 6817 4387 6851
rect 5641 6817 5675 6851
rect 7389 6817 7423 6851
rect 7941 6817 7975 6851
rect 8125 6817 8159 6851
rect 18889 6817 18923 6851
rect 19257 6817 19291 6851
rect 19901 6817 19935 6851
rect 20177 6817 20211 6851
rect 20294 6817 20328 6851
rect 22017 6817 22051 6851
rect 23949 6817 23983 6851
rect 24133 6817 24167 6851
rect 25329 6817 25363 6851
rect 25605 6817 25639 6851
rect 26249 6817 26283 6851
rect 26801 6817 26835 6851
rect 26893 6817 26927 6851
rect 27813 6817 27847 6851
rect 30021 6817 30055 6851
rect 30113 6817 30147 6851
rect 30481 6817 30515 6851
rect 31033 6817 31067 6851
rect 33885 6817 33919 6851
rect 36277 6817 36311 6851
rect 37565 6817 37599 6851
rect 40417 6817 40451 6851
rect 42211 6817 42245 6851
rect 42349 6817 42383 6851
rect 42625 6817 42659 6851
rect 43269 6817 43303 6851
rect 46673 6817 46707 6851
rect 47409 6817 47443 6851
rect 51825 6817 51859 6851
rect 52745 6817 52779 6851
rect 54217 6817 54251 6851
rect 56241 6817 56275 6851
rect 56793 6817 56827 6851
rect 4721 6749 4755 6783
rect 4997 6749 5031 6783
rect 6837 6749 6871 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 10333 6749 10367 6783
rect 12357 6749 12391 6783
rect 12613 6749 12647 6783
rect 14657 6749 14691 6783
rect 15393 6749 15427 6783
rect 16221 6749 16255 6783
rect 16865 6749 16899 6783
rect 19441 6749 19475 6783
rect 20453 6749 20487 6783
rect 21925 6749 21959 6783
rect 25053 6749 25087 6783
rect 25191 6749 25225 6783
rect 26065 6749 26099 6783
rect 28549 6749 28583 6783
rect 29377 6749 29411 6783
rect 31769 6749 31803 6783
rect 33517 6749 33551 6783
rect 36001 6749 36035 6783
rect 36461 6749 36495 6783
rect 37013 6749 37047 6783
rect 39681 6749 39715 6783
rect 40325 6749 40359 6783
rect 41245 6749 41279 6783
rect 42073 6749 42107 6783
rect 43085 6749 43119 6783
rect 46305 6749 46339 6783
rect 47041 6749 47075 6783
rect 51917 6749 51951 6783
rect 53021 6749 53055 6783
rect 54033 6749 54067 6783
rect 54769 6749 54803 6783
rect 57069 6749 57103 6783
rect 58081 6749 58115 6783
rect 58541 6749 58575 6783
rect 3096 6681 3130 6715
rect 3801 6681 3835 6715
rect 5181 6681 5215 6715
rect 8585 6681 8619 6715
rect 10600 6681 10634 6715
rect 12265 6681 12299 6715
rect 17132 6681 17166 6715
rect 18705 6681 18739 6715
rect 22284 6681 22318 6715
rect 26709 6681 26743 6715
rect 27537 6681 27571 6715
rect 27997 6681 28031 6715
rect 29929 6681 29963 6715
rect 31217 6681 31251 6715
rect 33272 6681 33306 6715
rect 33701 6681 33735 6715
rect 34253 6681 34287 6715
rect 35357 6681 35391 6715
rect 37933 6681 37967 6715
rect 38669 6681 38703 6715
rect 40233 6681 40267 6715
rect 40693 6681 40727 6715
rect 45569 6681 45603 6715
rect 56057 6681 56091 6715
rect 1961 6613 1995 6647
rect 4905 6613 4939 6647
rect 6009 6613 6043 6647
rect 6653 6613 6687 6647
rect 7481 6613 7515 6647
rect 7849 6613 7883 6647
rect 10241 6613 10275 6647
rect 11713 6613 11747 6647
rect 13737 6613 13771 6647
rect 14841 6613 14875 6647
rect 15853 6613 15887 6647
rect 16773 6613 16807 6647
rect 18245 6613 18279 6647
rect 18337 6613 18371 6647
rect 18797 6613 18831 6647
rect 21097 6613 21131 6647
rect 23397 6613 23431 6647
rect 23857 6613 23891 6647
rect 24409 6613 24443 6647
rect 27169 6613 27203 6647
rect 27629 6613 27663 6647
rect 28733 6613 28767 6647
rect 29561 6613 29595 6647
rect 32137 6613 32171 6647
rect 35449 6613 35483 6647
rect 36553 6613 36587 6647
rect 38393 6613 38427 6647
rect 39037 6613 39071 6647
rect 39865 6613 39899 6647
rect 41429 6613 41463 6647
rect 43637 6613 43671 6647
rect 44741 6613 44775 6647
rect 45753 6613 45787 6647
rect 47777 6613 47811 6647
rect 48145 6613 48179 6647
rect 48973 6613 49007 6647
rect 50353 6613 50387 6647
rect 50905 6613 50939 6647
rect 51273 6613 51307 6647
rect 52561 6613 52595 6647
rect 52929 6613 52963 6647
rect 53389 6613 53423 6647
rect 55689 6613 55723 6647
rect 56149 6613 56183 6647
rect 56977 6613 57011 6647
rect 57437 6613 57471 6647
rect 57529 6613 57563 6647
rect 58357 6613 58391 6647
rect 6929 6409 6963 6443
rect 9873 6409 9907 6443
rect 11529 6409 11563 6443
rect 12449 6409 12483 6443
rect 14381 6409 14415 6443
rect 18153 6409 18187 6443
rect 18521 6409 18555 6443
rect 18981 6409 19015 6443
rect 19717 6409 19751 6443
rect 25237 6409 25271 6443
rect 29929 6409 29963 6443
rect 40233 6409 40267 6443
rect 43821 6409 43855 6443
rect 48789 6409 48823 6443
rect 51641 6409 51675 6443
rect 51825 6409 51859 6443
rect 52193 6409 52227 6443
rect 54125 6409 54159 6443
rect 6009 6341 6043 6375
rect 8134 6341 8168 6375
rect 10232 6341 10266 6375
rect 15516 6341 15550 6375
rect 15853 6341 15887 6375
rect 16926 6341 16960 6375
rect 18613 6341 18647 6375
rect 23121 6341 23155 6375
rect 26372 6341 26406 6375
rect 26985 6341 27019 6375
rect 34897 6341 34931 6375
rect 35440 6341 35474 6375
rect 38669 6341 38703 6375
rect 42257 6341 42291 6375
rect 42686 6341 42720 6375
rect 45376 6341 45410 6375
rect 49249 6341 49283 6375
rect 50537 6341 50571 6375
rect 53012 6341 53046 6375
rect 5365 6273 5399 6307
rect 8401 6273 8435 6307
rect 9505 6273 9539 6307
rect 9965 6273 9999 6307
rect 11897 6273 11931 6307
rect 13093 6273 13127 6307
rect 14289 6273 14323 6307
rect 16681 6273 16715 6307
rect 19625 6273 19659 6307
rect 20830 6273 20864 6307
rect 21097 6273 21131 6307
rect 22385 6273 22419 6307
rect 23029 6273 23063 6307
rect 23489 6273 23523 6307
rect 24133 6273 24167 6307
rect 24777 6273 24811 6307
rect 24961 6273 24995 6307
rect 27537 6273 27571 6307
rect 28805 6273 28839 6307
rect 31134 6273 31168 6307
rect 33250 6273 33284 6307
rect 33609 6273 33643 6307
rect 35173 6273 35207 6307
rect 36921 6273 36955 6307
rect 37841 6273 37875 6307
rect 39109 6273 39143 6307
rect 44465 6273 44499 6307
rect 45109 6273 45143 6307
rect 49341 6273 49375 6307
rect 52285 6273 52319 6307
rect 52745 6273 52779 6307
rect 54953 6273 54987 6307
rect 57457 6273 57491 6307
rect 57713 6273 57747 6307
rect 3341 6205 3375 6239
rect 4077 6205 4111 6239
rect 4997 6205 5031 6239
rect 9137 6205 9171 6239
rect 11989 6205 12023 6239
rect 12173 6205 12207 6239
rect 13231 6205 13265 6239
rect 13369 6205 13403 6239
rect 14105 6205 14139 6239
rect 15761 6205 15795 6239
rect 16405 6205 16439 6239
rect 18705 6205 18739 6239
rect 23213 6205 23247 6239
rect 26617 6205 26651 6239
rect 28549 6205 28583 6239
rect 31401 6205 31435 6239
rect 33517 6205 33551 6239
rect 34437 6205 34471 6239
rect 38853 6205 38887 6239
rect 40877 6205 40911 6239
rect 41705 6205 41739 6239
rect 42441 6205 42475 6239
rect 47133 6205 47167 6239
rect 49065 6205 49099 6239
rect 50353 6205 50387 6239
rect 51089 6205 51123 6239
rect 52377 6205 52411 6239
rect 55091 6205 55125 6239
rect 55229 6205 55263 6239
rect 55505 6205 55539 6239
rect 55965 6205 55999 6239
rect 56149 6205 56183 6239
rect 57897 6205 57931 6239
rect 58449 6205 58483 6239
rect 2329 6137 2363 6171
rect 11345 6137 11379 6171
rect 13645 6137 13679 6171
rect 18061 6137 18095 6171
rect 21649 6137 21683 6171
rect 24501 6137 24535 6171
rect 38209 6137 38243 6171
rect 46489 6137 46523 6171
rect 49709 6137 49743 6171
rect 2697 6069 2731 6103
rect 2789 6069 2823 6103
rect 3525 6069 3559 6103
rect 4445 6069 4479 6103
rect 7021 6069 7055 6103
rect 21833 6069 21867 6103
rect 22661 6069 22695 6103
rect 27905 6069 27939 6103
rect 28365 6069 28399 6103
rect 30021 6069 30055 6103
rect 31861 6069 31895 6103
rect 32137 6069 32171 6103
rect 36553 6069 36587 6103
rect 37289 6069 37323 6103
rect 40325 6069 40359 6103
rect 41245 6069 41279 6103
rect 43913 6069 43947 6103
rect 44833 6069 44867 6103
rect 46581 6069 46615 6103
rect 47777 6069 47811 6103
rect 48513 6069 48547 6103
rect 49801 6069 49835 6103
rect 54309 6069 54343 6103
rect 56333 6069 56367 6103
rect 3525 5865 3559 5899
rect 4261 5865 4295 5899
rect 6101 5865 6135 5899
rect 10701 5865 10735 5899
rect 11529 5865 11563 5899
rect 15209 5865 15243 5899
rect 17785 5865 17819 5899
rect 20913 5865 20947 5899
rect 22293 5865 22327 5899
rect 22477 5865 22511 5899
rect 28457 5865 28491 5899
rect 33701 5865 33735 5899
rect 38025 5865 38059 5899
rect 38485 5865 38519 5899
rect 38761 5865 38795 5899
rect 41153 5865 41187 5899
rect 42349 5865 42383 5899
rect 43729 5865 43763 5899
rect 46581 5865 46615 5899
rect 48605 5865 48639 5899
rect 53113 5865 53147 5899
rect 56701 5865 56735 5899
rect 56793 5865 56827 5899
rect 58449 5865 58483 5899
rect 5733 5797 5767 5831
rect 10609 5797 10643 5831
rect 13737 5797 13771 5831
rect 17233 5797 17267 5831
rect 18981 5797 19015 5831
rect 24685 5797 24719 5831
rect 25605 5797 25639 5831
rect 32137 5797 32171 5831
rect 35633 5797 35667 5831
rect 47869 5797 47903 5831
rect 50905 5797 50939 5831
rect 7113 5729 7147 5763
rect 7389 5729 7423 5763
rect 8033 5729 8067 5763
rect 9321 5729 9355 5763
rect 11253 5729 11287 5763
rect 12081 5729 12115 5763
rect 13185 5729 13219 5763
rect 14657 5729 14691 5763
rect 17601 5729 17635 5763
rect 18337 5729 18371 5763
rect 20177 5729 20211 5763
rect 23029 5729 23063 5763
rect 24961 5729 24995 5763
rect 26157 5729 26191 5763
rect 28825 5729 28859 5763
rect 31861 5729 31895 5763
rect 32597 5729 32631 5763
rect 33057 5729 33091 5763
rect 35265 5729 35299 5763
rect 39497 5729 39531 5763
rect 42993 5729 43027 5763
rect 44465 5729 44499 5763
rect 45201 5729 45235 5763
rect 47455 5729 47489 5763
rect 47593 5729 47627 5763
rect 48513 5729 48547 5763
rect 50261 5729 50295 5763
rect 51549 5729 51583 5763
rect 1685 5661 1719 5695
rect 2053 5661 2087 5695
rect 2145 5661 2179 5695
rect 4353 5661 4387 5695
rect 4609 5661 4643 5695
rect 6837 5661 6871 5695
rect 6996 5661 7030 5695
rect 7849 5661 7883 5695
rect 8125 5661 8159 5695
rect 9965 5661 9999 5695
rect 12357 5661 12391 5695
rect 14841 5661 14875 5695
rect 19901 5661 19935 5695
rect 20453 5661 20487 5695
rect 21465 5661 21499 5695
rect 25513 5661 25547 5695
rect 25973 5661 26007 5695
rect 26985 5661 27019 5695
rect 27445 5661 27479 5695
rect 29561 5661 29595 5695
rect 30389 5661 30423 5695
rect 31585 5661 31619 5695
rect 31744 5661 31778 5695
rect 32781 5661 32815 5695
rect 34253 5661 34287 5695
rect 36757 5661 36791 5695
rect 37013 5661 37047 5695
rect 37657 5661 37691 5695
rect 39313 5661 39347 5695
rect 39865 5661 39899 5695
rect 42717 5661 42751 5695
rect 47317 5661 47351 5695
rect 48329 5661 48363 5695
rect 49718 5661 49752 5695
rect 49985 5661 50019 5695
rect 50997 5661 51031 5695
rect 51733 5661 51767 5695
rect 54953 5661 54987 5695
rect 55321 5661 55355 5695
rect 57345 5661 57379 5695
rect 58081 5661 58115 5695
rect 58265 5661 58299 5695
rect 2412 5593 2446 5627
rect 13369 5593 13403 5627
rect 15577 5593 15611 5627
rect 15945 5593 15979 5627
rect 16497 5593 16531 5627
rect 16865 5593 16899 5627
rect 22017 5593 22051 5627
rect 23489 5593 23523 5627
rect 28917 5593 28951 5627
rect 33149 5593 33183 5627
rect 34713 5593 34747 5627
rect 37933 5593 37967 5627
rect 39405 5593 39439 5627
rect 44189 5593 44223 5627
rect 45468 5593 45502 5627
rect 52000 5593 52034 5627
rect 53205 5593 53239 5627
rect 55588 5593 55622 5627
rect 6193 5525 6227 5559
rect 8769 5525 8803 5559
rect 11069 5525 11103 5559
rect 11161 5525 11195 5559
rect 12909 5525 12943 5559
rect 13277 5525 13311 5559
rect 14289 5525 14323 5559
rect 14749 5525 14783 5559
rect 19441 5525 19475 5559
rect 20361 5525 20395 5559
rect 20821 5525 20855 5559
rect 24225 5525 24259 5559
rect 26065 5525 26099 5559
rect 26433 5525 26467 5559
rect 27721 5525 27755 5559
rect 28181 5525 28215 5559
rect 29009 5525 29043 5559
rect 29377 5525 29411 5559
rect 30941 5525 30975 5559
rect 33241 5525 33275 5559
rect 33609 5525 33643 5559
rect 37105 5525 37139 5559
rect 38945 5525 38979 5559
rect 41981 5525 42015 5559
rect 42809 5525 42843 5559
rect 43453 5525 43487 5559
rect 46673 5525 46707 5559
rect 50445 5525 50479 5559
rect 50537 5525 50571 5559
rect 57529 5525 57563 5559
rect 4353 5321 4387 5355
rect 6101 5321 6135 5355
rect 7481 5321 7515 5355
rect 10701 5321 10735 5355
rect 14841 5321 14875 5355
rect 16129 5321 16163 5355
rect 20637 5321 20671 5355
rect 21557 5321 21591 5355
rect 26709 5321 26743 5355
rect 27997 5321 28031 5355
rect 29561 5321 29595 5355
rect 30941 5321 30975 5355
rect 31309 5321 31343 5355
rect 35265 5321 35299 5355
rect 35725 5321 35759 5355
rect 36093 5321 36127 5355
rect 36185 5321 36219 5355
rect 37657 5321 37691 5355
rect 42165 5321 42199 5355
rect 43545 5321 43579 5355
rect 43913 5321 43947 5355
rect 44649 5321 44683 5355
rect 45661 5321 45695 5355
rect 46029 5321 46063 5355
rect 51089 5321 51123 5355
rect 52745 5321 52779 5355
rect 54033 5321 54067 5355
rect 54953 5321 54987 5355
rect 55689 5321 55723 5355
rect 56885 5321 56919 5355
rect 57621 5321 57655 5355
rect 3433 5253 3467 5287
rect 4813 5253 4847 5287
rect 5273 5253 5307 5287
rect 8697 5253 8731 5287
rect 11897 5253 11931 5287
rect 13584 5253 13618 5287
rect 13921 5253 13955 5287
rect 20361 5253 20395 5287
rect 23029 5253 23063 5287
rect 29469 5253 29503 5287
rect 32781 5253 32815 5287
rect 33977 5253 34011 5287
rect 34897 5253 34931 5287
rect 36737 5253 36771 5287
rect 38853 5253 38887 5287
rect 39190 5253 39224 5287
rect 42809 5253 42843 5287
rect 50016 5253 50050 5287
rect 54309 5253 54343 5287
rect 55229 5253 55263 5287
rect 2237 5185 2271 5219
rect 5365 5185 5399 5219
rect 6377 5185 6411 5219
rect 7021 5185 7055 5219
rect 8953 5185 8987 5219
rect 9689 5185 9723 5219
rect 10057 5185 10091 5219
rect 10609 5185 10643 5219
rect 11805 5185 11839 5219
rect 14473 5185 14507 5219
rect 16497 5185 16531 5219
rect 18429 5185 18463 5219
rect 19533 5185 19567 5219
rect 20821 5185 20855 5219
rect 21281 5185 21315 5219
rect 23121 5185 23155 5219
rect 23489 5185 23523 5219
rect 24133 5185 24167 5219
rect 25329 5185 25363 5219
rect 25596 5185 25630 5219
rect 30297 5185 30331 5219
rect 32689 5185 32723 5219
rect 33241 5185 33275 5219
rect 33793 5185 33827 5219
rect 34529 5185 34563 5219
rect 38945 5185 38979 5219
rect 44189 5185 44223 5219
rect 46857 5185 46891 5219
rect 46949 5185 46983 5219
rect 47593 5185 47627 5219
rect 48145 5185 48179 5219
rect 50261 5185 50295 5219
rect 50537 5185 50571 5219
rect 50905 5185 50939 5219
rect 53389 5185 53423 5219
rect 53573 5185 53607 5219
rect 54493 5185 54527 5219
rect 55597 5185 55631 5219
rect 56241 5185 56275 5219
rect 56977 5185 57011 5219
rect 57437 5185 57471 5219
rect 3525 5117 3559 5151
rect 3617 5117 3651 5151
rect 5457 5117 5491 5151
rect 11345 5117 11379 5151
rect 11713 5117 11747 5151
rect 13829 5117 13863 5151
rect 17233 5117 17267 5151
rect 18061 5117 18095 5151
rect 19257 5117 19291 5151
rect 19717 5117 19751 5151
rect 19993 5117 20027 5151
rect 22569 5117 22603 5151
rect 23213 5117 23247 5151
rect 24777 5117 24811 5151
rect 27169 5117 27203 5151
rect 27537 5117 27571 5151
rect 30205 5117 30239 5151
rect 31677 5117 31711 5151
rect 32597 5117 32631 5151
rect 36277 5117 36311 5151
rect 37749 5117 37783 5151
rect 37933 5117 37967 5151
rect 38301 5117 38335 5151
rect 41061 5117 41095 5151
rect 42533 5117 42567 5151
rect 42717 5117 42751 5151
rect 46121 5117 46155 5151
rect 46213 5117 46247 5151
rect 47133 5117 47167 5151
rect 50721 5117 50755 5151
rect 51641 5117 51675 5151
rect 56701 5117 56735 5151
rect 58449 5117 58483 5151
rect 1869 5049 1903 5083
rect 3065 5049 3099 5083
rect 15761 5049 15795 5083
rect 22661 5049 22695 5083
rect 28641 5049 28675 5083
rect 29101 5049 29135 5083
rect 33149 5049 33183 5083
rect 40325 5049 40359 5083
rect 41429 5049 41463 5083
rect 45293 5049 45327 5083
rect 48513 5049 48547 5083
rect 57345 5049 57379 5083
rect 2605 4981 2639 5015
rect 2881 4981 2915 5015
rect 4905 4981 4939 5015
rect 7573 4981 7607 5015
rect 9045 4981 9079 5015
rect 12265 4981 12299 5015
rect 12449 4981 12483 5015
rect 15393 4981 15427 5015
rect 16681 4981 16715 5015
rect 17509 4981 17543 5015
rect 18613 4981 18647 5015
rect 19349 4981 19383 5015
rect 20269 4981 20303 5015
rect 21925 4981 21959 5015
rect 24225 4981 24259 5015
rect 25237 4981 25271 5015
rect 28365 4981 28399 5015
rect 37289 4981 37323 5015
rect 40417 4981 40451 5015
rect 41797 4981 41831 5015
rect 43177 4981 43211 5015
rect 44925 4981 44959 5015
rect 46489 4981 46523 5015
rect 48881 4981 48915 5015
rect 52009 4981 52043 5015
rect 52469 4981 52503 5015
rect 53757 4981 53791 5015
rect 55137 4981 55171 5015
rect 55413 4981 55447 5015
rect 57897 4981 57931 5015
rect 1777 4777 1811 4811
rect 6377 4777 6411 4811
rect 7205 4777 7239 4811
rect 9321 4777 9355 4811
rect 9965 4777 9999 4811
rect 16037 4777 16071 4811
rect 19257 4777 19291 4811
rect 21833 4777 21867 4811
rect 23397 4777 23431 4811
rect 26433 4777 26467 4811
rect 27629 4777 27663 4811
rect 35081 4777 35115 4811
rect 35541 4777 35575 4811
rect 37657 4777 37691 4811
rect 38025 4777 38059 4811
rect 38853 4777 38887 4811
rect 39589 4777 39623 4811
rect 42441 4777 42475 4811
rect 46029 4777 46063 4811
rect 48789 4777 48823 4811
rect 51733 4777 51767 4811
rect 55137 4777 55171 4811
rect 6009 4709 6043 4743
rect 6745 4709 6779 4743
rect 9597 4709 9631 4743
rect 14841 4709 14875 4743
rect 17509 4709 17543 4743
rect 25605 4709 25639 4743
rect 31033 4709 31067 4743
rect 36461 4709 36495 4743
rect 41245 4709 41279 4743
rect 47685 4709 47719 4743
rect 49157 4709 49191 4743
rect 49525 4709 49559 4743
rect 56517 4709 56551 4743
rect 7757 4641 7791 4675
rect 8677 4641 8711 4675
rect 14289 4641 14323 4675
rect 19901 4641 19935 4675
rect 22017 4641 22051 4675
rect 24041 4641 24075 4675
rect 25191 4641 25225 4675
rect 25329 4641 25363 4675
rect 26249 4641 26283 4675
rect 29377 4641 29411 4675
rect 33333 4641 33367 4675
rect 34437 4641 34471 4675
rect 35817 4641 35851 4675
rect 36737 4641 36771 4675
rect 37013 4641 37047 4675
rect 40601 4641 40635 4675
rect 41521 4641 41555 4675
rect 41659 4641 41693 4675
rect 43913 4641 43947 4675
rect 46581 4641 46615 4675
rect 48053 4641 48087 4675
rect 48421 4641 48455 4675
rect 53297 4641 53331 4675
rect 55321 4641 55355 4675
rect 57897 4641 57931 4675
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 4905 4573 4939 4607
rect 5733 4573 5767 4607
rect 6561 4573 6595 4607
rect 7573 4573 7607 4607
rect 8401 4573 8435 4607
rect 11529 4573 11563 4607
rect 11621 4573 11655 4607
rect 13369 4573 13403 4607
rect 13461 4573 13495 4607
rect 14473 4573 14507 4607
rect 16129 4573 16163 4607
rect 17693 4573 17727 4607
rect 17960 4573 17994 4607
rect 20729 4573 20763 4607
rect 20821 4573 20855 4607
rect 22273 4573 22307 4607
rect 23857 4573 23891 4607
rect 25053 4573 25087 4607
rect 26065 4573 26099 4607
rect 26617 4573 26651 4607
rect 26709 4573 26743 4607
rect 27261 4573 27295 4607
rect 27997 4573 28031 4607
rect 28273 4573 28307 4607
rect 28365 4573 28399 4607
rect 28825 4573 28859 4607
rect 29561 4573 29595 4607
rect 32505 4573 32539 4607
rect 33149 4573 33183 4607
rect 33885 4573 33919 4607
rect 35357 4573 35391 4607
rect 36001 4573 36035 4607
rect 36854 4573 36888 4607
rect 39037 4573 39071 4607
rect 39405 4573 39439 4607
rect 40417 4573 40451 4607
rect 40785 4573 40819 4607
rect 41797 4573 41831 4607
rect 44649 4573 44683 4607
rect 45201 4573 45235 4607
rect 45937 4573 45971 4607
rect 47317 4573 47351 4607
rect 47501 4573 47535 4607
rect 48973 4573 49007 4607
rect 50169 4573 50203 4607
rect 51457 4573 51491 4607
rect 51917 4573 51951 4607
rect 52101 4573 52135 4607
rect 53113 4573 53147 4607
rect 54125 4573 54159 4607
rect 54585 4573 54619 4607
rect 55505 4573 55539 4607
rect 55689 4573 55723 4607
rect 55781 4573 55815 4607
rect 57641 4573 57675 4607
rect 58173 4573 58207 4607
rect 58265 4573 58299 4607
rect 2145 4505 2179 4539
rect 11284 4505 11318 4539
rect 15209 4505 15243 4539
rect 15485 4505 15519 4539
rect 16396 4505 16430 4539
rect 19625 4505 19659 4539
rect 28549 4505 28583 4539
rect 30389 4505 30423 4539
rect 32260 4505 32294 4539
rect 34161 4505 34195 4539
rect 35173 4505 35207 4539
rect 38669 4505 38703 4539
rect 43668 4505 43702 4539
rect 44005 4505 44039 4539
rect 49893 4505 49927 4539
rect 2237 4437 2271 4471
rect 3617 4437 3651 4471
rect 4261 4437 4295 4471
rect 4353 4437 4387 4471
rect 5089 4437 5123 4471
rect 7389 4437 7423 4471
rect 8033 4437 8067 4471
rect 8493 4437 8527 4471
rect 10149 4437 10183 4471
rect 13645 4437 13679 4471
rect 14381 4437 14415 4471
rect 15393 4437 15427 4471
rect 19073 4437 19107 4471
rect 19717 4437 19751 4471
rect 20085 4437 20119 4471
rect 21465 4437 21499 4471
rect 23489 4437 23523 4471
rect 23949 4437 23983 4471
rect 24409 4437 24443 4471
rect 26893 4437 26927 4471
rect 28641 4437 28675 4471
rect 31125 4437 31159 4471
rect 32597 4437 32631 4471
rect 38301 4437 38335 4471
rect 39865 4437 39899 4471
rect 42533 4437 42567 4471
rect 45017 4437 45051 4471
rect 45293 4437 45327 4471
rect 46765 4437 46799 4471
rect 49801 4437 49835 4471
rect 50813 4437 50847 4471
rect 50905 4437 50939 4471
rect 52653 4437 52687 4471
rect 52745 4437 52779 4471
rect 53205 4437 53239 4471
rect 53573 4437 53607 4471
rect 56425 4437 56459 4471
rect 57989 4437 58023 4471
rect 3249 4233 3283 4267
rect 3709 4233 3743 4267
rect 4353 4233 4387 4267
rect 4813 4233 4847 4267
rect 7481 4233 7515 4267
rect 7573 4233 7607 4267
rect 7941 4233 7975 4267
rect 9873 4233 9907 4267
rect 10149 4233 10183 4267
rect 11529 4233 11563 4267
rect 14105 4233 14139 4267
rect 16405 4233 16439 4267
rect 16957 4233 16991 4267
rect 17325 4233 17359 4267
rect 17417 4233 17451 4267
rect 20637 4233 20671 4267
rect 23397 4233 23431 4267
rect 24777 4233 24811 4267
rect 29837 4233 29871 4267
rect 32413 4233 32447 4267
rect 33333 4233 33367 4267
rect 40049 4233 40083 4267
rect 40509 4233 40543 4267
rect 42809 4233 42843 4267
rect 43269 4233 43303 4267
rect 46121 4233 46155 4267
rect 46581 4233 46615 4267
rect 47961 4233 47995 4267
rect 49065 4233 49099 4267
rect 50813 4233 50847 4267
rect 51273 4233 51307 4267
rect 56057 4233 56091 4267
rect 57253 4233 57287 4267
rect 2044 4165 2078 4199
rect 4721 4165 4755 4199
rect 8033 4165 8067 4199
rect 8769 4165 8803 4199
rect 10609 4165 10643 4199
rect 20545 4165 20579 4199
rect 27353 4165 27387 4199
rect 35633 4165 35667 4199
rect 36093 4165 36127 4199
rect 38844 4165 38878 4199
rect 41245 4165 41279 4199
rect 41429 4165 41463 4199
rect 44916 4165 44950 4199
rect 48881 4165 48915 4199
rect 50200 4165 50234 4199
rect 53113 4165 53147 4199
rect 57161 4165 57195 4199
rect 1777 4097 1811 4131
rect 3617 4097 3651 4131
rect 4077 4097 4111 4131
rect 6101 4097 6135 4131
rect 6561 4097 6595 4131
rect 6929 4097 6963 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 9413 4097 9447 4131
rect 9689 4097 9723 4131
rect 10885 4097 10919 4131
rect 12265 4097 12299 4131
rect 13461 4097 13495 4131
rect 15117 4097 15151 4131
rect 17969 4097 18003 4131
rect 18981 4097 19015 4131
rect 19257 4097 19291 4131
rect 19993 4097 20027 4131
rect 21649 4097 21683 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 25605 4097 25639 4131
rect 26065 4097 26099 4131
rect 27261 4097 27295 4131
rect 27629 4097 27663 4131
rect 27997 4097 28031 4131
rect 28264 4097 28298 4131
rect 29469 4097 29503 4131
rect 30021 4097 30055 4131
rect 30757 4097 30791 4131
rect 32505 4097 32539 4131
rect 33241 4097 33275 4131
rect 33793 4097 33827 4131
rect 33977 4097 34011 4131
rect 35725 4097 35759 4131
rect 37105 4097 37139 4131
rect 38209 4097 38243 4131
rect 38577 4097 38611 4131
rect 40417 4097 40451 4131
rect 41797 4097 41831 4131
rect 42073 4097 42107 4131
rect 43821 4097 43855 4131
rect 44281 4097 44315 4131
rect 44373 4097 44407 4131
rect 44649 4097 44683 4131
rect 46489 4097 46523 4131
rect 47225 4097 47259 4131
rect 48605 4097 48639 4131
rect 50445 4097 50479 4131
rect 50905 4097 50939 4131
rect 51641 4097 51675 4131
rect 52561 4097 52595 4131
rect 53849 4097 53883 4131
rect 54769 4097 54803 4131
rect 55965 4097 55999 4131
rect 56425 4097 56459 4131
rect 3801 4029 3835 4063
rect 4997 4029 5031 4063
rect 5825 4029 5859 4063
rect 6745 4029 6779 4063
rect 7113 4029 7147 4063
rect 7389 4029 7423 4063
rect 12173 4029 12207 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 13185 4029 13219 4063
rect 13323 4029 13357 4063
rect 14749 4029 14783 4063
rect 15301 4029 15335 4063
rect 17509 4029 17543 4063
rect 19119 4029 19153 4063
rect 20177 4029 20211 4063
rect 20453 4029 20487 4063
rect 21281 4029 21315 4063
rect 23765 4029 23799 4063
rect 24869 4029 24903 4063
rect 24961 4029 24995 4063
rect 25697 4029 25731 4063
rect 25789 4029 25823 4063
rect 26617 4029 26651 4063
rect 27445 4029 27479 4063
rect 30113 4029 30147 4063
rect 30895 4029 30929 4063
rect 31033 4029 31067 4063
rect 31309 4029 31343 4063
rect 31769 4029 31803 4063
rect 31953 4029 31987 4063
rect 32321 4029 32355 4063
rect 33149 4029 33183 4063
rect 34161 4029 34195 4063
rect 35173 4029 35207 4063
rect 35817 4029 35851 4063
rect 36645 4029 36679 4063
rect 37841 4029 37875 4063
rect 40601 4029 40635 4063
rect 41061 4029 41095 4063
rect 41981 4029 42015 4063
rect 42625 4029 42659 4063
rect 42717 4029 42751 4063
rect 46673 4029 46707 4063
rect 47685 4029 47719 4063
rect 47869 4029 47903 4063
rect 48789 4029 48823 4063
rect 50721 4029 50755 4063
rect 51457 4029 51491 4063
rect 51825 4029 51859 4063
rect 52929 4029 52963 4063
rect 53021 4029 53055 4063
rect 53665 4029 53699 4063
rect 54907 4029 54941 4063
rect 55045 4029 55079 4063
rect 55321 4029 55355 4063
rect 55781 4029 55815 4063
rect 56517 4029 56551 4063
rect 56701 4029 56735 4063
rect 57069 4029 57103 4063
rect 58449 4029 58483 4063
rect 3157 3961 3191 3995
rect 8217 3961 8251 3995
rect 15669 3961 15703 3995
rect 19533 3961 19567 3995
rect 21005 3961 21039 3995
rect 25237 3961 25271 3995
rect 29653 3961 29687 3995
rect 32873 3961 32907 3995
rect 35265 3961 35299 3995
rect 38025 3961 38059 3995
rect 39957 3961 39991 3995
rect 43177 3961 43211 3995
rect 46029 3961 46063 3995
rect 48421 3961 48455 3995
rect 53481 3961 53515 3995
rect 57621 3961 57655 3995
rect 1685 3893 1719 3927
rect 4261 3893 4295 3927
rect 6469 3893 6503 3927
rect 8033 3893 8067 3927
rect 11253 3893 11287 3927
rect 14197 3893 14231 3927
rect 14933 3893 14967 3927
rect 16037 3893 16071 3927
rect 18153 3893 18187 3927
rect 18337 3893 18371 3927
rect 21465 3893 21499 3927
rect 24317 3893 24351 3927
rect 24409 3893 24443 3927
rect 27077 3893 27111 3927
rect 27353 3893 27387 3927
rect 27813 3893 27847 3927
rect 29377 3893 29411 3927
rect 33701 3893 33735 3927
rect 34529 3893 34563 3927
rect 36921 3893 36955 3927
rect 37289 3893 37323 3927
rect 41613 3893 41647 3927
rect 42257 3893 42291 3927
rect 44557 3893 44591 3927
rect 47041 3893 47075 3927
rect 48329 3893 48363 3927
rect 48697 3893 48731 3927
rect 51917 3893 51951 3927
rect 54033 3893 54067 3927
rect 54125 3893 54159 3927
rect 57897 3893 57931 3927
rect 3525 3689 3559 3723
rect 7849 3689 7883 3723
rect 10609 3689 10643 3723
rect 15669 3689 15703 3723
rect 16221 3689 16255 3723
rect 17417 3689 17451 3723
rect 22937 3689 22971 3723
rect 25973 3689 26007 3723
rect 26249 3689 26283 3723
rect 28733 3689 28767 3723
rect 36093 3689 36127 3723
rect 36185 3689 36219 3723
rect 37657 3689 37691 3723
rect 42901 3689 42935 3723
rect 46213 3689 46247 3723
rect 48329 3689 48363 3723
rect 51641 3689 51675 3723
rect 53573 3689 53607 3723
rect 54309 3689 54343 3723
rect 55413 3689 55447 3723
rect 1961 3621 1995 3655
rect 5365 3621 5399 3655
rect 6101 3621 6135 3655
rect 7021 3621 7055 3655
rect 7481 3621 7515 3655
rect 9689 3621 9723 3655
rect 15025 3621 15059 3655
rect 21465 3621 21499 3655
rect 27905 3621 27939 3655
rect 29561 3621 29595 3655
rect 40601 3621 40635 3655
rect 43453 3621 43487 3655
rect 45293 3621 45327 3655
rect 47409 3621 47443 3655
rect 49157 3621 49191 3655
rect 51825 3621 51859 3655
rect 53481 3621 53515 3655
rect 2145 3553 2179 3587
rect 2973 3553 3007 3587
rect 4813 3553 4847 3587
rect 4951 3553 4985 3587
rect 5070 3553 5104 3587
rect 5825 3553 5859 3587
rect 6653 3553 6687 3587
rect 8125 3553 8159 3587
rect 9045 3553 9079 3587
rect 9229 3553 9263 3587
rect 10333 3553 10367 3587
rect 12265 3553 12299 3587
rect 13277 3553 13311 3587
rect 16405 3553 16439 3587
rect 16865 3553 16899 3587
rect 19717 3553 19751 3587
rect 20821 3553 20855 3587
rect 22109 3553 22143 3587
rect 23489 3553 23523 3587
rect 23765 3553 23799 3587
rect 24593 3553 24627 3587
rect 26709 3553 26743 3587
rect 29377 3553 29411 3587
rect 30113 3553 30147 3587
rect 30941 3553 30975 3587
rect 32229 3553 32263 3587
rect 33517 3553 33551 3587
rect 33977 3553 34011 3587
rect 38117 3553 38151 3587
rect 38301 3553 38335 3587
rect 39037 3553 39071 3587
rect 39957 3553 39991 3587
rect 40141 3553 40175 3587
rect 41245 3553 41279 3587
rect 43085 3553 43119 3587
rect 43177 3553 43211 3587
rect 43729 3553 43763 3587
rect 44281 3553 44315 3587
rect 45845 3553 45879 3587
rect 46857 3553 46891 3587
rect 47133 3553 47167 3587
rect 48053 3553 48087 3587
rect 48513 3553 48547 3587
rect 49065 3553 49099 3587
rect 49709 3553 49743 3587
rect 54217 3553 54251 3587
rect 56609 3553 56643 3587
rect 57621 3553 57655 3587
rect 3065 3485 3099 3519
rect 6009 3485 6043 3519
rect 8033 3485 8067 3519
rect 10793 3485 10827 3519
rect 11529 3485 11563 3519
rect 13001 3485 13035 3519
rect 14657 3485 14691 3519
rect 14841 3485 14875 3519
rect 15301 3485 15335 3519
rect 15393 3485 15427 3519
rect 15853 3485 15887 3519
rect 16221 3485 16255 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 17601 3485 17635 3519
rect 18337 3485 18371 3519
rect 18981 3485 19015 3519
rect 19349 3485 19383 3519
rect 21005 3485 21039 3519
rect 21097 3485 21131 3519
rect 22293 3485 22327 3519
rect 22569 3485 22603 3519
rect 23949 3485 23983 3519
rect 26985 3485 27019 3519
rect 27169 3485 27203 3519
rect 27353 3485 27387 3519
rect 28089 3485 28123 3519
rect 31309 3485 31343 3519
rect 31953 3485 31987 3519
rect 32413 3485 32447 3519
rect 34069 3485 34103 3519
rect 34713 3485 34747 3519
rect 37565 3485 37599 3519
rect 39221 3485 39255 3519
rect 39405 3485 39439 3519
rect 41981 3485 42015 3519
rect 42165 3485 42199 3519
rect 42809 3485 42843 3519
rect 43637 3485 43671 3519
rect 43913 3485 43947 3519
rect 45201 3485 45235 3519
rect 45753 3485 45787 3519
rect 47016 3485 47050 3519
rect 47869 3485 47903 3519
rect 48145 3485 48179 3519
rect 50721 3485 50755 3519
rect 50997 3485 51031 3519
rect 52009 3485 52043 3519
rect 52101 3485 52135 3519
rect 54861 3485 54895 3519
rect 55597 3485 55631 3519
rect 57069 3485 57103 3519
rect 57161 3485 57195 3519
rect 2697 3417 2731 3451
rect 3157 3417 3191 3451
rect 3893 3417 3927 3451
rect 7297 3417 7331 3451
rect 8769 3417 8803 3451
rect 9321 3417 9355 3451
rect 16497 3417 16531 3451
rect 24838 3417 24872 3451
rect 26157 3417 26191 3451
rect 29929 3417 29963 3451
rect 32505 3417 32539 3451
rect 32965 3417 32999 3451
rect 34253 3417 34287 3451
rect 34958 3417 34992 3451
rect 37320 3417 37354 3451
rect 38025 3417 38059 3451
rect 38485 3417 38519 3451
rect 40233 3417 40267 3451
rect 41429 3417 41463 3451
rect 42901 3417 42935 3451
rect 43269 3417 43303 3451
rect 49525 3417 49559 3451
rect 50169 3417 50203 3451
rect 52346 3417 52380 3451
rect 3985 3349 4019 3383
rect 4169 3349 4203 3383
rect 9781 3349 9815 3383
rect 10885 3349 10919 3383
rect 11713 3349 11747 3383
rect 12449 3349 12483 3383
rect 13921 3349 13955 3383
rect 14105 3349 14139 3383
rect 15117 3349 15151 3383
rect 16037 3349 16071 3383
rect 16589 3349 16623 3383
rect 17233 3349 17267 3383
rect 17693 3349 17727 3383
rect 18429 3349 18463 3383
rect 21557 3349 21591 3383
rect 22477 3349 22511 3383
rect 22753 3349 22787 3383
rect 24133 3349 24167 3383
rect 26801 3349 26835 3383
rect 28641 3349 28675 3383
rect 30021 3349 30055 3383
rect 30389 3349 30423 3383
rect 31125 3349 31159 3383
rect 31401 3349 31435 3383
rect 32873 3349 32907 3383
rect 39589 3349 39623 3383
rect 40693 3349 40727 3383
rect 44097 3349 44131 3383
rect 44833 3349 44867 3383
rect 45017 3349 45051 3383
rect 45661 3349 45695 3383
rect 49617 3349 49651 3383
rect 1869 3145 1903 3179
rect 1961 3145 1995 3179
rect 5365 3145 5399 3179
rect 6653 3145 6687 3179
rect 7389 3145 7423 3179
rect 7573 3145 7607 3179
rect 7941 3145 7975 3179
rect 11345 3145 11379 3179
rect 11529 3145 11563 3179
rect 11897 3145 11931 3179
rect 11989 3145 12023 3179
rect 16405 3145 16439 3179
rect 18245 3145 18279 3179
rect 18337 3145 18371 3179
rect 18705 3145 18739 3179
rect 19901 3145 19935 3179
rect 20177 3145 20211 3179
rect 22937 3145 22971 3179
rect 23489 3145 23523 3179
rect 26801 3145 26835 3179
rect 27629 3145 27663 3179
rect 29101 3145 29135 3179
rect 32137 3145 32171 3179
rect 35081 3145 35115 3179
rect 36277 3145 36311 3179
rect 42441 3145 42475 3179
rect 43177 3145 43211 3179
rect 44373 3145 44407 3179
rect 47593 3145 47627 3179
rect 50169 3145 50203 3179
rect 54125 3145 54159 3179
rect 55965 3145 55999 3179
rect 57897 3145 57931 3179
rect 4252 3077 4286 3111
rect 6745 3077 6779 3111
rect 9076 3077 9110 3111
rect 10232 3077 10266 3111
rect 17132 3077 17166 3111
rect 19165 3077 19199 3111
rect 21312 3077 21346 3111
rect 27966 3077 28000 3111
rect 34989 3077 35023 3111
rect 39396 3077 39430 3111
rect 43637 3077 43671 3111
rect 44824 3077 44858 3111
rect 53012 3077 53046 3111
rect 57100 3077 57134 3111
rect 1685 3009 1719 3043
rect 3085 3009 3119 3043
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 3985 3009 4019 3043
rect 5457 3009 5491 3043
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 7113 3009 7147 3043
rect 7481 3009 7515 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 9597 3009 9631 3043
rect 9965 3009 9999 3043
rect 12541 3009 12575 3043
rect 13941 3009 13975 3043
rect 14197 3009 14231 3043
rect 15485 3009 15519 3043
rect 20085 3009 20119 3043
rect 21557 3009 21591 3043
rect 22109 3009 22143 3043
rect 22569 3009 22603 3043
rect 22661 3009 22695 3043
rect 23121 3009 23155 3043
rect 23397 3009 23431 3043
rect 24225 3009 24259 3043
rect 25881 3009 25915 3043
rect 27721 3009 27755 3043
rect 29193 3009 29227 3043
rect 31677 3009 31711 3043
rect 33261 3009 33295 3043
rect 33517 3009 33551 3043
rect 34161 3009 34195 3043
rect 35265 3009 35299 3043
rect 35541 3009 35575 3043
rect 35909 3009 35943 3043
rect 36093 3009 36127 3043
rect 36461 3009 36495 3043
rect 36737 3009 36771 3043
rect 36829 3009 36863 3043
rect 37013 3009 37047 3043
rect 37473 3009 37507 3043
rect 39129 3009 39163 3043
rect 41981 3009 42015 3043
rect 43361 3009 43395 3043
rect 43913 3009 43947 3043
rect 44097 3009 44131 3043
rect 44189 3009 44223 3043
rect 44557 3009 44591 3043
rect 46029 3009 46063 3043
rect 48237 3009 48271 3043
rect 48513 3009 48547 3043
rect 48789 3009 48823 3043
rect 49056 3009 49090 3043
rect 50445 3009 50479 3043
rect 50629 3009 50663 3043
rect 52101 3009 52135 3043
rect 52193 3009 52227 3043
rect 52377 3009 52411 3043
rect 52745 3009 52779 3043
rect 54217 3009 54251 3043
rect 55873 3009 55907 3043
rect 57345 3009 57379 3043
rect 57713 3009 57747 3043
rect 6009 2941 6043 2975
rect 12081 2941 12115 2975
rect 12725 2941 12759 2975
rect 14473 2941 14507 2975
rect 15761 2941 15795 2975
rect 16865 2941 16899 2975
rect 18797 2941 18831 2975
rect 18889 2941 18923 2975
rect 19717 2941 19751 2975
rect 21925 2941 21959 2975
rect 23305 2941 23339 2975
rect 24041 2941 24075 2975
rect 24685 2941 24719 2975
rect 25697 2941 25731 2975
rect 26249 2941 26283 2975
rect 27077 2941 27111 2975
rect 29653 2941 29687 2975
rect 30757 2941 30791 2975
rect 31861 2941 31895 2975
rect 33609 2941 33643 2975
rect 34345 2941 34379 2975
rect 35357 2941 35391 2975
rect 35725 2941 35759 2975
rect 37933 2941 37967 2975
rect 40969 2941 41003 2975
rect 42993 2941 43027 2975
rect 43545 2941 43579 2975
rect 46489 2941 46523 2975
rect 48697 2941 48731 2975
rect 50905 2941 50939 2975
rect 52561 2941 52595 2975
rect 54677 2941 54711 2975
rect 58449 2941 58483 2975
rect 7205 2873 7239 2907
rect 31401 2873 31435 2907
rect 3801 2805 3835 2839
rect 7757 2805 7791 2839
rect 9781 2805 9815 2839
rect 12357 2805 12391 2839
rect 12817 2805 12851 2839
rect 22293 2805 22327 2839
rect 22385 2805 22419 2839
rect 23121 2805 23155 2839
rect 26065 2805 26099 2839
rect 31493 2805 31527 2839
rect 35541 2805 35575 2839
rect 40509 2805 40543 2839
rect 43361 2805 43395 2839
rect 43729 2805 43763 2839
rect 45937 2805 45971 2839
rect 48329 2805 48363 2839
rect 50261 2805 50295 2839
rect 55689 2805 55723 2839
rect 57529 2805 57563 2839
rect 1961 2601 1995 2635
rect 9781 2601 9815 2635
rect 14105 2601 14139 2635
rect 17509 2601 17543 2635
rect 19441 2601 19475 2635
rect 21833 2601 21867 2635
rect 24041 2601 24075 2635
rect 25329 2601 25363 2635
rect 26985 2601 27019 2635
rect 27445 2601 27479 2635
rect 29561 2601 29595 2635
rect 32321 2601 32355 2635
rect 36921 2601 36955 2635
rect 38761 2601 38795 2635
rect 44557 2601 44591 2635
rect 46489 2601 46523 2635
rect 49801 2601 49835 2635
rect 51641 2601 51675 2635
rect 52377 2601 52411 2635
rect 54585 2601 54619 2635
rect 57161 2601 57195 2635
rect 57897 2601 57931 2635
rect 7297 2533 7331 2567
rect 13829 2533 13863 2567
rect 20177 2533 20211 2567
rect 24409 2533 24443 2567
rect 39497 2533 39531 2567
rect 42073 2533 42107 2567
rect 44649 2533 44683 2567
rect 54309 2533 54343 2567
rect 7849 2465 7883 2499
rect 10333 2465 10367 2499
rect 12541 2465 12575 2499
rect 14565 2465 14599 2499
rect 14657 2465 14691 2499
rect 15853 2465 15887 2499
rect 18061 2465 18095 2499
rect 23029 2465 23063 2499
rect 27997 2465 28031 2499
rect 30021 2465 30055 2499
rect 30113 2465 30147 2499
rect 34345 2465 34379 2499
rect 35173 2465 35207 2499
rect 40325 2465 40359 2499
rect 45569 2465 45603 2499
rect 47041 2465 47075 2499
rect 50629 2465 50663 2499
rect 53205 2465 53239 2499
rect 54953 2465 54987 2499
rect 56149 2465 56183 2499
rect 58449 2465 58483 2499
rect 3525 2397 3559 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 6193 2397 6227 2431
rect 6377 2397 6411 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 9229 2397 9263 2431
rect 9873 2397 9907 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13645 2397 13679 2431
rect 14473 2397 14507 2431
rect 15209 2397 15243 2431
rect 16957 2397 16991 2431
rect 17601 2397 17635 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 21649 2397 21683 2431
rect 22385 2397 22419 2431
rect 22569 2397 22603 2431
rect 24225 2397 24259 2431
rect 24593 2397 24627 2431
rect 24777 2397 24811 2431
rect 26801 2397 26835 2431
rect 27169 2397 27203 2431
rect 27261 2397 27295 2431
rect 27721 2397 27755 2431
rect 29101 2397 29135 2431
rect 29929 2397 29963 2431
rect 31769 2397 31803 2431
rect 32137 2397 32171 2431
rect 33885 2397 33919 2431
rect 33977 2397 34011 2431
rect 34161 2397 34195 2431
rect 34713 2397 34747 2431
rect 36737 2397 36771 2431
rect 37105 2397 37139 2431
rect 37473 2397 37507 2431
rect 38209 2397 38243 2431
rect 39313 2397 39347 2431
rect 39681 2397 39715 2431
rect 39865 2397 39899 2431
rect 41889 2397 41923 2431
rect 42257 2397 42291 2431
rect 43729 2397 43763 2431
rect 43913 2397 43947 2431
rect 44833 2397 44867 2431
rect 45017 2397 45051 2431
rect 48789 2397 48823 2431
rect 49065 2397 49099 2431
rect 49985 2397 50019 2431
rect 50261 2397 50295 2431
rect 52193 2397 52227 2431
rect 52561 2397 52595 2431
rect 52745 2397 52779 2431
rect 54493 2397 54527 2431
rect 54861 2397 54895 2431
rect 55597 2397 55631 2431
rect 55689 2397 55723 2431
rect 57345 2397 57379 2431
rect 57529 2397 57563 2431
rect 1685 2329 1719 2363
rect 2329 2329 2363 2363
rect 5273 2329 5307 2363
rect 20729 2329 20763 2363
rect 25789 2329 25823 2363
rect 26985 2329 27019 2363
rect 30757 2329 30791 2363
rect 32689 2329 32723 2363
rect 41337 2329 41371 2363
rect 42809 2329 42843 2363
rect 47777 2329 47811 2363
rect 6561 2261 6595 2295
rect 11713 2261 11747 2295
rect 29285 2261 29319 2295
rect 36185 2261 36219 2295
rect 49709 2261 49743 2295
rect 55413 2261 55447 2295
<< metal1 >>
rect 1104 21786 59040 21808
rect 1104 21734 15394 21786
rect 15446 21734 15458 21786
rect 15510 21734 15522 21786
rect 15574 21734 15586 21786
rect 15638 21734 15650 21786
rect 15702 21734 29838 21786
rect 29890 21734 29902 21786
rect 29954 21734 29966 21786
rect 30018 21734 30030 21786
rect 30082 21734 30094 21786
rect 30146 21734 44282 21786
rect 44334 21734 44346 21786
rect 44398 21734 44410 21786
rect 44462 21734 44474 21786
rect 44526 21734 44538 21786
rect 44590 21734 58726 21786
rect 58778 21734 58790 21786
rect 58842 21734 58854 21786
rect 58906 21734 58918 21786
rect 58970 21734 58982 21786
rect 59034 21734 59040 21786
rect 1104 21712 59040 21734
rect 37001 21539 37059 21545
rect 37001 21536 37013 21539
rect 32968 21508 37013 21536
rect 32968 21480 32996 21508
rect 37001 21505 37013 21508
rect 37047 21536 37059 21539
rect 38378 21536 38384 21548
rect 37047 21508 38384 21536
rect 37047 21505 37059 21508
rect 37001 21499 37059 21505
rect 38378 21496 38384 21508
rect 38436 21496 38442 21548
rect 5626 21428 5632 21480
rect 5684 21428 5690 21480
rect 9490 21428 9496 21480
rect 9548 21428 9554 21480
rect 12158 21428 12164 21480
rect 12216 21428 12222 21480
rect 12897 21471 12955 21477
rect 12897 21437 12909 21471
rect 12943 21468 12955 21471
rect 13446 21468 13452 21480
rect 12943 21440 13452 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 15381 21471 15439 21477
rect 15381 21468 15393 21471
rect 15252 21440 15393 21468
rect 15252 21428 15258 21440
rect 15381 21437 15393 21440
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 18598 21428 18604 21480
rect 18656 21428 18662 21480
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28350 21428 28356 21480
rect 28408 21468 28414 21480
rect 28629 21471 28687 21477
rect 28629 21468 28641 21471
rect 28408 21440 28641 21468
rect 28408 21428 28414 21440
rect 28629 21437 28641 21440
rect 28675 21437 28687 21471
rect 28629 21431 28687 21437
rect 30742 21428 30748 21480
rect 30800 21468 30806 21480
rect 31570 21468 31576 21480
rect 30800 21440 31576 21468
rect 30800 21428 30806 21440
rect 31570 21428 31576 21440
rect 31628 21428 31634 21480
rect 32950 21428 32956 21480
rect 33008 21428 33014 21480
rect 33410 21428 33416 21480
rect 33468 21428 33474 21480
rect 37829 21471 37887 21477
rect 37829 21468 37841 21471
rect 37660 21440 37841 21468
rect 37660 21412 37688 21440
rect 37829 21437 37841 21440
rect 37875 21437 37887 21471
rect 37829 21431 37887 21437
rect 38654 21428 38660 21480
rect 38712 21428 38718 21480
rect 39850 21428 39856 21480
rect 39908 21468 39914 21480
rect 40497 21471 40555 21477
rect 40497 21468 40509 21471
rect 39908 21440 40509 21468
rect 39908 21428 39914 21440
rect 40497 21437 40509 21440
rect 40543 21437 40555 21471
rect 40497 21431 40555 21437
rect 43254 21428 43260 21480
rect 43312 21428 43318 21480
rect 43990 21428 43996 21480
rect 44048 21428 44054 21480
rect 44082 21428 44088 21480
rect 44140 21468 44146 21480
rect 44177 21471 44235 21477
rect 44177 21468 44189 21471
rect 44140 21440 44189 21468
rect 44140 21428 44146 21440
rect 44177 21437 44189 21440
rect 44223 21437 44235 21471
rect 44177 21431 44235 21437
rect 46106 21428 46112 21480
rect 46164 21428 46170 21480
rect 48222 21428 48228 21480
rect 48280 21428 48286 21480
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 53374 21428 53380 21480
rect 53432 21428 53438 21480
rect 56594 21428 56600 21480
rect 56652 21428 56658 21480
rect 31662 21360 31668 21412
rect 31720 21400 31726 21412
rect 36357 21403 36415 21409
rect 36357 21400 36369 21403
rect 31720 21372 36369 21400
rect 31720 21360 31726 21372
rect 36357 21369 36369 21372
rect 36403 21400 36415 21403
rect 36906 21400 36912 21412
rect 36403 21372 36912 21400
rect 36403 21369 36415 21372
rect 36357 21363 36415 21369
rect 36906 21360 36912 21372
rect 36964 21360 36970 21412
rect 37277 21403 37335 21409
rect 37277 21369 37289 21403
rect 37323 21369 37335 21403
rect 37277 21363 37335 21369
rect 4982 21292 4988 21344
rect 5040 21292 5046 21344
rect 5166 21292 5172 21344
rect 5224 21332 5230 21344
rect 5905 21335 5963 21341
rect 5905 21332 5917 21335
rect 5224 21304 5917 21332
rect 5224 21292 5230 21304
rect 5905 21301 5917 21304
rect 5951 21301 5963 21335
rect 5905 21295 5963 21301
rect 8662 21292 8668 21344
rect 8720 21292 8726 21344
rect 8938 21292 8944 21344
rect 8996 21292 9002 21344
rect 11514 21292 11520 21344
rect 11572 21292 11578 21344
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 12253 21335 12311 21341
rect 12253 21332 12265 21335
rect 11664 21304 12265 21332
rect 11664 21292 11670 21304
rect 12253 21301 12265 21304
rect 12299 21301 12311 21335
rect 12253 21295 12311 21301
rect 14826 21292 14832 21344
rect 14884 21292 14890 21344
rect 18046 21292 18052 21344
rect 18104 21292 18110 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 22370 21332 22376 21344
rect 22143 21304 22376 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 24857 21335 24915 21341
rect 24857 21301 24869 21335
rect 24903 21332 24915 21335
rect 25590 21332 25596 21344
rect 24903 21304 25596 21332
rect 24903 21301 24915 21304
rect 24857 21295 24915 21301
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 27246 21292 27252 21344
rect 27304 21292 27310 21344
rect 28074 21292 28080 21344
rect 28132 21292 28138 21344
rect 30285 21335 30343 21341
rect 30285 21301 30297 21335
rect 30331 21332 30343 21335
rect 31294 21332 31300 21344
rect 30331 21304 31300 21332
rect 30331 21301 30343 21304
rect 30285 21295 30343 21301
rect 31294 21292 31300 21304
rect 31352 21292 31358 21344
rect 31386 21292 31392 21344
rect 31444 21292 31450 21344
rect 32401 21335 32459 21341
rect 32401 21301 32413 21335
rect 32447 21332 32459 21335
rect 32950 21332 32956 21344
rect 32447 21304 32956 21332
rect 32447 21301 32459 21304
rect 32401 21295 32459 21301
rect 32950 21292 32956 21304
rect 33008 21292 33014 21344
rect 33962 21292 33968 21344
rect 34020 21292 34026 21344
rect 34425 21335 34483 21341
rect 34425 21301 34437 21335
rect 34471 21332 34483 21335
rect 34514 21332 34520 21344
rect 34471 21304 34520 21332
rect 34471 21301 34483 21304
rect 34425 21295 34483 21301
rect 34514 21292 34520 21304
rect 34572 21292 34578 21344
rect 36722 21292 36728 21344
rect 36780 21332 36786 21344
rect 37292 21332 37320 21363
rect 37642 21360 37648 21412
rect 37700 21360 37706 21412
rect 46934 21360 46940 21412
rect 46992 21400 46998 21412
rect 47121 21403 47179 21409
rect 47121 21400 47133 21403
rect 46992 21372 47133 21400
rect 46992 21360 46998 21372
rect 47121 21369 47133 21372
rect 47167 21400 47179 21403
rect 51994 21400 52000 21412
rect 47167 21372 52000 21400
rect 47167 21369 47179 21372
rect 47121 21363 47179 21369
rect 51994 21360 52000 21372
rect 52052 21360 52058 21412
rect 36780 21304 37320 21332
rect 36780 21292 36786 21304
rect 38010 21292 38016 21344
rect 38068 21292 38074 21344
rect 39025 21335 39083 21341
rect 39025 21301 39037 21335
rect 39071 21332 39083 21335
rect 39206 21332 39212 21344
rect 39071 21304 39212 21332
rect 39071 21301 39083 21304
rect 39025 21295 39083 21301
rect 39206 21292 39212 21304
rect 39264 21292 39270 21344
rect 39945 21335 40003 21341
rect 39945 21301 39957 21335
rect 39991 21332 40003 21335
rect 40034 21332 40040 21344
rect 39991 21304 40040 21332
rect 39991 21301 40003 21304
rect 39945 21295 40003 21301
rect 40034 21292 40040 21304
rect 40092 21292 40098 21344
rect 42702 21292 42708 21344
rect 42760 21292 42766 21344
rect 43438 21292 43444 21344
rect 43496 21292 43502 21344
rect 44818 21292 44824 21344
rect 44876 21292 44882 21344
rect 45830 21292 45836 21344
rect 45888 21332 45894 21344
rect 46474 21332 46480 21344
rect 45888 21304 46480 21332
rect 45888 21292 45894 21304
rect 46474 21292 46480 21304
rect 46532 21292 46538 21344
rect 46750 21292 46756 21344
rect 46808 21292 46814 21344
rect 47578 21292 47584 21344
rect 47636 21292 47642 21344
rect 48498 21292 48504 21344
rect 48556 21292 48562 21344
rect 52822 21292 52828 21344
rect 52880 21292 52886 21344
rect 53837 21335 53895 21341
rect 53837 21301 53849 21335
rect 53883 21332 53895 21335
rect 54478 21332 54484 21344
rect 53883 21304 54484 21332
rect 53883 21301 53895 21304
rect 53837 21295 53895 21301
rect 54478 21292 54484 21304
rect 54536 21292 54542 21344
rect 55950 21292 55956 21344
rect 56008 21292 56014 21344
rect 56042 21292 56048 21344
rect 56100 21292 56106 21344
rect 1104 21242 58880 21264
rect 1104 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 22616 21242
rect 22668 21190 22680 21242
rect 22732 21190 22744 21242
rect 22796 21190 22808 21242
rect 22860 21190 22872 21242
rect 22924 21190 37060 21242
rect 37112 21190 37124 21242
rect 37176 21190 37188 21242
rect 37240 21190 37252 21242
rect 37304 21190 37316 21242
rect 37368 21190 51504 21242
rect 51556 21190 51568 21242
rect 51620 21190 51632 21242
rect 51684 21190 51696 21242
rect 51748 21190 51760 21242
rect 51812 21190 58880 21242
rect 1104 21168 58880 21190
rect 5626 21088 5632 21140
rect 5684 21128 5690 21140
rect 5813 21131 5871 21137
rect 5813 21128 5825 21131
rect 5684 21100 5825 21128
rect 5684 21088 5690 21100
rect 5813 21097 5825 21100
rect 5859 21097 5871 21131
rect 8938 21128 8944 21140
rect 5813 21091 5871 21097
rect 8220 21100 8944 21128
rect 4908 21032 6960 21060
rect 4908 21001 4936 21032
rect 4893 20995 4951 21001
rect 4893 20961 4905 20995
rect 4939 20961 4951 20995
rect 4893 20955 4951 20961
rect 5166 20952 5172 21004
rect 5224 20952 5230 21004
rect 4617 20927 4675 20933
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 5626 20924 5632 20936
rect 4663 20896 5632 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 5626 20884 5632 20896
rect 5684 20884 5690 20936
rect 6546 20884 6552 20936
rect 6604 20884 6610 20936
rect 6932 20933 6960 21032
rect 8220 21001 8248 21100
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 12161 21131 12219 21137
rect 10796 21100 12020 21128
rect 10796 21072 10824 21100
rect 10689 21063 10747 21069
rect 10689 21060 10701 21063
rect 8312 21032 10701 21060
rect 8205 20995 8263 21001
rect 8205 20961 8217 20995
rect 8251 20961 8263 20995
rect 8205 20955 8263 20961
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 8312 20924 8340 21032
rect 10689 21029 10701 21032
rect 10735 21060 10747 21063
rect 10778 21060 10784 21072
rect 10735 21032 10784 21060
rect 10735 21029 10747 21032
rect 10689 21023 10747 21029
rect 10778 21020 10784 21032
rect 10836 21020 10842 21072
rect 11992 21060 12020 21100
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 13446 21128 13452 21140
rect 12207 21100 13452 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 18785 21131 18843 21137
rect 18785 21128 18797 21131
rect 15028 21100 18797 21128
rect 15028 21060 15056 21100
rect 18785 21097 18797 21100
rect 18831 21128 18843 21131
rect 19150 21128 19156 21140
rect 18831 21100 19156 21128
rect 18831 21097 18843 21100
rect 18785 21091 18843 21097
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 27065 21131 27123 21137
rect 27065 21128 27077 21131
rect 22388 21100 27077 21128
rect 22388 21072 22416 21100
rect 27065 21097 27077 21100
rect 27111 21097 27123 21131
rect 27065 21091 27123 21097
rect 27249 21131 27307 21137
rect 27249 21097 27261 21131
rect 27295 21128 27307 21131
rect 27798 21128 27804 21140
rect 27295 21100 27804 21128
rect 27295 21097 27307 21100
rect 27249 21091 27307 21097
rect 11992 21032 15056 21060
rect 15289 21063 15347 21069
rect 15289 21029 15301 21063
rect 15335 21029 15347 21063
rect 15289 21023 15347 21029
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20992 8447 20995
rect 8662 20992 8668 21004
rect 8435 20964 8668 20992
rect 8435 20961 8447 20964
rect 8389 20955 8447 20961
rect 8662 20952 8668 20964
rect 8720 20992 8726 21004
rect 9398 20992 9404 21004
rect 8720 20964 9404 20992
rect 8720 20952 8726 20964
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 14645 20995 14703 21001
rect 14645 20992 14657 20995
rect 14384 20964 14657 20992
rect 6963 20896 8340 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 9122 20884 9128 20936
rect 9180 20884 9186 20936
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20893 10195 20927
rect 10137 20887 10195 20893
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 10870 20924 10876 20936
rect 10827 20896 10876 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 5353 20859 5411 20865
rect 5353 20825 5365 20859
rect 5399 20856 5411 20859
rect 5905 20859 5963 20865
rect 5905 20856 5917 20859
rect 5399 20828 5917 20856
rect 5399 20825 5411 20828
rect 5353 20819 5411 20825
rect 5905 20825 5917 20828
rect 5951 20825 5963 20859
rect 10152 20856 10180 20887
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 12526 20924 12532 20936
rect 10980 20896 12532 20924
rect 10980 20856 11008 20896
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 12802 20884 12808 20936
rect 12860 20884 12866 20936
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13228 20896 13553 20924
rect 13228 20884 13234 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 5905 20819 5963 20825
rect 6104 20828 8156 20856
rect 10152 20828 11008 20856
rect 11048 20859 11106 20865
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 4212 20760 4261 20788
rect 4212 20748 4218 20760
rect 4249 20757 4261 20760
rect 4295 20757 4307 20791
rect 4249 20751 4307 20757
rect 4709 20791 4767 20797
rect 4709 20757 4721 20791
rect 4755 20788 4767 20791
rect 5445 20791 5503 20797
rect 5445 20788 5457 20791
rect 4755 20760 5457 20788
rect 4755 20757 4767 20760
rect 4709 20751 4767 20757
rect 5445 20757 5457 20760
rect 5491 20788 5503 20791
rect 6104 20788 6132 20828
rect 5491 20760 6132 20788
rect 5491 20757 5503 20760
rect 5445 20751 5503 20757
rect 7742 20748 7748 20800
rect 7800 20748 7806 20800
rect 8128 20797 8156 20828
rect 11048 20825 11060 20859
rect 11094 20856 11106 20859
rect 12989 20859 13047 20865
rect 12989 20856 13001 20859
rect 11094 20828 13001 20856
rect 11094 20825 11106 20828
rect 11048 20819 11106 20825
rect 12989 20825 13001 20828
rect 13035 20825 13047 20859
rect 12989 20819 13047 20825
rect 14384 20800 14412 20964
rect 14645 20961 14657 20964
rect 14691 20961 14703 20995
rect 14645 20955 14703 20961
rect 14826 20952 14832 21004
rect 14884 20952 14890 21004
rect 15304 20992 15332 21023
rect 22370 21020 22376 21072
rect 22428 21020 22434 21072
rect 24397 21063 24455 21069
rect 24397 21029 24409 21063
rect 24443 21029 24455 21063
rect 24397 21023 24455 21029
rect 15381 20995 15439 21001
rect 15381 20992 15393 20995
rect 15304 20964 15393 20992
rect 15381 20961 15393 20964
rect 15427 20961 15439 20995
rect 15381 20955 15439 20961
rect 15746 20952 15752 21004
rect 15804 20992 15810 21004
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 15804 20964 17693 20992
rect 15804 20952 15810 20964
rect 17681 20961 17693 20964
rect 17727 20992 17739 20995
rect 18325 20995 18383 21001
rect 18325 20992 18337 20995
rect 17727 20964 18337 20992
rect 17727 20961 17739 20964
rect 17681 20955 17739 20961
rect 18325 20961 18337 20964
rect 18371 20961 18383 20995
rect 18325 20955 18383 20961
rect 24213 20995 24271 21001
rect 24213 20961 24225 20995
rect 24259 20992 24271 20995
rect 24412 20992 24440 21023
rect 24259 20964 24440 20992
rect 24259 20961 24271 20964
rect 24213 20955 24271 20961
rect 24578 20952 24584 21004
rect 24636 20992 24642 21004
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 24636 20964 24961 20992
rect 24636 20952 24642 20964
rect 24949 20961 24961 20964
rect 24995 20961 25007 20995
rect 27080 20992 27108 21091
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 28074 21088 28080 21140
rect 28132 21088 28138 21140
rect 35621 21131 35679 21137
rect 35621 21128 35633 21131
rect 31726 21100 35633 21128
rect 27801 20995 27859 21001
rect 27801 20992 27813 20995
rect 27080 20964 27813 20992
rect 24949 20955 25007 20961
rect 27801 20961 27813 20964
rect 27847 20961 27859 20995
rect 27801 20955 27859 20961
rect 14844 20924 14872 20952
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14844 20896 14933 20924
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 19794 20884 19800 20936
rect 19852 20884 19858 20936
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 22094 20884 22100 20936
rect 22152 20884 22158 20936
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22520 20896 22845 20924
rect 22520 20884 22526 20896
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 24596 20924 24624 20952
rect 23523 20896 24624 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 25222 20884 25228 20936
rect 25280 20884 25286 20936
rect 25866 20884 25872 20936
rect 25924 20884 25930 20936
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20924 27675 20927
rect 28092 20924 28120 21088
rect 30377 21063 30435 21069
rect 30377 21029 30389 21063
rect 30423 21029 30435 21063
rect 30377 21023 30435 21029
rect 30285 20995 30343 21001
rect 30285 20961 30297 20995
rect 30331 20992 30343 20995
rect 30392 20992 30420 21023
rect 30331 20964 30420 20992
rect 31021 20995 31079 21001
rect 30331 20961 30343 20964
rect 30285 20955 30343 20961
rect 31021 20961 31033 20995
rect 31067 20992 31079 20995
rect 31294 20992 31300 21004
rect 31067 20964 31300 20992
rect 31067 20961 31079 20964
rect 31021 20955 31079 20961
rect 31294 20952 31300 20964
rect 31352 20992 31358 21004
rect 31726 20992 31754 21100
rect 35621 21097 35633 21100
rect 35667 21128 35679 21131
rect 35667 21100 37228 21128
rect 35667 21097 35679 21100
rect 35621 21091 35679 21097
rect 36541 21063 36599 21069
rect 36541 21029 36553 21063
rect 36587 21029 36599 21063
rect 36541 21023 36599 21029
rect 31352 20964 31754 20992
rect 36449 20995 36507 21001
rect 31352 20952 31358 20964
rect 36449 20961 36461 20995
rect 36495 20992 36507 20995
rect 36556 20992 36584 21023
rect 36722 21020 36728 21072
rect 36780 21060 36786 21072
rect 36780 21032 36952 21060
rect 36780 21020 36786 21032
rect 36495 20964 36584 20992
rect 36495 20961 36507 20964
rect 36449 20955 36507 20961
rect 27663 20896 28120 20924
rect 27663 20893 27675 20896
rect 27617 20887 27675 20893
rect 28626 20884 28632 20936
rect 28684 20884 28690 20936
rect 31846 20884 31852 20936
rect 31904 20884 31910 20936
rect 34241 20927 34299 20933
rect 34241 20924 34253 20927
rect 32140 20896 34253 20924
rect 18141 20859 18199 20865
rect 18141 20825 18153 20859
rect 18187 20856 18199 20859
rect 20340 20859 20398 20865
rect 18187 20828 18736 20856
rect 18187 20825 18199 20828
rect 18141 20819 18199 20825
rect 18708 20800 18736 20828
rect 20340 20825 20352 20859
rect 20386 20856 20398 20859
rect 22281 20859 22339 20865
rect 22281 20856 22293 20859
rect 20386 20828 22293 20856
rect 20386 20825 20398 20828
rect 20340 20819 20398 20825
rect 22281 20825 22293 20828
rect 22327 20825 22339 20859
rect 22281 20819 22339 20825
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 25038 20856 25044 20868
rect 24811 20828 25044 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 25038 20816 25044 20828
rect 25096 20816 25102 20868
rect 27709 20859 27767 20865
rect 27709 20856 27721 20859
rect 26804 20828 27721 20856
rect 8113 20791 8171 20797
rect 8113 20757 8125 20791
rect 8159 20788 8171 20791
rect 9030 20788 9036 20800
rect 8159 20760 9036 20788
rect 8159 20757 8171 20760
rect 8113 20751 8171 20757
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 9766 20748 9772 20800
rect 9824 20748 9830 20800
rect 12250 20748 12256 20800
rect 12308 20748 12314 20800
rect 14366 20748 14372 20800
rect 14424 20748 14430 20800
rect 14826 20748 14832 20800
rect 14884 20748 14890 20800
rect 16022 20748 16028 20800
rect 16080 20748 16086 20800
rect 17770 20748 17776 20800
rect 17828 20748 17834 20800
rect 18230 20748 18236 20800
rect 18288 20748 18294 20800
rect 18690 20748 18696 20800
rect 18748 20748 18754 20800
rect 19242 20748 19248 20800
rect 19300 20748 19306 20800
rect 21450 20748 21456 20800
rect 21508 20748 21514 20800
rect 21542 20748 21548 20800
rect 21600 20748 21606 20800
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20788 23627 20791
rect 23658 20788 23664 20800
rect 23615 20760 23664 20788
rect 23615 20757 23627 20760
rect 23569 20751 23627 20757
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 24670 20748 24676 20800
rect 24728 20788 24734 20800
rect 24857 20791 24915 20797
rect 24857 20788 24869 20791
rect 24728 20760 24869 20788
rect 24728 20748 24734 20760
rect 24857 20757 24869 20760
rect 24903 20788 24915 20791
rect 26804 20788 26832 20828
rect 27709 20825 27721 20828
rect 27755 20856 27767 20859
rect 27890 20856 27896 20868
rect 27755 20828 27896 20856
rect 27755 20825 27767 20828
rect 27709 20819 27767 20825
rect 27890 20816 27896 20828
rect 27948 20816 27954 20868
rect 30745 20859 30803 20865
rect 30745 20825 30757 20859
rect 30791 20856 30803 20859
rect 31478 20856 31484 20868
rect 30791 20828 31484 20856
rect 30791 20825 30803 20828
rect 30745 20819 30803 20825
rect 31478 20816 31484 20828
rect 31536 20816 31542 20868
rect 32140 20800 32168 20896
rect 34241 20893 34253 20896
rect 34287 20924 34299 20927
rect 34514 20924 34520 20936
rect 34287 20896 34520 20924
rect 34287 20893 34299 20896
rect 34241 20887 34299 20893
rect 34514 20884 34520 20896
rect 34572 20884 34578 20936
rect 35250 20884 35256 20936
rect 35308 20884 35314 20936
rect 36924 20933 36952 21032
rect 36998 20952 37004 21004
rect 37056 20992 37062 21004
rect 37093 20995 37151 21001
rect 37093 20992 37105 20995
rect 37056 20964 37105 20992
rect 37056 20952 37062 20964
rect 37093 20961 37105 20964
rect 37139 20961 37151 20995
rect 37200 20992 37228 21100
rect 38010 21088 38016 21140
rect 38068 21088 38074 21140
rect 39850 21088 39856 21140
rect 39908 21088 39914 21140
rect 43438 21088 43444 21140
rect 43496 21088 43502 21140
rect 45925 21131 45983 21137
rect 45925 21097 45937 21131
rect 45971 21128 45983 21131
rect 46106 21128 46112 21140
rect 45971 21100 46112 21128
rect 45971 21097 45983 21100
rect 45925 21091 45983 21097
rect 46106 21088 46112 21100
rect 46164 21088 46170 21140
rect 47578 21128 47584 21140
rect 46308 21100 47584 21128
rect 37461 20995 37519 21001
rect 37461 20992 37473 20995
rect 37200 20964 37473 20992
rect 37093 20955 37151 20961
rect 37461 20961 37473 20964
rect 37507 20961 37519 20995
rect 37461 20955 37519 20961
rect 37645 20995 37703 21001
rect 37645 20961 37657 20995
rect 37691 20992 37703 20995
rect 38028 20992 38056 21088
rect 37691 20964 38056 20992
rect 37691 20961 37703 20964
rect 37645 20955 37703 20961
rect 39206 20952 39212 21004
rect 39264 20952 39270 21004
rect 41386 20964 42380 20992
rect 36909 20927 36967 20933
rect 36909 20893 36921 20927
rect 36955 20893 36967 20927
rect 36909 20887 36967 20893
rect 41233 20927 41291 20933
rect 41233 20893 41245 20927
rect 41279 20924 41291 20927
rect 41386 20924 41414 20964
rect 41279 20896 41414 20924
rect 41279 20893 41291 20896
rect 41233 20887 41291 20893
rect 41874 20884 41880 20936
rect 41932 20884 41938 20936
rect 42352 20933 42380 20964
rect 42337 20927 42395 20933
rect 42337 20893 42349 20927
rect 42383 20924 42395 20927
rect 42426 20924 42432 20936
rect 42383 20896 42432 20924
rect 42383 20893 42395 20896
rect 42337 20887 42395 20893
rect 42426 20884 42432 20896
rect 42484 20884 42490 20936
rect 42604 20927 42662 20933
rect 42604 20893 42616 20927
rect 42650 20924 42662 20927
rect 43456 20924 43484 21088
rect 43717 21063 43775 21069
rect 43717 21029 43729 21063
rect 43763 21060 43775 21063
rect 43763 21032 44128 21060
rect 43763 21029 43775 21032
rect 43717 21023 43775 21029
rect 44100 21004 44128 21032
rect 44082 20952 44088 21004
rect 44140 20952 44146 21004
rect 42650 20896 43484 20924
rect 42650 20893 42662 20896
rect 42604 20887 42662 20893
rect 44174 20884 44180 20936
rect 44232 20924 44238 20936
rect 46308 20933 46336 21100
rect 47578 21088 47584 21100
rect 47636 21088 47642 21140
rect 49142 21088 49148 21140
rect 49200 21128 49206 21140
rect 49329 21131 49387 21137
rect 49329 21128 49341 21131
rect 49200 21100 49341 21128
rect 49200 21088 49206 21100
rect 49329 21097 49341 21100
rect 49375 21097 49387 21131
rect 49329 21091 49387 21097
rect 51994 21088 52000 21140
rect 52052 21088 52058 21140
rect 52822 21088 52828 21140
rect 52880 21088 52886 21140
rect 56045 21131 56103 21137
rect 56045 21097 56057 21131
rect 56091 21128 56103 21131
rect 56594 21128 56600 21140
rect 56091 21100 56600 21128
rect 56091 21097 56103 21100
rect 56045 21091 56103 21097
rect 56594 21088 56600 21100
rect 56652 21088 56658 21140
rect 46474 20952 46480 21004
rect 46532 20952 46538 21004
rect 46934 20952 46940 21004
rect 46992 20952 46998 21004
rect 48774 20952 48780 21004
rect 48832 20992 48838 21004
rect 49605 20995 49663 21001
rect 49605 20992 49617 20995
rect 48832 20964 49617 20992
rect 48832 20952 48838 20964
rect 49605 20961 49617 20964
rect 49651 20961 49663 20995
rect 52012 20992 52040 21088
rect 52273 20995 52331 21001
rect 52273 20992 52285 20995
rect 52012 20964 52285 20992
rect 49605 20955 49663 20961
rect 52273 20961 52285 20964
rect 52319 20961 52331 20995
rect 52273 20955 52331 20961
rect 52457 20995 52515 21001
rect 52457 20961 52469 20995
rect 52503 20992 52515 20995
rect 52840 20992 52868 21088
rect 52503 20964 52868 20992
rect 52503 20961 52515 20964
rect 52457 20955 52515 20961
rect 53834 20952 53840 21004
rect 53892 20992 53898 21004
rect 54389 20995 54447 21001
rect 54389 20992 54401 20995
rect 53892 20964 54401 20992
rect 53892 20952 53898 20964
rect 54389 20961 54401 20964
rect 54435 20992 54447 20995
rect 54662 20992 54668 21004
rect 54435 20964 54668 20992
rect 54435 20961 54447 20964
rect 54389 20955 54447 20961
rect 54662 20952 54668 20964
rect 54720 20952 54726 21004
rect 55401 20995 55459 21001
rect 55401 20992 55413 20995
rect 55048 20964 55413 20992
rect 44361 20927 44419 20933
rect 44361 20924 44373 20927
rect 44232 20896 44373 20924
rect 44232 20884 44238 20896
rect 44361 20893 44373 20896
rect 44407 20893 44419 20927
rect 44361 20887 44419 20893
rect 46293 20927 46351 20933
rect 46293 20893 46305 20927
rect 46339 20893 46351 20927
rect 46293 20887 46351 20893
rect 46385 20927 46443 20933
rect 46385 20893 46397 20927
rect 46431 20924 46443 20927
rect 47121 20927 47179 20933
rect 47121 20924 47133 20927
rect 46431 20896 47133 20924
rect 46431 20893 46443 20896
rect 46385 20887 46443 20893
rect 47121 20893 47133 20896
rect 47167 20924 47179 20927
rect 47167 20896 47716 20924
rect 47167 20893 47179 20896
rect 47121 20887 47179 20893
rect 32585 20859 32643 20865
rect 32585 20825 32597 20859
rect 32631 20856 32643 20859
rect 33502 20856 33508 20868
rect 32631 20828 33508 20856
rect 32631 20825 32643 20828
rect 32585 20819 32643 20825
rect 33502 20816 33508 20828
rect 33560 20816 33566 20868
rect 33996 20859 34054 20865
rect 33996 20825 34008 20859
rect 34042 20856 34054 20859
rect 34606 20856 34612 20868
rect 34042 20828 34612 20856
rect 34042 20825 34054 20828
rect 33996 20819 34054 20825
rect 34606 20816 34612 20828
rect 34664 20816 34670 20868
rect 38933 20859 38991 20865
rect 38933 20856 38945 20859
rect 37752 20828 38945 20856
rect 24903 20760 26832 20788
rect 24903 20757 24915 20760
rect 24857 20751 24915 20757
rect 28074 20748 28080 20800
rect 28132 20748 28138 20800
rect 28994 20748 29000 20800
rect 29052 20748 29058 20800
rect 29638 20748 29644 20800
rect 29696 20748 29702 20800
rect 30834 20748 30840 20800
rect 30892 20748 30898 20800
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 32122 20748 32128 20800
rect 32180 20748 32186 20800
rect 32861 20791 32919 20797
rect 32861 20757 32873 20791
rect 32907 20788 32919 20791
rect 33410 20788 33416 20800
rect 32907 20760 33416 20788
rect 32907 20757 32919 20760
rect 32861 20751 32919 20757
rect 33410 20748 33416 20760
rect 33468 20788 33474 20800
rect 33778 20788 33784 20800
rect 33468 20760 33784 20788
rect 33468 20748 33474 20760
rect 33778 20748 33784 20760
rect 33836 20748 33842 20800
rect 34698 20748 34704 20800
rect 34756 20748 34762 20800
rect 35805 20791 35863 20797
rect 35805 20757 35817 20791
rect 35851 20788 35863 20791
rect 35986 20788 35992 20800
rect 35851 20760 35992 20788
rect 35851 20757 35863 20760
rect 35805 20751 35863 20757
rect 35986 20748 35992 20760
rect 36044 20748 36050 20800
rect 37001 20791 37059 20797
rect 37001 20757 37013 20791
rect 37047 20788 37059 20791
rect 37550 20788 37556 20800
rect 37047 20760 37556 20788
rect 37047 20757 37059 20760
rect 37001 20751 37059 20757
rect 37550 20748 37556 20760
rect 37608 20788 37614 20800
rect 37752 20797 37780 20828
rect 38933 20825 38945 20828
rect 38979 20856 38991 20859
rect 39942 20856 39948 20868
rect 38979 20828 39948 20856
rect 38979 20825 38991 20828
rect 38933 20819 38991 20825
rect 39942 20816 39948 20828
rect 40000 20816 40006 20868
rect 40988 20859 41046 20865
rect 40988 20825 41000 20859
rect 41034 20856 41046 20859
rect 41325 20859 41383 20865
rect 41325 20856 41337 20859
rect 41034 20828 41337 20856
rect 41034 20825 41046 20828
rect 40988 20819 41046 20825
rect 41325 20825 41337 20828
rect 41371 20825 41383 20859
rect 41325 20819 41383 20825
rect 47029 20859 47087 20865
rect 47029 20825 47041 20859
rect 47075 20856 47087 20859
rect 47581 20859 47639 20865
rect 47581 20856 47593 20859
rect 47075 20828 47593 20856
rect 47075 20825 47087 20828
rect 47029 20819 47087 20825
rect 47581 20825 47593 20828
rect 47627 20825 47639 20859
rect 47688 20856 47716 20896
rect 47762 20884 47768 20936
rect 47820 20924 47826 20936
rect 48133 20927 48191 20933
rect 48133 20924 48145 20927
rect 47820 20896 48145 20924
rect 47820 20884 47826 20896
rect 48133 20893 48145 20896
rect 48179 20893 48191 20927
rect 48133 20887 48191 20893
rect 49418 20884 49424 20936
rect 49476 20924 49482 20936
rect 50709 20927 50767 20933
rect 50709 20924 50721 20927
rect 49476 20896 50721 20924
rect 49476 20884 49482 20896
rect 50709 20893 50721 20896
rect 50755 20893 50767 20927
rect 50709 20887 50767 20893
rect 51258 20884 51264 20936
rect 51316 20924 51322 20936
rect 51445 20927 51503 20933
rect 51445 20924 51457 20927
rect 51316 20896 51457 20924
rect 51316 20884 51322 20896
rect 51445 20893 51457 20896
rect 51491 20893 51503 20927
rect 51445 20887 51503 20893
rect 53466 20884 53472 20936
rect 53524 20924 53530 20936
rect 53561 20927 53619 20933
rect 53561 20924 53573 20927
rect 53524 20896 53573 20924
rect 53524 20884 53530 20896
rect 53561 20893 53573 20896
rect 53607 20893 53619 20927
rect 53561 20887 53619 20893
rect 48869 20859 48927 20865
rect 47688 20828 47900 20856
rect 47581 20819 47639 20825
rect 37737 20791 37795 20797
rect 37737 20788 37749 20791
rect 37608 20760 37749 20788
rect 37608 20748 37614 20760
rect 37737 20757 37749 20760
rect 37783 20757 37795 20791
rect 37737 20751 37795 20757
rect 38102 20748 38108 20800
rect 38160 20748 38166 20800
rect 38470 20748 38476 20800
rect 38528 20748 38534 20800
rect 38562 20748 38568 20800
rect 38620 20748 38626 20800
rect 39022 20748 39028 20800
rect 39080 20748 39086 20800
rect 39669 20791 39727 20797
rect 39669 20757 39681 20791
rect 39715 20788 39727 20791
rect 39758 20788 39764 20800
rect 39715 20760 39764 20788
rect 39715 20757 39727 20760
rect 39669 20751 39727 20757
rect 39758 20748 39764 20760
rect 39816 20748 39822 20800
rect 43806 20748 43812 20800
rect 43864 20748 43870 20800
rect 44821 20791 44879 20797
rect 44821 20757 44833 20791
rect 44867 20788 44879 20791
rect 45002 20788 45008 20800
rect 44867 20760 45008 20788
rect 44867 20757 44879 20760
rect 44821 20751 44879 20757
rect 45002 20748 45008 20760
rect 45060 20788 45066 20800
rect 45189 20791 45247 20797
rect 45189 20788 45201 20791
rect 45060 20760 45201 20788
rect 45060 20748 45066 20760
rect 45189 20757 45201 20760
rect 45235 20788 45247 20791
rect 45741 20791 45799 20797
rect 45741 20788 45753 20791
rect 45235 20760 45753 20788
rect 45235 20757 45247 20760
rect 45189 20751 45247 20757
rect 45741 20757 45753 20760
rect 45787 20757 45799 20791
rect 45741 20751 45799 20757
rect 47486 20748 47492 20800
rect 47544 20748 47550 20800
rect 47872 20788 47900 20828
rect 48869 20825 48881 20859
rect 48915 20856 48927 20859
rect 50157 20859 50215 20865
rect 50157 20856 50169 20859
rect 48915 20828 50169 20856
rect 48915 20825 48927 20828
rect 48869 20819 48927 20825
rect 50157 20825 50169 20828
rect 50203 20825 50215 20859
rect 50157 20819 50215 20825
rect 55048 20800 55076 20964
rect 55401 20961 55413 20964
rect 55447 20961 55459 20995
rect 55401 20955 55459 20961
rect 55950 20952 55956 21004
rect 56008 20992 56014 21004
rect 56689 20995 56747 21001
rect 56689 20992 56701 20995
rect 56008 20964 56701 20992
rect 56008 20952 56014 20964
rect 56689 20961 56701 20964
rect 56735 20961 56747 20995
rect 56689 20955 56747 20961
rect 55585 20927 55643 20933
rect 55585 20893 55597 20927
rect 55631 20924 55643 20927
rect 56965 20927 57023 20933
rect 56965 20924 56977 20927
rect 55631 20896 56977 20924
rect 55631 20893 55643 20896
rect 55585 20887 55643 20893
rect 56965 20893 56977 20896
rect 57011 20893 57023 20927
rect 56965 20887 57023 20893
rect 57514 20884 57520 20936
rect 57572 20884 57578 20936
rect 56505 20859 56563 20865
rect 55692 20828 56272 20856
rect 48961 20791 49019 20797
rect 48961 20788 48973 20791
rect 47872 20760 48973 20788
rect 48961 20757 48973 20760
rect 49007 20788 49019 20791
rect 49326 20788 49332 20800
rect 49007 20760 49332 20788
rect 49007 20757 49019 20760
rect 48961 20751 49019 20757
rect 49326 20748 49332 20760
rect 49384 20748 49390 20800
rect 50890 20748 50896 20800
rect 50948 20748 50954 20800
rect 51902 20748 51908 20800
rect 51960 20748 51966 20800
rect 52546 20748 52552 20800
rect 52604 20748 52610 20800
rect 52914 20748 52920 20800
rect 52972 20748 52978 20800
rect 53006 20748 53012 20800
rect 53064 20748 53070 20800
rect 53742 20748 53748 20800
rect 53800 20748 53806 20800
rect 55030 20748 55036 20800
rect 55088 20748 55094 20800
rect 55582 20748 55588 20800
rect 55640 20788 55646 20800
rect 55692 20797 55720 20828
rect 55677 20791 55735 20797
rect 55677 20788 55689 20791
rect 55640 20760 55689 20788
rect 55640 20748 55646 20760
rect 55677 20757 55689 20760
rect 55723 20757 55735 20791
rect 55677 20751 55735 20757
rect 56134 20748 56140 20800
rect 56192 20748 56198 20800
rect 56244 20788 56272 20828
rect 56505 20825 56517 20859
rect 56551 20856 56563 20859
rect 56778 20856 56784 20868
rect 56551 20828 56784 20856
rect 56551 20825 56563 20828
rect 56505 20819 56563 20825
rect 56778 20816 56784 20828
rect 56836 20816 56842 20868
rect 56597 20791 56655 20797
rect 56597 20788 56609 20791
rect 56244 20760 56609 20788
rect 56597 20757 56609 20760
rect 56643 20757 56655 20791
rect 56597 20751 56655 20757
rect 1104 20698 59040 20720
rect 1104 20646 15394 20698
rect 15446 20646 15458 20698
rect 15510 20646 15522 20698
rect 15574 20646 15586 20698
rect 15638 20646 15650 20698
rect 15702 20646 29838 20698
rect 29890 20646 29902 20698
rect 29954 20646 29966 20698
rect 30018 20646 30030 20698
rect 30082 20646 30094 20698
rect 30146 20646 44282 20698
rect 44334 20646 44346 20698
rect 44398 20646 44410 20698
rect 44462 20646 44474 20698
rect 44526 20646 44538 20698
rect 44590 20646 58726 20698
rect 58778 20646 58790 20698
rect 58842 20646 58854 20698
rect 58906 20646 58918 20698
rect 58970 20646 58982 20698
rect 59034 20646 59040 20698
rect 1104 20624 59040 20646
rect 6917 20587 6975 20593
rect 6917 20553 6929 20587
rect 6963 20584 6975 20587
rect 8570 20584 8576 20596
rect 6963 20556 8576 20584
rect 6963 20553 6975 20556
rect 6917 20547 6975 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 8849 20587 8907 20593
rect 8849 20553 8861 20587
rect 8895 20584 8907 20587
rect 9122 20584 9128 20596
rect 8895 20556 9128 20584
rect 8895 20553 8907 20556
rect 8849 20547 8907 20553
rect 4792 20519 4850 20525
rect 4792 20485 4804 20519
rect 4838 20516 4850 20519
rect 4982 20516 4988 20528
rect 4838 20488 4988 20516
rect 4838 20485 4850 20488
rect 4792 20479 4850 20485
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 8864 20448 8892 20547
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11606 20584 11612 20596
rect 11011 20556 11612 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 11793 20587 11851 20593
rect 11793 20553 11805 20587
rect 11839 20584 11851 20587
rect 12250 20584 12256 20596
rect 11839 20556 12256 20584
rect 11839 20553 11851 20556
rect 11793 20547 11851 20553
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 14366 20584 14372 20596
rect 12406 20556 14372 20584
rect 10870 20516 10876 20528
rect 10244 20488 10876 20516
rect 9490 20448 9496 20460
rect 8619 20420 8892 20448
rect 8956 20420 9496 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4154 20380 4160 20392
rect 3927 20352 4160 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 4525 20383 4583 20389
rect 4525 20380 4537 20383
rect 4304 20352 4537 20380
rect 4304 20340 4310 20352
rect 4525 20349 4537 20352
rect 4571 20349 4583 20383
rect 4525 20343 4583 20349
rect 7558 20340 7564 20392
rect 7616 20340 7622 20392
rect 7650 20340 7656 20392
rect 7708 20389 7714 20392
rect 7708 20383 7757 20389
rect 7708 20349 7711 20383
rect 7745 20349 7757 20383
rect 7708 20343 7757 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20380 7895 20383
rect 7883 20352 8064 20380
rect 7883 20349 7895 20352
rect 7837 20343 7895 20349
rect 7708 20340 7714 20343
rect 5905 20315 5963 20321
rect 5905 20281 5917 20315
rect 5951 20312 5963 20315
rect 6546 20312 6552 20324
rect 5951 20284 6552 20312
rect 5951 20281 5963 20284
rect 5905 20275 5963 20281
rect 6546 20272 6552 20284
rect 6604 20312 6610 20324
rect 6604 20284 7052 20312
rect 6604 20272 6610 20284
rect 4430 20204 4436 20256
rect 4488 20204 4494 20256
rect 7024 20244 7052 20284
rect 8036 20244 8064 20352
rect 8754 20340 8760 20392
rect 8812 20380 8818 20392
rect 8956 20380 8984 20420
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 9973 20451 10031 20457
rect 9973 20417 9985 20451
rect 10019 20448 10031 20451
rect 10134 20448 10140 20460
rect 10019 20420 10140 20448
rect 10019 20417 10031 20420
rect 9973 20411 10031 20417
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 10244 20457 10272 20488
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 12406 20516 12434 20556
rect 14366 20544 14372 20556
rect 14424 20544 14430 20596
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 15194 20584 15200 20596
rect 14691 20556 15200 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 11112 20488 12434 20516
rect 11112 20476 11118 20488
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 11698 20448 11704 20460
rect 10229 20411 10287 20417
rect 10888 20420 11704 20448
rect 8812 20352 8984 20380
rect 8812 20340 8818 20352
rect 10778 20340 10784 20392
rect 10836 20340 10842 20392
rect 10888 20389 10916 20420
rect 11698 20408 11704 20420
rect 11756 20448 11762 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11756 20420 11897 20448
rect 11756 20408 11762 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 13446 20408 13452 20460
rect 13504 20457 13510 20460
rect 13504 20451 13553 20457
rect 13504 20417 13507 20451
rect 13541 20417 13553 20451
rect 13504 20411 13553 20417
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20448 14427 20451
rect 14660 20448 14688 20547
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 18598 20544 18604 20596
rect 18656 20544 18662 20596
rect 18969 20587 19027 20593
rect 18969 20553 18981 20587
rect 19015 20584 19027 20587
rect 19242 20584 19248 20596
rect 19015 20556 19248 20584
rect 19015 20553 19027 20556
rect 18969 20547 19027 20553
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 20530 20584 20536 20596
rect 19852 20556 20536 20584
rect 19852 20544 19858 20556
rect 20530 20544 20536 20556
rect 20588 20544 20594 20596
rect 21821 20587 21879 20593
rect 21821 20553 21833 20587
rect 21867 20584 21879 20587
rect 22094 20584 22100 20596
rect 21867 20556 22100 20584
rect 21867 20553 21879 20556
rect 21821 20547 21879 20553
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 24857 20587 24915 20593
rect 24857 20553 24869 20587
rect 24903 20584 24915 20587
rect 25866 20584 25872 20596
rect 24903 20556 25872 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 28350 20584 28356 20596
rect 26620 20556 28356 20584
rect 15780 20519 15838 20525
rect 15780 20485 15792 20519
rect 15826 20516 15838 20519
rect 16040 20516 16068 20544
rect 15826 20488 16068 20516
rect 17396 20519 17454 20525
rect 15826 20485 15838 20488
rect 15780 20479 15838 20485
rect 17396 20485 17408 20519
rect 17442 20516 17454 20519
rect 18046 20516 18052 20528
rect 17442 20488 18052 20516
rect 17442 20485 17454 20488
rect 17396 20479 17454 20485
rect 18046 20476 18052 20488
rect 18104 20476 18110 20528
rect 14415 20420 14688 20448
rect 14415 20417 14427 20420
rect 14369 20411 14427 20417
rect 13504 20408 13510 20411
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 20530 20457 20536 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15988 20420 16037 20448
rect 15988 20408 15994 20420
rect 16025 20417 16037 20420
rect 16071 20448 16083 20451
rect 17129 20451 17187 20457
rect 17129 20448 17141 20451
rect 16071 20420 17141 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 17129 20417 17141 20420
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 20508 20451 20536 20457
rect 20508 20417 20520 20451
rect 20508 20411 20536 20417
rect 20530 20408 20536 20411
rect 20588 20408 20594 20460
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 21545 20451 21603 20457
rect 21545 20448 21557 20451
rect 21508 20420 21557 20448
rect 21508 20408 21514 20420
rect 21545 20417 21557 20420
rect 21591 20417 21603 20451
rect 21545 20411 21603 20417
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22235 20420 22661 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 23566 20408 23572 20460
rect 23624 20448 23630 20460
rect 23733 20451 23791 20457
rect 23733 20448 23745 20451
rect 23624 20420 23745 20448
rect 23624 20408 23630 20420
rect 23733 20417 23745 20420
rect 23779 20417 23791 20451
rect 23733 20411 23791 20417
rect 25590 20408 25596 20460
rect 25648 20408 25654 20460
rect 25866 20408 25872 20460
rect 25924 20408 25930 20460
rect 26620 20457 26648 20556
rect 28350 20544 28356 20556
rect 28408 20544 28414 20596
rect 28445 20587 28503 20593
rect 28445 20553 28457 20587
rect 28491 20584 28503 20587
rect 28626 20584 28632 20596
rect 28491 20556 28632 20584
rect 28491 20553 28503 20556
rect 28445 20547 28503 20553
rect 28626 20544 28632 20556
rect 28684 20544 28690 20596
rect 29733 20587 29791 20593
rect 29733 20553 29745 20587
rect 29779 20584 29791 20587
rect 30742 20584 30748 20596
rect 29779 20556 30748 20584
rect 29779 20553 29791 20556
rect 29733 20547 29791 20553
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 31202 20584 31208 20596
rect 31036 20556 31208 20584
rect 27246 20525 27252 20528
rect 27240 20516 27252 20525
rect 27207 20488 27252 20516
rect 27240 20479 27252 20488
rect 27246 20476 27252 20479
rect 27304 20476 27310 20528
rect 27890 20476 27896 20528
rect 27948 20516 27954 20528
rect 28813 20519 28871 20525
rect 28813 20516 28825 20519
rect 27948 20488 28825 20516
rect 27948 20476 27954 20488
rect 28813 20485 28825 20488
rect 28859 20485 28871 20519
rect 28813 20479 28871 20485
rect 30190 20476 30196 20528
rect 30248 20476 30254 20528
rect 30868 20519 30926 20525
rect 30868 20485 30880 20519
rect 30914 20516 30926 20519
rect 31036 20516 31064 20556
rect 31202 20544 31208 20556
rect 31260 20544 31266 20596
rect 31386 20544 31392 20596
rect 31444 20584 31450 20596
rect 31573 20587 31631 20593
rect 31573 20584 31585 20587
rect 31444 20556 31585 20584
rect 31444 20544 31450 20556
rect 31573 20553 31585 20556
rect 31619 20553 31631 20587
rect 31573 20547 31631 20553
rect 31846 20544 31852 20596
rect 31904 20584 31910 20596
rect 31941 20587 31999 20593
rect 31941 20584 31953 20587
rect 31904 20556 31953 20584
rect 31904 20544 31910 20556
rect 31941 20553 31953 20556
rect 31987 20553 31999 20587
rect 35250 20584 35256 20596
rect 31941 20547 31999 20553
rect 34164 20556 35256 20584
rect 32122 20516 32128 20528
rect 30914 20488 31064 20516
rect 31128 20488 32128 20516
rect 30914 20485 30926 20488
rect 30868 20479 30926 20485
rect 26605 20451 26663 20457
rect 26605 20417 26617 20451
rect 26651 20417 26663 20451
rect 26605 20411 26663 20417
rect 26789 20451 26847 20457
rect 26789 20417 26801 20451
rect 26835 20448 26847 20451
rect 27706 20448 27712 20460
rect 26835 20420 27712 20448
rect 26835 20417 26847 20420
rect 26789 20411 26847 20417
rect 27706 20408 27712 20420
rect 27764 20408 27770 20460
rect 29641 20451 29699 20457
rect 29641 20417 29653 20451
rect 29687 20448 29699 20451
rect 30208 20448 30236 20476
rect 31128 20457 31156 20488
rect 32122 20476 32128 20488
rect 32180 20476 32186 20528
rect 34164 20460 34192 20556
rect 35250 20544 35256 20556
rect 35308 20544 35314 20596
rect 37093 20587 37151 20593
rect 37093 20553 37105 20587
rect 37139 20584 37151 20587
rect 37642 20584 37648 20596
rect 37139 20556 37648 20584
rect 37139 20553 37151 20556
rect 37093 20547 37151 20553
rect 37642 20544 37648 20556
rect 37700 20544 37706 20596
rect 37918 20544 37924 20596
rect 37976 20584 37982 20596
rect 38470 20584 38476 20596
rect 37976 20556 38476 20584
rect 37976 20544 37982 20556
rect 38470 20544 38476 20556
rect 38528 20584 38534 20596
rect 38838 20584 38844 20596
rect 38528 20556 38844 20584
rect 38528 20544 38534 20556
rect 38838 20544 38844 20556
rect 38896 20544 38902 20596
rect 39942 20544 39948 20596
rect 40000 20544 40006 20596
rect 40034 20544 40040 20596
rect 40092 20544 40098 20596
rect 40405 20587 40463 20593
rect 40405 20553 40417 20587
rect 40451 20584 40463 20587
rect 41874 20584 41880 20596
rect 40451 20556 41880 20584
rect 40451 20553 40463 20556
rect 40405 20547 40463 20553
rect 41874 20544 41880 20556
rect 41932 20544 41938 20596
rect 43809 20587 43867 20593
rect 43809 20553 43821 20587
rect 43855 20584 43867 20587
rect 44174 20584 44180 20596
rect 43855 20556 44180 20584
rect 43855 20553 43867 20556
rect 43809 20547 43867 20553
rect 44174 20544 44180 20556
rect 44232 20544 44238 20596
rect 47305 20587 47363 20593
rect 44284 20556 46980 20584
rect 34514 20476 34520 20528
rect 34572 20516 34578 20528
rect 37461 20519 37519 20525
rect 37461 20516 37473 20519
rect 34572 20488 37473 20516
rect 34572 20476 34578 20488
rect 35728 20460 35756 20488
rect 37461 20485 37473 20488
rect 37507 20485 37519 20519
rect 37461 20479 37519 20485
rect 31113 20451 31171 20457
rect 29687 20420 31064 20448
rect 29687 20417 29699 20420
rect 29641 20411 29699 20417
rect 10873 20383 10931 20389
rect 10873 20349 10885 20383
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 11609 20383 11667 20389
rect 11609 20349 11621 20383
rect 11655 20380 11667 20383
rect 12066 20380 12072 20392
rect 11655 20352 12072 20380
rect 11655 20349 11667 20352
rect 11609 20343 11667 20349
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 13170 20380 13176 20392
rect 12406 20352 13176 20380
rect 8110 20272 8116 20324
rect 8168 20272 8174 20324
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 12406 20312 12434 20352
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 13354 20340 13360 20392
rect 13412 20340 13418 20392
rect 13630 20340 13636 20392
rect 13688 20340 13694 20392
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 11379 20284 12434 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 13909 20315 13967 20321
rect 13909 20312 13921 20315
rect 13872 20284 13921 20312
rect 13872 20272 13878 20284
rect 13909 20281 13921 20284
rect 13955 20281 13967 20315
rect 13909 20275 13967 20281
rect 14090 20272 14096 20324
rect 14148 20312 14154 20324
rect 14568 20312 14596 20343
rect 18690 20340 18696 20392
rect 18748 20380 18754 20392
rect 19061 20383 19119 20389
rect 19061 20380 19073 20383
rect 18748 20352 19073 20380
rect 18748 20340 18754 20352
rect 19061 20349 19073 20352
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 19150 20340 19156 20392
rect 19208 20340 19214 20392
rect 20346 20340 20352 20392
rect 20404 20380 20410 20392
rect 20404 20352 20449 20380
rect 20404 20340 20410 20352
rect 20622 20340 20628 20392
rect 20680 20340 20686 20392
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21726 20380 21732 20392
rect 21407 20352 21732 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 21726 20340 21732 20352
rect 21784 20380 21790 20392
rect 21784 20352 22094 20380
rect 21784 20340 21790 20352
rect 14148 20284 14596 20312
rect 14148 20272 14154 20284
rect 7024 20216 8064 20244
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 12253 20247 12311 20253
rect 12253 20244 12265 20247
rect 12216 20216 12265 20244
rect 12216 20204 12222 20216
rect 12253 20213 12265 20216
rect 12299 20213 12311 20247
rect 12253 20207 12311 20213
rect 12618 20204 12624 20256
rect 12676 20204 12682 20256
rect 12713 20247 12771 20253
rect 12713 20213 12725 20247
rect 12759 20244 12771 20247
rect 14458 20244 14464 20256
rect 12759 20216 14464 20244
rect 12759 20213 12771 20216
rect 12713 20207 12771 20213
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 14568 20244 14596 20284
rect 18509 20315 18567 20321
rect 18509 20281 18521 20315
rect 18555 20312 18567 20315
rect 19794 20312 19800 20324
rect 18555 20284 19800 20312
rect 18555 20281 18567 20284
rect 18509 20275 18567 20281
rect 19794 20272 19800 20284
rect 19852 20272 19858 20324
rect 20806 20272 20812 20324
rect 20864 20312 20870 20324
rect 20901 20315 20959 20321
rect 20901 20312 20913 20315
rect 20864 20284 20913 20312
rect 20864 20272 20870 20284
rect 20901 20281 20913 20284
rect 20947 20281 20959 20315
rect 22066 20312 22094 20352
rect 22278 20340 22284 20392
rect 22336 20340 22342 20392
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 23216 20312 23244 20343
rect 23474 20340 23480 20392
rect 23532 20340 23538 20392
rect 25774 20389 25780 20392
rect 25752 20383 25780 20389
rect 25752 20349 25764 20383
rect 25752 20343 25780 20349
rect 25774 20340 25780 20343
rect 25832 20340 25838 20392
rect 26973 20383 27031 20389
rect 26973 20349 26985 20383
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 22066 20284 23244 20312
rect 20901 20275 20959 20281
rect 26142 20272 26148 20324
rect 26200 20272 26206 20324
rect 26988 20256 27016 20343
rect 28902 20340 28908 20392
rect 28960 20340 28966 20392
rect 28994 20340 29000 20392
rect 29052 20340 29058 20392
rect 31036 20380 31064 20420
rect 31113 20417 31125 20451
rect 31159 20417 31171 20451
rect 31113 20411 31171 20417
rect 31478 20408 31484 20460
rect 31536 20408 31542 20460
rect 31662 20448 31668 20460
rect 31588 20420 31668 20448
rect 31389 20383 31447 20389
rect 31389 20380 31401 20383
rect 31036 20352 31401 20380
rect 31389 20349 31401 20352
rect 31435 20380 31447 20383
rect 31588 20380 31616 20420
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 32950 20408 32956 20460
rect 33008 20408 33014 20460
rect 33778 20408 33784 20460
rect 33836 20448 33842 20460
rect 33965 20451 34023 20457
rect 33965 20448 33977 20451
rect 33836 20420 33977 20448
rect 33836 20408 33842 20420
rect 33965 20417 33977 20420
rect 34011 20417 34023 20451
rect 33965 20411 34023 20417
rect 34146 20408 34152 20460
rect 34204 20408 34210 20460
rect 34609 20451 34667 20457
rect 34609 20448 34621 20451
rect 34256 20420 34621 20448
rect 33091 20383 33149 20389
rect 33091 20380 33103 20383
rect 31435 20352 31616 20380
rect 31726 20352 33103 20380
rect 31435 20349 31447 20352
rect 31389 20343 31447 20349
rect 28166 20272 28172 20324
rect 28224 20312 28230 20324
rect 29012 20312 29040 20340
rect 28224 20284 29040 20312
rect 28224 20272 28230 20284
rect 31570 20272 31576 20324
rect 31628 20312 31634 20324
rect 31726 20312 31754 20352
rect 33091 20349 33103 20352
rect 33137 20349 33149 20383
rect 33091 20343 33149 20349
rect 33226 20340 33232 20392
rect 33284 20340 33290 20392
rect 33502 20340 33508 20392
rect 33560 20380 33566 20392
rect 33870 20380 33876 20392
rect 33560 20352 33876 20380
rect 33560 20340 33566 20352
rect 33870 20340 33876 20352
rect 33928 20340 33934 20392
rect 31628 20284 31754 20312
rect 31628 20272 31634 20284
rect 33594 20272 33600 20324
rect 33652 20312 33658 20324
rect 34256 20312 34284 20420
rect 34609 20417 34621 20420
rect 34655 20417 34667 20451
rect 34609 20411 34667 20417
rect 34698 20408 34704 20460
rect 34756 20408 34762 20460
rect 35710 20408 35716 20460
rect 35768 20408 35774 20460
rect 35986 20457 35992 20460
rect 35980 20448 35992 20457
rect 35947 20420 35992 20448
rect 35980 20411 35992 20420
rect 35986 20408 35992 20411
rect 36044 20408 36050 20460
rect 34425 20383 34483 20389
rect 34425 20349 34437 20383
rect 34471 20349 34483 20383
rect 34425 20343 34483 20349
rect 34517 20383 34575 20389
rect 34517 20349 34529 20383
rect 34563 20380 34575 20383
rect 34716 20380 34744 20408
rect 34563 20352 34744 20380
rect 37660 20380 37688 20544
rect 42702 20525 42708 20528
rect 42696 20516 42708 20525
rect 42663 20488 42708 20516
rect 42696 20479 42708 20488
rect 42702 20476 42708 20479
rect 42760 20476 42766 20528
rect 43070 20476 43076 20528
rect 43128 20516 43134 20528
rect 44284 20516 44312 20556
rect 46952 20528 46980 20556
rect 47305 20553 47317 20587
rect 47351 20584 47363 20587
rect 48222 20584 48228 20596
rect 47351 20556 48228 20584
rect 47351 20553 47363 20556
rect 47305 20547 47363 20553
rect 48222 20544 48228 20556
rect 48280 20544 48286 20596
rect 51902 20584 51908 20596
rect 51046 20556 51908 20584
rect 43128 20488 44312 20516
rect 46192 20519 46250 20525
rect 43128 20476 43134 20488
rect 46192 20485 46204 20519
rect 46238 20516 46250 20519
rect 46750 20516 46756 20528
rect 46238 20488 46756 20516
rect 46238 20485 46250 20488
rect 46192 20479 46250 20485
rect 46750 20476 46756 20488
rect 46808 20476 46814 20528
rect 46934 20476 46940 20528
rect 46992 20476 46998 20528
rect 50648 20519 50706 20525
rect 50648 20485 50660 20519
rect 50694 20516 50706 20519
rect 50890 20516 50896 20528
rect 50694 20488 50896 20516
rect 50694 20485 50706 20488
rect 50648 20479 50706 20485
rect 50890 20476 50896 20488
rect 50948 20476 50954 20528
rect 38378 20408 38384 20460
rect 38436 20408 38442 20460
rect 39393 20451 39451 20457
rect 39393 20417 39405 20451
rect 39439 20448 39451 20451
rect 39850 20448 39856 20460
rect 39439 20420 39856 20448
rect 39439 20417 39451 20420
rect 39393 20411 39451 20417
rect 39850 20408 39856 20420
rect 39908 20408 39914 20460
rect 45738 20408 45744 20460
rect 45796 20448 45802 20460
rect 45833 20451 45891 20457
rect 45833 20448 45845 20451
rect 45796 20420 45845 20448
rect 45796 20408 45802 20420
rect 45833 20417 45845 20420
rect 45879 20417 45891 20451
rect 45833 20411 45891 20417
rect 48314 20408 48320 20460
rect 48372 20457 48378 20460
rect 48372 20451 48421 20457
rect 48372 20417 48375 20451
rect 48409 20417 48421 20451
rect 48372 20411 48421 20417
rect 48372 20408 48378 20411
rect 49418 20408 49424 20460
rect 49476 20408 49482 20460
rect 38519 20383 38577 20389
rect 38519 20380 38531 20383
rect 37660 20352 38531 20380
rect 34563 20349 34575 20352
rect 34517 20343 34575 20349
rect 38519 20349 38531 20352
rect 38565 20349 38577 20383
rect 38519 20343 38577 20349
rect 33652 20284 34284 20312
rect 34440 20312 34468 20343
rect 38654 20340 38660 20392
rect 38712 20340 38718 20392
rect 38838 20340 38844 20392
rect 38896 20380 38902 20392
rect 38933 20383 38991 20389
rect 38933 20380 38945 20383
rect 38896 20352 38945 20380
rect 38896 20340 38902 20352
rect 38933 20349 38945 20352
rect 38979 20349 38991 20383
rect 38933 20343 38991 20349
rect 39577 20383 39635 20389
rect 39577 20349 39589 20383
rect 39623 20349 39635 20383
rect 39577 20343 39635 20349
rect 35253 20315 35311 20321
rect 35253 20312 35265 20315
rect 34440 20284 35265 20312
rect 33652 20272 33658 20284
rect 35253 20281 35265 20284
rect 35299 20312 35311 20315
rect 35526 20312 35532 20324
rect 35299 20284 35532 20312
rect 35299 20281 35311 20284
rect 35253 20275 35311 20281
rect 35526 20272 35532 20284
rect 35584 20272 35590 20324
rect 39592 20256 39620 20343
rect 39758 20340 39764 20392
rect 39816 20380 39822 20392
rect 40034 20380 40040 20392
rect 39816 20352 40040 20380
rect 39816 20340 39822 20352
rect 40034 20340 40040 20352
rect 40092 20340 40098 20392
rect 42426 20340 42432 20392
rect 42484 20340 42490 20392
rect 45922 20340 45928 20392
rect 45980 20340 45986 20392
rect 48225 20383 48283 20389
rect 48225 20380 48237 20383
rect 47688 20352 48237 20380
rect 16114 20244 16120 20256
rect 14568 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 19705 20247 19763 20253
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 21358 20244 21364 20256
rect 19751 20216 21364 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 26234 20244 26240 20256
rect 24995 20216 26240 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 26234 20204 26240 20216
rect 26292 20204 26298 20256
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 32309 20247 32367 20253
rect 32309 20213 32321 20247
rect 32355 20244 32367 20247
rect 34698 20244 34704 20256
rect 32355 20216 34704 20244
rect 32355 20213 32367 20216
rect 32309 20207 32367 20213
rect 34698 20204 34704 20216
rect 34756 20204 34762 20256
rect 34974 20204 34980 20256
rect 35032 20204 35038 20256
rect 37737 20247 37795 20253
rect 37737 20213 37749 20247
rect 37783 20244 37795 20247
rect 38838 20244 38844 20256
rect 37783 20216 38844 20244
rect 37783 20213 37795 20216
rect 37737 20207 37795 20213
rect 38838 20204 38844 20216
rect 38896 20204 38902 20256
rect 39574 20204 39580 20256
rect 39632 20204 39638 20256
rect 41417 20247 41475 20253
rect 41417 20213 41429 20247
rect 41463 20244 41475 20247
rect 42444 20244 42472 20340
rect 47688 20256 47716 20352
rect 48225 20349 48237 20352
rect 48271 20349 48283 20383
rect 48225 20343 48283 20349
rect 48501 20383 48559 20389
rect 48501 20349 48513 20383
rect 48547 20380 48559 20383
rect 49237 20383 49295 20389
rect 48547 20352 48728 20380
rect 48547 20349 48559 20352
rect 48501 20343 48559 20349
rect 44545 20247 44603 20253
rect 44545 20244 44557 20247
rect 41463 20216 44557 20244
rect 41463 20213 41475 20216
rect 41417 20207 41475 20213
rect 44545 20213 44557 20216
rect 44591 20244 44603 20247
rect 45002 20244 45008 20256
rect 44591 20216 45008 20244
rect 44591 20213 44603 20216
rect 44545 20207 44603 20213
rect 45002 20204 45008 20216
rect 45060 20204 45066 20256
rect 47578 20204 47584 20256
rect 47636 20204 47642 20256
rect 47670 20204 47676 20256
rect 47728 20204 47734 20256
rect 47762 20204 47768 20256
rect 47820 20244 47826 20256
rect 48700 20244 48728 20352
rect 49237 20349 49249 20383
rect 49283 20349 49295 20383
rect 49237 20343 49295 20349
rect 50893 20383 50951 20389
rect 50893 20349 50905 20383
rect 50939 20380 50951 20383
rect 51046 20380 51074 20556
rect 51902 20544 51908 20556
rect 51960 20584 51966 20596
rect 57149 20587 57207 20593
rect 51960 20556 55536 20584
rect 51960 20544 51966 20556
rect 51436 20519 51494 20525
rect 51436 20485 51448 20519
rect 51482 20516 51494 20519
rect 53006 20516 53012 20528
rect 51482 20488 53012 20516
rect 51482 20485 51494 20488
rect 51436 20479 51494 20485
rect 53006 20476 53012 20488
rect 53064 20476 53070 20528
rect 53101 20519 53159 20525
rect 53101 20485 53113 20519
rect 53147 20516 53159 20519
rect 53742 20516 53748 20528
rect 53147 20488 53748 20516
rect 53147 20485 53159 20488
rect 53101 20479 53159 20485
rect 53742 20476 53748 20488
rect 53800 20476 53806 20528
rect 52546 20408 52552 20460
rect 52604 20448 52610 20460
rect 54662 20457 54668 20460
rect 54640 20451 54668 20457
rect 52604 20420 53052 20448
rect 52604 20408 52610 20420
rect 53024 20392 53052 20420
rect 54640 20417 54652 20451
rect 54640 20411 54668 20417
rect 54662 20408 54668 20411
rect 54720 20408 54726 20460
rect 55508 20448 55536 20556
rect 57149 20553 57161 20587
rect 57195 20584 57207 20587
rect 57514 20584 57520 20596
rect 57195 20556 57520 20584
rect 57195 20553 57207 20556
rect 57149 20547 57207 20553
rect 56042 20525 56048 20528
rect 56036 20516 56048 20525
rect 56003 20488 56048 20516
rect 56036 20479 56048 20488
rect 56042 20476 56048 20479
rect 56100 20476 56106 20528
rect 55769 20451 55827 20457
rect 55769 20448 55781 20451
rect 55416 20420 55781 20448
rect 55416 20392 55444 20420
rect 55769 20417 55781 20420
rect 55815 20417 55827 20451
rect 57164 20448 57192 20547
rect 57514 20544 57520 20556
rect 57572 20544 57578 20596
rect 55769 20411 55827 20417
rect 55876 20420 57192 20448
rect 51169 20383 51227 20389
rect 51169 20380 51181 20383
rect 50939 20352 51181 20380
rect 50939 20349 50951 20352
rect 50893 20343 50951 20349
rect 51169 20349 51181 20352
rect 51215 20349 51227 20383
rect 51169 20343 51227 20349
rect 48777 20315 48835 20321
rect 48777 20281 48789 20315
rect 48823 20312 48835 20315
rect 48866 20312 48872 20324
rect 48823 20284 48872 20312
rect 48823 20281 48835 20284
rect 48777 20275 48835 20281
rect 48866 20272 48872 20284
rect 48924 20272 48930 20324
rect 49252 20312 49280 20343
rect 52822 20340 52828 20392
rect 52880 20340 52886 20392
rect 53006 20340 53012 20392
rect 53064 20340 53070 20392
rect 53834 20380 53840 20392
rect 53392 20352 53840 20380
rect 52549 20315 52607 20321
rect 49252 20284 49556 20312
rect 49528 20253 49556 20284
rect 52549 20281 52561 20315
rect 52595 20312 52607 20315
rect 53392 20312 53420 20352
rect 53834 20340 53840 20352
rect 53892 20340 53898 20392
rect 54478 20340 54484 20392
rect 54536 20340 54542 20392
rect 54754 20340 54760 20392
rect 54812 20340 54818 20392
rect 55398 20340 55404 20392
rect 55456 20340 55462 20392
rect 55490 20340 55496 20392
rect 55548 20340 55554 20392
rect 55677 20383 55735 20389
rect 55677 20349 55689 20383
rect 55723 20380 55735 20383
rect 55876 20380 55904 20420
rect 55723 20352 55904 20380
rect 55723 20349 55735 20352
rect 55677 20343 55735 20349
rect 52595 20284 53420 20312
rect 52595 20281 52607 20284
rect 52549 20275 52607 20281
rect 53466 20272 53472 20324
rect 53524 20272 53530 20324
rect 54938 20272 54944 20324
rect 54996 20312 55002 20324
rect 55033 20315 55091 20321
rect 55033 20312 55045 20315
rect 54996 20284 55045 20312
rect 54996 20272 55002 20284
rect 55033 20281 55045 20284
rect 55079 20281 55091 20315
rect 55033 20275 55091 20281
rect 47820 20216 48728 20244
rect 49513 20247 49571 20253
rect 47820 20204 47826 20216
rect 49513 20213 49525 20247
rect 49559 20244 49571 20247
rect 50706 20244 50712 20256
rect 49559 20216 50712 20244
rect 49559 20213 49571 20216
rect 49513 20207 49571 20213
rect 50706 20204 50712 20216
rect 50764 20204 50770 20256
rect 53837 20247 53895 20253
rect 53837 20213 53849 20247
rect 53883 20244 53895 20247
rect 55766 20244 55772 20256
rect 53883 20216 55772 20244
rect 53883 20213 53895 20216
rect 53837 20207 53895 20213
rect 55766 20204 55772 20216
rect 55824 20204 55830 20256
rect 1104 20154 58880 20176
rect 1104 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 22616 20154
rect 22668 20102 22680 20154
rect 22732 20102 22744 20154
rect 22796 20102 22808 20154
rect 22860 20102 22872 20154
rect 22924 20102 37060 20154
rect 37112 20102 37124 20154
rect 37176 20102 37188 20154
rect 37240 20102 37252 20154
rect 37304 20102 37316 20154
rect 37368 20102 51504 20154
rect 51556 20102 51568 20154
rect 51620 20102 51632 20154
rect 51684 20102 51696 20154
rect 51748 20102 51760 20154
rect 51812 20102 58880 20154
rect 1104 20080 58880 20102
rect 5626 20000 5632 20052
rect 5684 20000 5690 20052
rect 7650 20040 7656 20052
rect 6472 20012 7656 20040
rect 5537 19975 5595 19981
rect 5537 19941 5549 19975
rect 5583 19972 5595 19975
rect 6472 19972 6500 20012
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8665 20043 8723 20049
rect 8665 20009 8677 20043
rect 8711 20040 8723 20043
rect 8754 20040 8760 20052
rect 8711 20012 8760 20040
rect 8711 20009 8723 20012
rect 8665 20003 8723 20009
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 10192 20012 10517 20040
rect 10192 20000 10198 20012
rect 10505 20009 10517 20012
rect 10551 20009 10563 20043
rect 10505 20003 10563 20009
rect 12253 20043 12311 20049
rect 12253 20009 12265 20043
rect 12299 20040 12311 20043
rect 12802 20040 12808 20052
rect 12299 20012 12808 20040
rect 12299 20009 12311 20012
rect 12253 20003 12311 20009
rect 12802 20000 12808 20012
rect 12860 20040 12866 20052
rect 13630 20040 13636 20052
rect 12860 20012 13636 20040
rect 12860 20000 12866 20012
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14090 20000 14096 20052
rect 14148 20000 14154 20052
rect 15746 20040 15752 20052
rect 14568 20012 15752 20040
rect 5583 19944 6500 19972
rect 5583 19941 5595 19944
rect 5537 19935 5595 19941
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4246 19836 4252 19848
rect 4203 19808 4252 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4246 19796 4252 19808
rect 4304 19836 4310 19848
rect 6273 19839 6331 19845
rect 4304 19808 6224 19836
rect 4304 19796 4310 19808
rect 4430 19777 4436 19780
rect 4424 19768 4436 19777
rect 4391 19740 4436 19768
rect 4424 19731 4436 19740
rect 4430 19728 4436 19731
rect 4488 19728 4494 19780
rect 6196 19768 6224 19808
rect 6273 19805 6285 19839
rect 6319 19836 6331 19839
rect 6472 19836 6500 19944
rect 9677 19975 9735 19981
rect 9677 19941 9689 19975
rect 9723 19941 9735 19975
rect 9677 19935 9735 19941
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19873 7343 19907
rect 7285 19867 7343 19873
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19873 9183 19907
rect 9692 19904 9720 19935
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 12989 19975 13047 19981
rect 12989 19972 13001 19975
rect 12124 19944 13001 19972
rect 12124 19932 12130 19944
rect 12989 19941 13001 19944
rect 13035 19972 13047 19975
rect 14568 19972 14596 20012
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 18288 20012 19257 20040
rect 18288 20000 18294 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 20622 20040 20628 20052
rect 19245 20003 19303 20009
rect 19996 20012 20628 20040
rect 13035 19944 14596 19972
rect 18509 19975 18567 19981
rect 13035 19941 13047 19944
rect 12989 19935 13047 19941
rect 18509 19941 18521 19975
rect 18555 19972 18567 19975
rect 19996 19972 20024 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21726 20000 21732 20052
rect 21784 20000 21790 20052
rect 23566 20000 23572 20052
rect 23624 20000 23630 20052
rect 25038 20000 25044 20052
rect 25096 20040 25102 20052
rect 25225 20043 25283 20049
rect 25225 20040 25237 20043
rect 25096 20012 25237 20040
rect 25096 20000 25102 20012
rect 25225 20009 25237 20012
rect 25271 20009 25283 20043
rect 25225 20003 25283 20009
rect 27706 20000 27712 20052
rect 27764 20000 27770 20052
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 28997 20043 29055 20049
rect 28997 20040 29009 20043
rect 28960 20012 29009 20040
rect 28960 20000 28966 20012
rect 28997 20009 29009 20012
rect 29043 20009 29055 20043
rect 28997 20003 29055 20009
rect 30834 20000 30840 20052
rect 30892 20040 30898 20052
rect 31205 20043 31263 20049
rect 31205 20040 31217 20043
rect 30892 20012 31217 20040
rect 30892 20000 30898 20012
rect 31205 20009 31217 20012
rect 31251 20009 31263 20043
rect 33226 20040 33232 20052
rect 31205 20003 31263 20009
rect 31726 20012 33232 20040
rect 18555 19944 20024 19972
rect 18555 19941 18567 19944
rect 18509 19935 18567 19941
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9692 19876 9873 19904
rect 9125 19867 9183 19873
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 12434 19904 12440 19916
rect 9861 19867 9919 19873
rect 11900 19876 12440 19904
rect 6319 19808 6500 19836
rect 6319 19805 6331 19808
rect 6273 19799 6331 19805
rect 7300 19780 7328 19867
rect 7282 19768 7288 19780
rect 6196 19740 7288 19768
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 7552 19771 7610 19777
rect 7552 19737 7564 19771
rect 7598 19768 7610 19771
rect 7650 19768 7656 19780
rect 7598 19740 7656 19768
rect 7598 19737 7610 19740
rect 7552 19731 7610 19737
rect 7650 19728 7656 19740
rect 7708 19728 7714 19780
rect 9140 19768 9168 19867
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9766 19836 9772 19848
rect 9355 19808 9772 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 11900 19836 11928 19876
rect 12434 19864 12440 19876
rect 12492 19904 12498 19916
rect 17126 19904 17132 19916
rect 12492 19876 12664 19904
rect 12492 19864 12498 19876
rect 10928 19808 11928 19836
rect 12636 19836 12664 19876
rect 15948 19876 17132 19904
rect 15948 19848 15976 19876
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 12636 19808 15485 19836
rect 10928 19796 10934 19808
rect 15473 19805 15485 19808
rect 15519 19836 15531 19839
rect 15930 19836 15936 19848
rect 15519 19808 15936 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16114 19796 16120 19848
rect 16172 19796 16178 19848
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 19996 19836 20024 19944
rect 20349 19907 20407 19913
rect 20349 19904 20361 19907
rect 20088 19876 20361 19904
rect 20088 19848 20116 19876
rect 20349 19873 20361 19876
rect 20395 19873 20407 19907
rect 20349 19867 20407 19873
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21913 19907 21971 19913
rect 21913 19904 21925 19907
rect 21508 19876 21925 19904
rect 21508 19864 21514 19876
rect 21913 19873 21925 19876
rect 21959 19873 21971 19907
rect 23750 19904 23756 19916
rect 21913 19867 21971 19873
rect 23492 19876 23756 19904
rect 19935 19808 20024 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 20616 19839 20674 19845
rect 20616 19805 20628 19839
rect 20662 19836 20674 19839
rect 21542 19836 21548 19848
rect 20662 19808 21548 19836
rect 20662 19805 20674 19808
rect 20616 19799 20674 19805
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 23492 19845 23520 19876
rect 23750 19864 23756 19876
rect 23808 19904 23814 19916
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 23808 19876 24961 19904
rect 23808 19864 23814 19876
rect 24949 19873 24961 19876
rect 24995 19873 25007 19907
rect 27724 19904 27752 20000
rect 31113 19975 31171 19981
rect 31113 19941 31125 19975
rect 31159 19972 31171 19975
rect 31726 19972 31754 20012
rect 33226 20000 33232 20012
rect 33284 20000 33290 20052
rect 33965 20043 34023 20049
rect 33965 20009 33977 20043
rect 34011 20040 34023 20043
rect 34146 20040 34152 20052
rect 34011 20012 34152 20040
rect 34011 20009 34023 20012
rect 33965 20003 34023 20009
rect 34146 20000 34152 20012
rect 34204 20000 34210 20052
rect 34606 20000 34612 20052
rect 34664 20040 34670 20052
rect 34701 20043 34759 20049
rect 34701 20040 34713 20043
rect 34664 20012 34713 20040
rect 34664 20000 34670 20012
rect 34701 20009 34713 20012
rect 34747 20009 34759 20043
rect 34701 20003 34759 20009
rect 37461 20043 37519 20049
rect 37461 20009 37473 20043
rect 37507 20040 37519 20043
rect 38654 20040 38660 20052
rect 37507 20012 38660 20040
rect 37507 20009 37519 20012
rect 37461 20003 37519 20009
rect 38654 20000 38660 20012
rect 38712 20000 38718 20052
rect 39022 20000 39028 20052
rect 39080 20040 39086 20052
rect 39853 20043 39911 20049
rect 39853 20040 39865 20043
rect 39080 20012 39865 20040
rect 39080 20000 39086 20012
rect 39853 20009 39865 20012
rect 39899 20009 39911 20043
rect 39853 20003 39911 20009
rect 42705 20043 42763 20049
rect 42705 20009 42717 20043
rect 42751 20040 42763 20043
rect 43254 20040 43260 20052
rect 42751 20012 43260 20040
rect 42751 20009 42763 20012
rect 42705 20003 42763 20009
rect 43254 20000 43260 20012
rect 43312 20000 43318 20052
rect 43901 20043 43959 20049
rect 43901 20009 43913 20043
rect 43947 20040 43959 20043
rect 43990 20040 43996 20052
rect 43947 20012 43996 20040
rect 43947 20009 43959 20012
rect 43901 20003 43959 20009
rect 43990 20000 43996 20012
rect 44048 20000 44054 20052
rect 46753 20043 46811 20049
rect 46753 20009 46765 20043
rect 46799 20040 46811 20043
rect 47762 20040 47768 20052
rect 46799 20012 47768 20040
rect 46799 20009 46811 20012
rect 46753 20003 46811 20009
rect 47762 20000 47768 20012
rect 47820 20000 47826 20052
rect 49050 20040 49056 20052
rect 48148 20012 49056 20040
rect 39393 19975 39451 19981
rect 31159 19944 31800 19972
rect 31159 19941 31171 19944
rect 31113 19935 31171 19941
rect 31772 19913 31800 19944
rect 39393 19941 39405 19975
rect 39439 19941 39451 19975
rect 39393 19935 39451 19941
rect 42153 19975 42211 19981
rect 42153 19941 42165 19975
rect 42199 19972 42211 19975
rect 42199 19944 43668 19972
rect 42199 19941 42211 19944
rect 42153 19935 42211 19941
rect 28353 19907 28411 19913
rect 28353 19904 28365 19907
rect 27724 19876 28365 19904
rect 24949 19867 25007 19873
rect 28353 19873 28365 19876
rect 28399 19873 28411 19907
rect 28353 19867 28411 19873
rect 31757 19907 31815 19913
rect 31757 19873 31769 19907
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 35710 19864 35716 19916
rect 35768 19904 35774 19916
rect 36081 19907 36139 19913
rect 36081 19904 36093 19907
rect 35768 19876 36093 19904
rect 35768 19864 35774 19876
rect 36081 19873 36093 19876
rect 36127 19873 36139 19907
rect 39408 19904 39436 19935
rect 43640 19916 43668 19944
rect 43714 19932 43720 19984
rect 43772 19972 43778 19984
rect 43772 19944 44588 19972
rect 43772 19932 43778 19944
rect 39574 19904 39580 19916
rect 39408 19876 39580 19904
rect 36081 19867 36139 19873
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19805 23535 19839
rect 23477 19799 23535 19805
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19836 24271 19839
rect 25777 19839 25835 19845
rect 24259 19808 24440 19836
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 11140 19771 11198 19777
rect 9140 19740 9904 19768
rect 9876 19712 9904 19740
rect 11140 19737 11152 19771
rect 11186 19768 11198 19771
rect 11514 19768 11520 19780
rect 11186 19740 11520 19768
rect 11186 19737 11198 19740
rect 11140 19731 11198 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 12618 19728 12624 19780
rect 12676 19768 12682 19780
rect 13354 19768 13360 19780
rect 12676 19740 13360 19768
rect 12676 19728 12682 19740
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 15228 19771 15286 19777
rect 15228 19737 15240 19771
rect 15274 19768 15286 19771
rect 15746 19768 15752 19780
rect 15274 19740 15752 19768
rect 15274 19737 15286 19740
rect 15228 19731 15286 19737
rect 15746 19728 15752 19740
rect 15804 19728 15810 19780
rect 17396 19771 17454 19777
rect 17396 19737 17408 19771
rect 17442 19768 17454 19771
rect 17586 19768 17592 19780
rect 17442 19740 17592 19768
rect 17442 19737 17454 19740
rect 17396 19731 17454 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 19061 19771 19119 19777
rect 19061 19737 19073 19771
rect 19107 19768 19119 19771
rect 19107 19740 20760 19768
rect 19107 19737 19119 19740
rect 19061 19731 19119 19737
rect 20732 19712 20760 19740
rect 9122 19660 9128 19712
rect 9180 19700 9186 19712
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 9180 19672 9229 19700
rect 9180 19660 9186 19672
rect 9217 19669 9229 19672
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 9858 19660 9864 19712
rect 9916 19660 9922 19712
rect 12526 19660 12532 19712
rect 12584 19660 12590 19712
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 15565 19703 15623 19709
rect 15565 19700 15577 19703
rect 14608 19672 15577 19700
rect 14608 19660 14614 19672
rect 15565 19669 15577 19672
rect 15611 19669 15623 19703
rect 15565 19663 15623 19669
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20165 19703 20223 19709
rect 20165 19700 20177 19703
rect 19944 19672 20177 19700
rect 19944 19660 19950 19672
rect 20165 19669 20177 19672
rect 20211 19700 20223 19703
rect 20346 19700 20352 19712
rect 20211 19672 20352 19700
rect 20211 19669 20223 19672
rect 20165 19663 20223 19669
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 20714 19660 20720 19712
rect 20772 19660 20778 19712
rect 22554 19660 22560 19712
rect 22612 19660 22618 19712
rect 24412 19709 24440 19808
rect 25777 19805 25789 19839
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26596 19839 26654 19845
rect 26596 19805 26608 19839
rect 26642 19836 26654 19839
rect 28074 19836 28080 19848
rect 26642 19808 28080 19836
rect 26642 19805 26654 19808
rect 26596 19799 26654 19805
rect 24857 19771 24915 19777
rect 24857 19737 24869 19771
rect 24903 19768 24915 19771
rect 25222 19768 25228 19780
rect 24903 19740 25228 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 25792 19712 25820 19799
rect 26344 19768 26372 19799
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 29638 19796 29644 19848
rect 29696 19796 29702 19848
rect 29730 19796 29736 19848
rect 29788 19796 29794 19848
rect 32585 19839 32643 19845
rect 32585 19836 32597 19839
rect 32140 19808 32597 19836
rect 26970 19768 26976 19780
rect 26344 19740 26976 19768
rect 26970 19728 26976 19740
rect 27028 19728 27034 19780
rect 29656 19768 29684 19796
rect 29978 19771 30036 19777
rect 29978 19768 29990 19771
rect 29656 19740 29990 19768
rect 29978 19737 29990 19740
rect 30024 19737 30036 19771
rect 29978 19731 30036 19737
rect 32140 19712 32168 19808
rect 32585 19805 32597 19808
rect 32631 19805 32643 19839
rect 32585 19799 32643 19805
rect 35250 19796 35256 19848
rect 35308 19796 35314 19848
rect 35526 19796 35532 19848
rect 35584 19796 35590 19848
rect 36096 19836 36124 19867
rect 39574 19864 39580 19876
rect 39632 19904 39638 19916
rect 40405 19907 40463 19913
rect 40405 19904 40417 19907
rect 39632 19876 40417 19904
rect 39632 19864 39638 19876
rect 40405 19873 40417 19876
rect 40451 19873 40463 19907
rect 40405 19867 40463 19873
rect 40494 19864 40500 19916
rect 40552 19904 40558 19916
rect 41785 19907 41843 19913
rect 41785 19904 41797 19907
rect 40552 19876 41797 19904
rect 40552 19864 40558 19876
rect 41785 19873 41797 19876
rect 41831 19904 41843 19907
rect 43346 19904 43352 19916
rect 41831 19876 43352 19904
rect 41831 19873 41843 19876
rect 41785 19867 41843 19873
rect 43346 19864 43352 19876
rect 43404 19864 43410 19916
rect 43622 19864 43628 19916
rect 43680 19864 43686 19916
rect 43806 19864 43812 19916
rect 43864 19864 43870 19916
rect 44560 19913 44588 19944
rect 47578 19932 47584 19984
rect 47636 19972 47642 19984
rect 48148 19972 48176 20012
rect 49050 20000 49056 20012
rect 49108 20000 49114 20052
rect 49418 20000 49424 20052
rect 49476 20040 49482 20052
rect 49513 20043 49571 20049
rect 49513 20040 49525 20043
rect 49476 20012 49525 20040
rect 49476 20000 49482 20012
rect 49513 20009 49525 20012
rect 49559 20009 49571 20043
rect 49513 20003 49571 20009
rect 51445 20043 51503 20049
rect 51445 20009 51457 20043
rect 51491 20040 51503 20043
rect 51902 20040 51908 20052
rect 51491 20012 51908 20040
rect 51491 20009 51503 20012
rect 51445 20003 51503 20009
rect 47636 19944 48176 19972
rect 47636 19932 47642 19944
rect 44545 19907 44603 19913
rect 44545 19873 44557 19907
rect 44591 19904 44603 19907
rect 44634 19904 44640 19916
rect 44591 19876 44640 19904
rect 44591 19873 44603 19876
rect 44545 19867 44603 19873
rect 44634 19864 44640 19876
rect 44692 19864 44698 19916
rect 47486 19864 47492 19916
rect 47544 19864 47550 19916
rect 50706 19864 50712 19916
rect 50764 19864 50770 19916
rect 51552 19913 51580 20012
rect 51902 20000 51908 20012
rect 51960 20000 51966 20052
rect 52822 20000 52828 20052
rect 52880 20040 52886 20052
rect 53929 20043 53987 20049
rect 53929 20040 53941 20043
rect 52880 20012 53941 20040
rect 52880 20000 52886 20012
rect 53929 20009 53941 20012
rect 53975 20009 53987 20043
rect 53929 20003 53987 20009
rect 55490 20000 55496 20052
rect 55548 20040 55554 20052
rect 56689 20043 56747 20049
rect 56689 20040 56701 20043
rect 55548 20012 56701 20040
rect 55548 20000 55554 20012
rect 56689 20009 56701 20012
rect 56735 20009 56747 20043
rect 56689 20003 56747 20009
rect 53374 19932 53380 19984
rect 53432 19972 53438 19984
rect 54754 19972 54760 19984
rect 53432 19944 54760 19972
rect 53432 19932 53438 19944
rect 54754 19932 54760 19944
rect 54812 19932 54818 19984
rect 51537 19907 51595 19913
rect 51537 19873 51549 19907
rect 51583 19873 51595 19907
rect 51537 19867 51595 19873
rect 37737 19839 37795 19845
rect 37737 19836 37749 19839
rect 36096 19808 37749 19836
rect 37737 19805 37749 19808
rect 37783 19836 37795 19839
rect 38013 19839 38071 19845
rect 38013 19836 38025 19839
rect 37783 19808 38025 19836
rect 37783 19805 37795 19808
rect 37737 19799 37795 19805
rect 38013 19805 38025 19808
rect 38059 19836 38071 19839
rect 39666 19836 39672 19848
rect 38059 19808 39672 19836
rect 38059 19805 38071 19808
rect 38013 19799 38071 19805
rect 39666 19796 39672 19808
rect 39724 19796 39730 19848
rect 32852 19771 32910 19777
rect 32852 19737 32864 19771
rect 32898 19768 32910 19771
rect 33502 19768 33508 19780
rect 32898 19740 33508 19768
rect 32898 19737 32910 19740
rect 32852 19731 32910 19737
rect 33502 19728 33508 19740
rect 33560 19728 33566 19780
rect 35544 19768 35572 19796
rect 36348 19771 36406 19777
rect 35544 19740 36308 19768
rect 24397 19703 24455 19709
rect 24397 19669 24409 19703
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 24762 19660 24768 19712
rect 24820 19660 24826 19712
rect 25774 19660 25780 19712
rect 25832 19660 25838 19712
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 34330 19660 34336 19712
rect 34388 19660 34394 19712
rect 35342 19660 35348 19712
rect 35400 19700 35406 19712
rect 35621 19703 35679 19709
rect 35621 19700 35633 19703
rect 35400 19672 35633 19700
rect 35400 19660 35406 19672
rect 35621 19669 35633 19672
rect 35667 19669 35679 19703
rect 36280 19700 36308 19740
rect 36348 19737 36360 19771
rect 36394 19768 36406 19771
rect 37274 19768 37280 19780
rect 36394 19740 37280 19768
rect 36394 19737 36406 19740
rect 36348 19731 36406 19737
rect 37274 19728 37280 19740
rect 37332 19728 37338 19780
rect 38280 19771 38338 19777
rect 38280 19737 38292 19771
rect 38326 19768 38338 19771
rect 38746 19768 38752 19780
rect 38326 19740 38752 19768
rect 38326 19737 38338 19740
rect 38280 19731 38338 19737
rect 38746 19728 38752 19740
rect 38804 19728 38810 19780
rect 39206 19700 39212 19712
rect 36280 19672 39212 19700
rect 35621 19663 35679 19669
rect 39206 19660 39212 19672
rect 39264 19700 39270 19712
rect 40512 19700 40540 19864
rect 42521 19839 42579 19845
rect 42521 19805 42533 19839
rect 42567 19836 42579 19839
rect 43070 19836 43076 19848
rect 42567 19808 43076 19836
rect 42567 19805 42579 19808
rect 42521 19799 42579 19805
rect 43070 19796 43076 19808
rect 43128 19796 43134 19848
rect 43165 19839 43223 19845
rect 43165 19805 43177 19839
rect 43211 19836 43223 19839
rect 43824 19836 43852 19864
rect 43211 19808 43852 19836
rect 44269 19839 44327 19845
rect 43211 19805 43223 19808
rect 43165 19799 43223 19805
rect 44269 19805 44281 19839
rect 44315 19836 44327 19839
rect 44818 19836 44824 19848
rect 44315 19808 44824 19836
rect 44315 19805 44327 19808
rect 44269 19799 44327 19805
rect 44818 19796 44824 19808
rect 44876 19796 44882 19848
rect 45002 19796 45008 19848
rect 45060 19836 45066 19848
rect 45281 19839 45339 19845
rect 45281 19836 45293 19839
rect 45060 19808 45293 19836
rect 45060 19796 45066 19808
rect 45281 19805 45293 19808
rect 45327 19836 45339 19839
rect 45373 19839 45431 19845
rect 45373 19836 45385 19839
rect 45327 19808 45385 19836
rect 45327 19805 45339 19808
rect 45281 19799 45339 19805
rect 45373 19805 45385 19808
rect 45419 19836 45431 19839
rect 45922 19836 45928 19848
rect 45419 19808 45928 19836
rect 45419 19805 45431 19808
rect 45373 19799 45431 19805
rect 45922 19796 45928 19808
rect 45980 19836 45986 19848
rect 47394 19836 47400 19848
rect 45980 19808 47400 19836
rect 45980 19796 45986 19808
rect 47394 19796 47400 19808
rect 47452 19836 47458 19848
rect 48133 19839 48191 19845
rect 48133 19836 48145 19839
rect 47452 19808 48145 19836
rect 47452 19796 47458 19808
rect 48133 19805 48145 19808
rect 48179 19836 48191 19839
rect 48958 19836 48964 19848
rect 48179 19808 48964 19836
rect 48179 19805 48191 19808
rect 48133 19799 48191 19805
rect 48958 19796 48964 19808
rect 49016 19836 49022 19848
rect 49789 19839 49847 19845
rect 49789 19836 49801 19839
rect 49016 19808 49801 19836
rect 49016 19796 49022 19808
rect 49789 19805 49801 19808
rect 49835 19836 49847 19839
rect 51552 19836 51580 19867
rect 52914 19864 52920 19916
rect 52972 19904 52978 19916
rect 53561 19907 53619 19913
rect 53561 19904 53573 19907
rect 52972 19876 53573 19904
rect 52972 19864 52978 19876
rect 53561 19873 53573 19876
rect 53607 19873 53619 19907
rect 56704 19904 56732 20003
rect 56778 20000 56784 20052
rect 56836 20000 56842 20052
rect 57333 19907 57391 19913
rect 57333 19904 57345 19907
rect 56704 19876 57345 19904
rect 53561 19867 53619 19873
rect 57333 19873 57345 19876
rect 57379 19873 57391 19907
rect 57333 19867 57391 19873
rect 49835 19808 51580 19836
rect 55125 19839 55183 19845
rect 49835 19805 49847 19808
rect 49789 19799 49847 19805
rect 55125 19805 55137 19839
rect 55171 19836 55183 19839
rect 55309 19839 55367 19845
rect 55309 19836 55321 19839
rect 55171 19808 55321 19836
rect 55171 19805 55183 19808
rect 55125 19799 55183 19805
rect 55309 19805 55321 19808
rect 55355 19836 55367 19839
rect 55398 19836 55404 19848
rect 55355 19808 55404 19836
rect 55355 19805 55367 19808
rect 55309 19799 55367 19805
rect 55398 19796 55404 19808
rect 55456 19796 55462 19848
rect 45640 19771 45698 19777
rect 45640 19737 45652 19771
rect 45686 19737 45698 19771
rect 45640 19731 45698 19737
rect 48400 19771 48458 19777
rect 48400 19737 48412 19771
rect 48446 19768 48458 19771
rect 48498 19768 48504 19780
rect 48446 19740 48504 19768
rect 48446 19737 48458 19740
rect 48400 19731 48458 19737
rect 39264 19672 40540 19700
rect 39264 19660 39270 19672
rect 42978 19660 42984 19712
rect 43036 19700 43042 19712
rect 43073 19703 43131 19709
rect 43073 19700 43085 19703
rect 43036 19672 43085 19700
rect 43036 19660 43042 19672
rect 43073 19669 43085 19672
rect 43119 19700 43131 19703
rect 44361 19703 44419 19709
rect 44361 19700 44373 19703
rect 43119 19672 44373 19700
rect 43119 19669 43131 19672
rect 43073 19663 43131 19669
rect 44361 19669 44373 19672
rect 44407 19669 44419 19703
rect 45664 19700 45692 19731
rect 48498 19728 48504 19740
rect 48556 19728 48562 19780
rect 51804 19771 51862 19777
rect 51804 19737 51816 19771
rect 51850 19768 51862 19771
rect 53009 19771 53067 19777
rect 53009 19768 53021 19771
rect 51850 19740 53021 19768
rect 51850 19737 51862 19740
rect 51804 19731 51862 19737
rect 53009 19737 53021 19740
rect 53055 19737 53067 19771
rect 53009 19731 53067 19737
rect 55576 19771 55634 19777
rect 55576 19737 55588 19771
rect 55622 19768 55634 19771
rect 55858 19768 55864 19780
rect 55622 19740 55864 19768
rect 55622 19737 55634 19740
rect 55576 19731 55634 19737
rect 55858 19728 55864 19740
rect 55916 19728 55922 19780
rect 46845 19703 46903 19709
rect 46845 19700 46857 19703
rect 45664 19672 46857 19700
rect 44361 19663 44419 19669
rect 46845 19669 46857 19672
rect 46891 19669 46903 19703
rect 46845 19663 46903 19669
rect 47857 19703 47915 19709
rect 47857 19669 47869 19703
rect 47903 19700 47915 19703
rect 48314 19700 48320 19712
rect 47903 19672 48320 19700
rect 47903 19669 47915 19672
rect 47857 19663 47915 19669
rect 48314 19660 48320 19672
rect 48372 19660 48378 19712
rect 50154 19660 50160 19712
rect 50212 19660 50218 19712
rect 52917 19703 52975 19709
rect 52917 19669 52929 19703
rect 52963 19700 52975 19703
rect 53374 19700 53380 19712
rect 52963 19672 53380 19700
rect 52963 19669 52975 19672
rect 52917 19663 52975 19669
rect 53374 19660 53380 19672
rect 53432 19660 53438 19712
rect 54294 19660 54300 19712
rect 54352 19700 54358 19712
rect 54938 19700 54944 19712
rect 54352 19672 54944 19700
rect 54352 19660 54358 19672
rect 54938 19660 54944 19672
rect 54996 19660 55002 19712
rect 1104 19610 59040 19632
rect 1104 19558 15394 19610
rect 15446 19558 15458 19610
rect 15510 19558 15522 19610
rect 15574 19558 15586 19610
rect 15638 19558 15650 19610
rect 15702 19558 29838 19610
rect 29890 19558 29902 19610
rect 29954 19558 29966 19610
rect 30018 19558 30030 19610
rect 30082 19558 30094 19610
rect 30146 19558 44282 19610
rect 44334 19558 44346 19610
rect 44398 19558 44410 19610
rect 44462 19558 44474 19610
rect 44526 19558 44538 19610
rect 44590 19558 58726 19610
rect 58778 19558 58790 19610
rect 58842 19558 58854 19610
rect 58906 19558 58918 19610
rect 58970 19558 58982 19610
rect 59034 19558 59040 19610
rect 1104 19536 59040 19558
rect 7650 19456 7656 19508
rect 7708 19456 7714 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10962 19496 10968 19508
rect 9916 19468 10968 19496
rect 9916 19456 9922 19468
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 14550 19456 14556 19508
rect 14608 19456 14614 19508
rect 15746 19456 15752 19508
rect 15804 19456 15810 19508
rect 17586 19456 17592 19508
rect 17644 19456 17650 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22554 19496 22560 19508
rect 22143 19468 22560 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 23658 19456 23664 19508
rect 23716 19456 23722 19508
rect 24857 19499 24915 19505
rect 24857 19465 24869 19499
rect 24903 19496 24915 19499
rect 25774 19496 25780 19508
rect 24903 19468 25780 19496
rect 24903 19465 24915 19468
rect 24857 19459 24915 19465
rect 25774 19456 25780 19468
rect 25832 19456 25838 19508
rect 33502 19456 33508 19508
rect 33560 19456 33566 19508
rect 33689 19499 33747 19505
rect 33689 19465 33701 19499
rect 33735 19496 33747 19499
rect 33962 19496 33968 19508
rect 33735 19468 33968 19496
rect 33735 19465 33747 19468
rect 33689 19459 33747 19465
rect 33962 19456 33968 19468
rect 34020 19456 34026 19508
rect 34057 19499 34115 19505
rect 34057 19465 34069 19499
rect 34103 19496 34115 19499
rect 35250 19496 35256 19508
rect 34103 19468 35256 19496
rect 34103 19465 34115 19468
rect 34057 19459 34115 19465
rect 35250 19456 35256 19468
rect 35308 19456 35314 19508
rect 37274 19456 37280 19508
rect 37332 19456 37338 19508
rect 38746 19456 38752 19508
rect 38804 19456 38810 19508
rect 39666 19456 39672 19508
rect 39724 19456 39730 19508
rect 43346 19456 43352 19508
rect 43404 19496 43410 19508
rect 48774 19496 48780 19508
rect 43404 19468 48780 19496
rect 43404 19456 43410 19468
rect 48774 19456 48780 19468
rect 48832 19456 48838 19508
rect 48958 19456 48964 19508
rect 49016 19456 49022 19508
rect 49513 19499 49571 19505
rect 49513 19465 49525 19499
rect 49559 19496 49571 19499
rect 50154 19496 50160 19508
rect 49559 19468 50160 19496
rect 49559 19465 49571 19468
rect 49513 19459 49571 19465
rect 50154 19456 50160 19468
rect 50212 19456 50218 19508
rect 55398 19456 55404 19508
rect 55456 19496 55462 19508
rect 55585 19499 55643 19505
rect 55585 19496 55597 19499
rect 55456 19468 55597 19496
rect 55456 19456 55462 19468
rect 55585 19465 55597 19468
rect 55631 19465 55643 19499
rect 55585 19459 55643 19465
rect 55858 19456 55864 19508
rect 55916 19456 55922 19508
rect 22189 19431 22247 19437
rect 22189 19397 22201 19431
rect 22235 19428 22247 19431
rect 22278 19428 22284 19440
rect 22235 19400 22284 19428
rect 22235 19397 22247 19400
rect 22189 19391 22247 19397
rect 22278 19388 22284 19400
rect 22336 19388 22342 19440
rect 22462 19388 22468 19440
rect 22520 19388 22526 19440
rect 7006 19320 7012 19372
rect 7064 19320 7070 19372
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 13722 19360 13728 19372
rect 12584 19332 13728 19360
rect 12584 19320 12590 19332
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14645 19363 14703 19369
rect 14645 19360 14657 19363
rect 14016 19332 14657 19360
rect 4154 19252 4160 19304
rect 4212 19252 4218 19304
rect 4614 19252 4620 19304
rect 4672 19252 4678 19304
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8297 19295 8355 19301
rect 8297 19292 8309 19295
rect 7800 19264 8309 19292
rect 7800 19252 7806 19264
rect 8297 19261 8309 19264
rect 8343 19261 8355 19295
rect 8297 19255 8355 19261
rect 8846 19252 8852 19304
rect 8904 19252 8910 19304
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 11330 19252 11336 19304
rect 11388 19292 11394 19304
rect 12069 19295 12127 19301
rect 12069 19292 12081 19295
rect 11388 19264 12081 19292
rect 11388 19252 11394 19264
rect 12069 19261 12081 19264
rect 12115 19261 12127 19295
rect 12069 19255 12127 19261
rect 12406 19264 13492 19292
rect 9398 19184 9404 19236
rect 9456 19224 9462 19236
rect 12406 19224 12434 19264
rect 9456 19196 12434 19224
rect 9456 19184 9462 19196
rect 3510 19116 3516 19168
rect 3568 19116 3574 19168
rect 5258 19116 5264 19168
rect 5316 19116 5322 19168
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 10686 19116 10692 19168
rect 10744 19116 10750 19168
rect 11514 19116 11520 19168
rect 11572 19116 11578 19168
rect 12894 19116 12900 19168
rect 12952 19116 12958 19168
rect 13464 19156 13492 19264
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 14016 19292 14044 19332
rect 14645 19329 14657 19332
rect 14691 19360 14703 19363
rect 14826 19360 14832 19372
rect 14691 19332 14832 19360
rect 14691 19329 14703 19332
rect 14645 19323 14703 19329
rect 14826 19320 14832 19332
rect 14884 19360 14890 19372
rect 21177 19363 21235 19369
rect 14884 19332 15240 19360
rect 14884 19320 14890 19332
rect 13596 19264 14044 19292
rect 14461 19295 14519 19301
rect 13596 19252 13602 19264
rect 14461 19261 14473 19295
rect 14507 19292 14519 19295
rect 15105 19295 15163 19301
rect 14507 19264 14872 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 14182 19224 14188 19236
rect 13832 19196 14188 19224
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13464 19128 13645 19156
rect 13633 19125 13645 19128
rect 13679 19156 13691 19159
rect 13832 19156 13860 19196
rect 14182 19184 14188 19196
rect 14240 19224 14246 19236
rect 14476 19224 14504 19255
rect 14240 19196 14504 19224
rect 14240 19184 14246 19196
rect 13679 19128 13860 19156
rect 13679 19125 13691 19128
rect 13633 19119 13691 19125
rect 13906 19116 13912 19168
rect 13964 19116 13970 19168
rect 14844 19156 14872 19264
rect 15105 19261 15117 19295
rect 15151 19261 15163 19295
rect 15212 19292 15240 19332
rect 21177 19329 21189 19363
rect 21223 19329 21235 19363
rect 22480 19360 22508 19388
rect 23676 19360 23704 19456
rect 33520 19428 33548 19456
rect 34149 19431 34207 19437
rect 34149 19428 34161 19431
rect 33520 19400 34161 19428
rect 34149 19397 34161 19400
rect 34195 19397 34207 19431
rect 34149 19391 34207 19397
rect 44634 19388 44640 19440
rect 44692 19428 44698 19440
rect 49421 19431 49479 19437
rect 44692 19400 49280 19428
rect 44692 19388 44698 19400
rect 23733 19363 23791 19369
rect 23733 19360 23745 19363
rect 22480 19332 22600 19360
rect 23676 19332 23745 19360
rect 21177 19323 21235 19329
rect 15286 19292 15292 19304
rect 15212 19264 15292 19292
rect 15105 19255 15163 19261
rect 15013 19227 15071 19233
rect 15013 19193 15025 19227
rect 15059 19224 15071 19227
rect 15120 19224 15148 19255
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17828 19264 18153 19292
rect 17828 19252 17834 19264
rect 18141 19261 18153 19264
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 21192 19292 21220 19323
rect 19392 19264 21220 19292
rect 22005 19295 22063 19301
rect 19392 19252 19398 19264
rect 22005 19261 22017 19295
rect 22051 19292 22063 19295
rect 22462 19292 22468 19304
rect 22051 19264 22468 19292
rect 22051 19261 22063 19264
rect 22005 19255 22063 19261
rect 15059 19196 15148 19224
rect 17144 19224 17172 19252
rect 19702 19224 19708 19236
rect 17144 19196 19708 19224
rect 15059 19193 15071 19196
rect 15013 19187 15071 19193
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 22020 19224 22048 19255
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 22572 19233 22600 19332
rect 23733 19329 23745 19332
rect 23779 19329 23791 19363
rect 23733 19323 23791 19329
rect 34793 19363 34851 19369
rect 34793 19329 34805 19363
rect 34839 19360 34851 19363
rect 34974 19360 34980 19372
rect 34839 19332 34980 19360
rect 34839 19329 34851 19332
rect 34793 19323 34851 19329
rect 34974 19320 34980 19332
rect 35032 19320 35038 19372
rect 40034 19360 40040 19372
rect 35866 19332 40040 19360
rect 23474 19252 23480 19304
rect 23532 19252 23538 19304
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 26142 19292 26148 19304
rect 25271 19264 26148 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 27982 19252 27988 19304
rect 28040 19252 28046 19304
rect 28534 19252 28540 19304
rect 28592 19292 28598 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28592 19264 28825 19292
rect 28592 19252 28598 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 31110 19252 31116 19304
rect 31168 19252 31174 19304
rect 32769 19295 32827 19301
rect 32769 19261 32781 19295
rect 32815 19261 32827 19295
rect 32769 19255 32827 19261
rect 33505 19295 33563 19301
rect 33505 19261 33517 19295
rect 33551 19261 33563 19295
rect 33505 19255 33563 19261
rect 19812 19196 22048 19224
rect 22557 19227 22615 19233
rect 19812 19156 19840 19196
rect 22557 19193 22569 19227
rect 22603 19193 22615 19227
rect 22557 19187 22615 19193
rect 22756 19196 23520 19224
rect 14844 19128 19840 19156
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 21232 19128 21465 19156
rect 21232 19116 21238 19128
rect 21453 19125 21465 19128
rect 21499 19156 21511 19159
rect 22756 19156 22784 19196
rect 21499 19128 22784 19156
rect 21499 19125 21511 19128
rect 21453 19119 21511 19125
rect 22830 19116 22836 19168
rect 22888 19156 22894 19168
rect 22925 19159 22983 19165
rect 22925 19156 22937 19159
rect 22888 19128 22937 19156
rect 22888 19116 22894 19128
rect 22925 19125 22937 19128
rect 22971 19156 22983 19159
rect 23382 19156 23388 19168
rect 22971 19128 23388 19156
rect 22971 19125 22983 19128
rect 22925 19119 22983 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 23492 19156 23520 19196
rect 32784 19168 32812 19255
rect 33520 19224 33548 19255
rect 33594 19252 33600 19304
rect 33652 19252 33658 19304
rect 34330 19252 34336 19304
rect 34388 19292 34394 19304
rect 35866 19292 35894 19332
rect 40034 19320 40040 19332
rect 40092 19320 40098 19372
rect 44082 19320 44088 19372
rect 44140 19320 44146 19372
rect 44174 19320 44180 19372
rect 44232 19360 44238 19372
rect 44269 19363 44327 19369
rect 44269 19360 44281 19363
rect 44232 19332 44281 19360
rect 44232 19320 44238 19332
rect 44269 19329 44281 19332
rect 44315 19329 44327 19363
rect 44269 19323 44327 19329
rect 45278 19320 45284 19372
rect 45336 19360 45342 19372
rect 45465 19363 45523 19369
rect 45465 19360 45477 19363
rect 45336 19332 45477 19360
rect 45336 19320 45342 19332
rect 45465 19329 45477 19332
rect 45511 19329 45523 19363
rect 45465 19323 45523 19329
rect 34388 19264 35894 19292
rect 37921 19295 37979 19301
rect 34388 19252 34394 19264
rect 37921 19261 37933 19295
rect 37967 19292 37979 19295
rect 38102 19292 38108 19304
rect 37967 19264 38108 19292
rect 37967 19261 37979 19264
rect 37921 19255 37979 19261
rect 38102 19252 38108 19264
rect 38160 19252 38166 19304
rect 38562 19252 38568 19304
rect 38620 19252 38626 19304
rect 38654 19252 38660 19304
rect 38712 19252 38718 19304
rect 39301 19295 39359 19301
rect 39301 19261 39313 19295
rect 39347 19261 39359 19295
rect 39301 19255 39359 19261
rect 34348 19224 34376 19252
rect 33520 19196 34376 19224
rect 38580 19224 38608 19252
rect 39316 19224 39344 19255
rect 42242 19252 42248 19304
rect 42300 19252 42306 19304
rect 42702 19252 42708 19304
rect 42760 19292 42766 19304
rect 43254 19301 43260 19304
rect 43073 19295 43131 19301
rect 43073 19292 43085 19295
rect 42760 19264 43085 19292
rect 42760 19252 42766 19264
rect 43073 19261 43085 19264
rect 43119 19261 43131 19295
rect 43073 19255 43131 19261
rect 43232 19295 43260 19301
rect 43232 19261 43244 19295
rect 43232 19255 43260 19261
rect 43254 19252 43260 19255
rect 43312 19252 43318 19304
rect 43349 19295 43407 19301
rect 43349 19261 43361 19295
rect 43395 19292 43407 19295
rect 43395 19264 43852 19292
rect 43395 19261 43407 19264
rect 43349 19255 43407 19261
rect 38580 19196 39344 19224
rect 41509 19227 41567 19233
rect 41509 19193 41521 19227
rect 41555 19224 41567 19227
rect 42720 19224 42748 19252
rect 41555 19196 42748 19224
rect 41555 19193 41567 19196
rect 41509 19187 41567 19193
rect 43622 19184 43628 19236
rect 43680 19184 43686 19236
rect 43824 19168 43852 19264
rect 46014 19252 46020 19304
rect 46072 19252 46078 19304
rect 47305 19295 47363 19301
rect 47305 19261 47317 19295
rect 47351 19292 47363 19295
rect 48314 19292 48320 19304
rect 47351 19264 48320 19292
rect 47351 19261 47363 19264
rect 47305 19255 47363 19261
rect 48314 19252 48320 19264
rect 48372 19292 48378 19304
rect 48774 19292 48780 19304
rect 48372 19264 48780 19292
rect 48372 19252 48378 19264
rect 48774 19252 48780 19264
rect 48832 19252 48838 19304
rect 49252 19301 49280 19400
rect 49421 19397 49433 19431
rect 49467 19397 49479 19431
rect 51258 19428 51264 19440
rect 49421 19391 49479 19397
rect 49896 19400 51264 19428
rect 49326 19320 49332 19372
rect 49384 19360 49390 19372
rect 49436 19360 49464 19391
rect 49384 19332 49464 19360
rect 49384 19320 49390 19332
rect 49237 19295 49295 19301
rect 49237 19261 49249 19295
rect 49283 19292 49295 19295
rect 49283 19264 49832 19292
rect 49283 19261 49295 19264
rect 49237 19255 49295 19261
rect 45738 19224 45744 19236
rect 44560 19196 45744 19224
rect 27246 19156 27252 19168
rect 23492 19128 27252 19156
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 27430 19116 27436 19168
rect 27488 19116 27494 19168
rect 28258 19116 28264 19168
rect 28316 19116 28322 19168
rect 30558 19116 30564 19168
rect 30616 19116 30622 19168
rect 31570 19116 31576 19168
rect 31628 19116 31634 19168
rect 31938 19116 31944 19168
rect 31996 19156 32002 19168
rect 32125 19159 32183 19165
rect 32125 19156 32137 19159
rect 31996 19128 32137 19156
rect 31996 19116 32002 19128
rect 32125 19125 32137 19128
rect 32171 19125 32183 19159
rect 32125 19119 32183 19125
rect 32766 19116 32772 19168
rect 32824 19116 32830 19168
rect 33134 19116 33140 19168
rect 33192 19116 33198 19168
rect 34882 19116 34888 19168
rect 34940 19156 34946 19168
rect 35069 19159 35127 19165
rect 35069 19156 35081 19159
rect 34940 19128 35081 19156
rect 34940 19116 34946 19128
rect 35069 19125 35081 19128
rect 35115 19125 35127 19159
rect 35069 19119 35127 19125
rect 36906 19116 36912 19168
rect 36964 19116 36970 19168
rect 38010 19116 38016 19168
rect 38068 19116 38074 19168
rect 41598 19116 41604 19168
rect 41656 19116 41662 19168
rect 42429 19159 42487 19165
rect 42429 19125 42441 19159
rect 42475 19156 42487 19159
rect 43714 19156 43720 19168
rect 42475 19128 43720 19156
rect 42475 19125 42487 19128
rect 42429 19119 42487 19125
rect 43714 19116 43720 19128
rect 43772 19116 43778 19168
rect 43806 19116 43812 19168
rect 43864 19116 43870 19168
rect 44174 19116 44180 19168
rect 44232 19156 44238 19168
rect 44560 19165 44588 19196
rect 45738 19184 45744 19196
rect 45796 19224 45802 19236
rect 49694 19224 49700 19236
rect 45796 19196 49700 19224
rect 45796 19184 45802 19196
rect 49694 19184 49700 19196
rect 49752 19184 49758 19236
rect 44545 19159 44603 19165
rect 44545 19156 44557 19159
rect 44232 19128 44557 19156
rect 44232 19116 44238 19128
rect 44545 19125 44557 19128
rect 44591 19125 44603 19159
rect 44545 19119 44603 19125
rect 44910 19116 44916 19168
rect 44968 19156 44974 19168
rect 46845 19159 46903 19165
rect 46845 19156 46857 19159
rect 44968 19128 46857 19156
rect 44968 19116 44974 19128
rect 46845 19125 46857 19128
rect 46891 19156 46903 19159
rect 47670 19156 47676 19168
rect 46891 19128 47676 19156
rect 46891 19125 46903 19128
rect 46845 19119 46903 19125
rect 47670 19116 47676 19128
rect 47728 19156 47734 19168
rect 47765 19159 47823 19165
rect 47765 19156 47777 19159
rect 47728 19128 47777 19156
rect 47728 19116 47734 19128
rect 47765 19125 47777 19128
rect 47811 19125 47823 19159
rect 47765 19119 47823 19125
rect 48222 19116 48228 19168
rect 48280 19116 48286 19168
rect 48590 19116 48596 19168
rect 48648 19116 48654 19168
rect 49804 19156 49832 19264
rect 49896 19233 49924 19400
rect 51258 19388 51264 19400
rect 51316 19388 51322 19440
rect 53469 19295 53527 19301
rect 53469 19292 53481 19295
rect 52564 19264 53481 19292
rect 49881 19227 49939 19233
rect 49881 19193 49893 19227
rect 49927 19193 49939 19227
rect 49881 19187 49939 19193
rect 52564 19168 52592 19264
rect 53469 19261 53481 19264
rect 53515 19261 53527 19295
rect 53469 19255 53527 19261
rect 56134 19252 56140 19304
rect 56192 19292 56198 19304
rect 56413 19295 56471 19301
rect 56413 19292 56425 19295
rect 56192 19264 56425 19292
rect 56192 19252 56198 19264
rect 56413 19261 56425 19264
rect 56459 19261 56471 19295
rect 56413 19255 56471 19261
rect 50157 19159 50215 19165
rect 50157 19156 50169 19159
rect 49804 19128 50169 19156
rect 50157 19125 50169 19128
rect 50203 19156 50215 19159
rect 51350 19156 51356 19168
rect 50203 19128 51356 19156
rect 50203 19125 50215 19128
rect 50157 19119 50215 19125
rect 51350 19116 51356 19128
rect 51408 19116 51414 19168
rect 52178 19116 52184 19168
rect 52236 19116 52242 19168
rect 52546 19116 52552 19168
rect 52604 19116 52610 19168
rect 52914 19116 52920 19168
rect 52972 19116 52978 19168
rect 1104 19066 58880 19088
rect 1104 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 22616 19066
rect 22668 19014 22680 19066
rect 22732 19014 22744 19066
rect 22796 19014 22808 19066
rect 22860 19014 22872 19066
rect 22924 19014 37060 19066
rect 37112 19014 37124 19066
rect 37176 19014 37188 19066
rect 37240 19014 37252 19066
rect 37304 19014 37316 19066
rect 37368 19014 51504 19066
rect 51556 19014 51568 19066
rect 51620 19014 51632 19066
rect 51684 19014 51696 19066
rect 51748 19014 51760 19066
rect 51812 19014 58880 19066
rect 1104 18992 58880 19014
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 4614 18952 4620 18964
rect 4571 18924 4620 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 6454 18912 6460 18964
rect 6512 18912 6518 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 8018 18952 8024 18964
rect 7156 18924 8024 18952
rect 7156 18912 7162 18924
rect 8018 18912 8024 18924
rect 8076 18952 8082 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 8076 18924 8493 18952
rect 8076 18912 8082 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 11149 18955 11207 18961
rect 11149 18921 11161 18955
rect 11195 18952 11207 18955
rect 11238 18952 11244 18964
rect 11195 18924 11244 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11698 18952 11704 18964
rect 11624 18924 11704 18952
rect 4706 18884 4712 18896
rect 3988 18856 4712 18884
rect 3988 18825 4016 18856
rect 4706 18844 4712 18856
rect 4764 18884 4770 18896
rect 4801 18887 4859 18893
rect 4801 18884 4813 18887
rect 4764 18856 4813 18884
rect 4764 18844 4770 18856
rect 4801 18853 4813 18856
rect 4847 18853 4859 18887
rect 4801 18847 4859 18853
rect 9677 18887 9735 18893
rect 9677 18853 9689 18887
rect 9723 18884 9735 18887
rect 10318 18884 10324 18896
rect 9723 18856 10324 18884
rect 9723 18853 9735 18856
rect 9677 18847 9735 18853
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18785 4031 18819
rect 4430 18816 4436 18828
rect 3973 18779 4031 18785
rect 4172 18788 4436 18816
rect 4172 18757 4200 18788
rect 4430 18776 4436 18788
rect 4488 18816 4494 18828
rect 4488 18788 5948 18816
rect 4488 18776 4494 18788
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 5675 18720 5856 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 4065 18683 4123 18689
rect 4065 18649 4077 18683
rect 4111 18680 4123 18683
rect 4985 18683 5043 18689
rect 4985 18680 4997 18683
rect 4111 18652 4997 18680
rect 4111 18649 4123 18652
rect 4065 18643 4123 18649
rect 4985 18649 4997 18652
rect 5031 18649 5043 18683
rect 4985 18643 5043 18649
rect 5828 18624 5856 18720
rect 5920 18680 5948 18788
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 7009 18819 7067 18825
rect 7009 18816 7021 18819
rect 6512 18788 7021 18816
rect 6512 18776 6518 18788
rect 7009 18785 7021 18788
rect 7055 18785 7067 18819
rect 7009 18779 7067 18785
rect 9125 18819 9183 18825
rect 9125 18785 9137 18819
rect 9171 18816 9183 18819
rect 10042 18816 10048 18828
rect 9171 18788 10048 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11624 18825 11652 18924
rect 11698 18912 11704 18924
rect 11756 18952 11762 18964
rect 13538 18952 13544 18964
rect 11756 18924 13544 18952
rect 11756 18912 11762 18924
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 27433 18955 27491 18961
rect 18340 18924 21036 18952
rect 13906 18884 13912 18896
rect 11716 18856 13912 18884
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 7837 18751 7895 18757
rect 7837 18748 7849 18751
rect 6420 18720 7849 18748
rect 6420 18708 6426 18720
rect 7837 18717 7849 18720
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8628 18720 9321 18748
rect 8628 18708 8634 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 6825 18683 6883 18689
rect 6825 18680 6837 18683
rect 5920 18652 6837 18680
rect 6825 18649 6837 18652
rect 6871 18680 6883 18683
rect 10060 18680 10088 18776
rect 11054 18708 11060 18760
rect 11112 18708 11118 18760
rect 11514 18708 11520 18760
rect 11572 18708 11578 18760
rect 11716 18680 11744 18856
rect 13906 18844 13912 18856
rect 13964 18884 13970 18896
rect 17589 18887 17647 18893
rect 13964 18856 14228 18884
rect 13964 18844 13970 18856
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12894 18816 12900 18828
rect 11839 18788 12900 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 14200 18825 14228 18856
rect 17589 18853 17601 18887
rect 17635 18884 17647 18887
rect 17954 18884 17960 18896
rect 17635 18856 17960 18884
rect 17635 18853 17647 18856
rect 17589 18847 17647 18853
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 13004 18788 13737 18816
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 6871 18652 9168 18680
rect 10060 18652 11744 18680
rect 6871 18649 6883 18652
rect 6825 18643 6883 18649
rect 9140 18624 9168 18652
rect 5810 18572 5816 18624
rect 5868 18572 5874 18624
rect 6365 18615 6423 18621
rect 6365 18581 6377 18615
rect 6411 18612 6423 18615
rect 6454 18612 6460 18624
rect 6411 18584 6460 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 6963 18584 7297 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 9122 18572 9128 18624
rect 9180 18572 9186 18624
rect 9214 18572 9220 18624
rect 9272 18572 9278 18624
rect 10410 18572 10416 18624
rect 10468 18572 10474 18624
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13004 18621 13032 18788
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 14185 18819 14243 18825
rect 14185 18785 14197 18819
rect 14231 18785 14243 18819
rect 14185 18779 14243 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 18230 18816 18236 18828
rect 17543 18788 18236 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 18230 18776 18236 18788
rect 18288 18816 18294 18828
rect 18340 18816 18368 18924
rect 18288 18788 18368 18816
rect 18288 18776 18294 18788
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 19978 18816 19984 18828
rect 19760 18788 19984 18816
rect 19760 18776 19766 18788
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 14918 18708 14924 18760
rect 14976 18708 14982 18760
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18690 18748 18696 18760
rect 18003 18720 18696 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19058 18708 19064 18760
rect 19116 18708 19122 18760
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18717 19855 18751
rect 19996 18748 20024 18776
rect 20806 18748 20812 18760
rect 19996 18720 20812 18748
rect 19797 18711 19855 18717
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 19812 18680 19840 18711
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 20254 18689 20260 18692
rect 14056 18652 14872 18680
rect 14056 18640 14062 18652
rect 12989 18615 13047 18621
rect 12989 18612 13001 18615
rect 12860 18584 13001 18612
rect 12860 18572 12866 18584
rect 12989 18581 13001 18584
rect 13035 18581 13047 18615
rect 12989 18575 13047 18581
rect 13170 18572 13176 18624
rect 13228 18572 13234 18624
rect 13538 18572 13544 18624
rect 13596 18572 13602 18624
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 14090 18612 14096 18624
rect 13679 18584 14096 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14366 18572 14372 18624
rect 14424 18572 14430 18624
rect 14844 18621 14872 18652
rect 18340 18652 19840 18680
rect 18340 18624 18368 18652
rect 14829 18615 14887 18621
rect 14829 18581 14841 18615
rect 14875 18581 14887 18615
rect 14829 18575 14887 18581
rect 15565 18615 15623 18621
rect 15565 18581 15577 18615
rect 15611 18612 15623 18615
rect 15746 18612 15752 18624
rect 15611 18584 15752 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 18046 18572 18052 18624
rect 18104 18572 18110 18624
rect 18322 18572 18328 18624
rect 18380 18572 18386 18624
rect 18414 18572 18420 18624
rect 18472 18572 18478 18624
rect 18782 18572 18788 18624
rect 18840 18612 18846 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 18840 18584 19257 18612
rect 18840 18572 18846 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 19812 18612 19840 18652
rect 20248 18643 20260 18689
rect 20254 18640 20260 18643
rect 20312 18640 20318 18692
rect 21008 18680 21036 18924
rect 27433 18921 27445 18955
rect 27479 18952 27491 18955
rect 27982 18952 27988 18964
rect 27479 18924 27988 18952
rect 27479 18921 27491 18924
rect 27433 18915 27491 18921
rect 27982 18912 27988 18924
rect 28040 18912 28046 18964
rect 30745 18955 30803 18961
rect 30745 18921 30757 18955
rect 30791 18952 30803 18955
rect 31110 18952 31116 18964
rect 30791 18924 31116 18952
rect 30791 18921 30803 18924
rect 30745 18915 30803 18921
rect 31110 18912 31116 18924
rect 31168 18912 31174 18964
rect 36906 18952 36912 18964
rect 32232 18924 36912 18952
rect 21361 18887 21419 18893
rect 21361 18853 21373 18887
rect 21407 18884 21419 18887
rect 22094 18884 22100 18896
rect 21407 18856 22100 18884
rect 21407 18853 21419 18856
rect 21361 18847 21419 18853
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 22189 18887 22247 18893
rect 22189 18853 22201 18887
rect 22235 18884 22247 18887
rect 24397 18887 24455 18893
rect 22235 18856 22876 18884
rect 22235 18853 22247 18856
rect 22189 18847 22247 18853
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 22848 18825 22876 18856
rect 24397 18853 24409 18887
rect 24443 18853 24455 18887
rect 24397 18847 24455 18853
rect 21545 18819 21603 18825
rect 21545 18816 21557 18819
rect 21232 18788 21557 18816
rect 21232 18776 21238 18788
rect 21545 18785 21557 18788
rect 21591 18785 21603 18819
rect 21545 18779 21603 18785
rect 22833 18819 22891 18825
rect 22833 18785 22845 18819
rect 22879 18785 22891 18819
rect 22833 18779 22891 18785
rect 24213 18819 24271 18825
rect 24213 18785 24225 18819
rect 24259 18816 24271 18819
rect 24412 18816 24440 18847
rect 30926 18844 30932 18896
rect 30984 18884 30990 18896
rect 31570 18884 31576 18896
rect 30984 18856 31576 18884
rect 30984 18844 30990 18856
rect 31570 18844 31576 18856
rect 31628 18884 31634 18896
rect 32232 18884 32260 18924
rect 36906 18912 36912 18924
rect 36964 18912 36970 18964
rect 39666 18912 39672 18964
rect 39724 18952 39730 18964
rect 40957 18955 41015 18961
rect 40957 18952 40969 18955
rect 39724 18924 40969 18952
rect 39724 18912 39730 18924
rect 40957 18921 40969 18924
rect 41003 18952 41015 18955
rect 41414 18952 41420 18964
rect 41003 18924 41420 18952
rect 41003 18921 41015 18924
rect 40957 18915 41015 18921
rect 35437 18887 35495 18893
rect 31628 18856 32260 18884
rect 31628 18844 31634 18856
rect 24259 18788 24440 18816
rect 25041 18819 25099 18825
rect 24259 18785 24271 18788
rect 24213 18779 24271 18785
rect 25041 18785 25053 18819
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 26513 18819 26571 18825
rect 26513 18785 26525 18819
rect 26559 18816 26571 18819
rect 27157 18819 27215 18825
rect 27157 18816 27169 18819
rect 26559 18788 27169 18816
rect 26559 18785 26571 18788
rect 26513 18779 26571 18785
rect 27157 18785 27169 18788
rect 27203 18785 27215 18819
rect 27157 18779 27215 18785
rect 21910 18708 21916 18760
rect 21968 18748 21974 18760
rect 22278 18748 22284 18760
rect 21968 18720 22284 18748
rect 21968 18708 21974 18720
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18748 23535 18751
rect 25056 18748 25084 18779
rect 25222 18748 25228 18760
rect 23523 18720 25228 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 23492 18680 23520 18711
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 21008 18652 23520 18680
rect 25884 18624 25912 18711
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 26292 18720 26985 18748
rect 26292 18708 26298 18720
rect 26973 18717 26985 18720
rect 27019 18717 27031 18751
rect 27172 18748 27200 18779
rect 27246 18776 27252 18828
rect 27304 18816 27310 18828
rect 32232 18825 32260 18856
rect 34808 18856 35204 18884
rect 27985 18819 28043 18825
rect 27985 18816 27997 18819
rect 27304 18788 27997 18816
rect 27304 18776 27310 18788
rect 27985 18785 27997 18788
rect 28031 18785 28043 18819
rect 31297 18819 31355 18825
rect 31297 18816 31309 18819
rect 27985 18779 28043 18785
rect 31036 18788 31309 18816
rect 27801 18751 27859 18757
rect 27172 18720 27292 18748
rect 26973 18711 27031 18717
rect 27264 18624 27292 18720
rect 27801 18717 27813 18751
rect 27847 18748 27859 18751
rect 28258 18748 28264 18760
rect 27847 18720 28264 18748
rect 27847 18717 27859 18720
rect 27801 18711 27859 18717
rect 28258 18708 28264 18720
rect 28316 18708 28322 18760
rect 28810 18708 28816 18760
rect 28868 18708 28874 18760
rect 28902 18708 28908 18760
rect 28960 18748 28966 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 28960 18720 30113 18748
rect 28960 18708 28966 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 27890 18640 27896 18692
rect 27948 18680 27954 18692
rect 28718 18680 28724 18692
rect 27948 18652 28724 18680
rect 27948 18640 27954 18652
rect 28718 18640 28724 18652
rect 28776 18640 28782 18692
rect 20346 18612 20352 18624
rect 19812 18584 20352 18612
rect 19245 18575 19303 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 20898 18572 20904 18624
rect 20956 18612 20962 18624
rect 21726 18612 21732 18624
rect 20956 18584 21732 18612
rect 20956 18572 20962 18584
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 21818 18572 21824 18624
rect 21876 18572 21882 18624
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22244 18584 22293 18612
rect 22244 18572 22250 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 23566 18572 23572 18624
rect 23624 18572 23630 18624
rect 24762 18572 24768 18624
rect 24820 18572 24826 18624
rect 24857 18615 24915 18621
rect 24857 18581 24869 18615
rect 24903 18612 24915 18615
rect 25225 18615 25283 18621
rect 25225 18612 25237 18615
rect 24903 18584 25237 18612
rect 24903 18581 24915 18584
rect 24857 18575 24915 18581
rect 25225 18581 25237 18584
rect 25271 18581 25283 18615
rect 25225 18575 25283 18581
rect 25866 18572 25872 18624
rect 25924 18572 25930 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 26605 18615 26663 18621
rect 26605 18612 26617 18615
rect 26292 18584 26617 18612
rect 26292 18572 26298 18584
rect 26605 18581 26617 18584
rect 26651 18581 26663 18615
rect 26605 18575 26663 18581
rect 27062 18572 27068 18624
rect 27120 18572 27126 18624
rect 27246 18572 27252 18624
rect 27304 18572 27310 18624
rect 28258 18572 28264 18624
rect 28316 18572 28322 18624
rect 29546 18572 29552 18624
rect 29604 18572 29610 18624
rect 30653 18615 30711 18621
rect 30653 18581 30665 18615
rect 30699 18612 30711 18615
rect 31036 18612 31064 18788
rect 31297 18785 31309 18788
rect 31343 18785 31355 18819
rect 31297 18779 31355 18785
rect 32217 18819 32275 18825
rect 32217 18785 32229 18819
rect 32263 18785 32275 18819
rect 32217 18779 32275 18785
rect 33045 18819 33103 18825
rect 33045 18785 33057 18819
rect 33091 18816 33103 18819
rect 33134 18816 33140 18828
rect 33091 18788 33140 18816
rect 33091 18785 33103 18788
rect 33045 18779 33103 18785
rect 33134 18776 33140 18788
rect 33192 18816 33198 18828
rect 34808 18816 34836 18856
rect 35176 18828 35204 18856
rect 35437 18853 35449 18887
rect 35483 18853 35495 18887
rect 35437 18847 35495 18853
rect 33192 18788 34836 18816
rect 33192 18776 33198 18788
rect 34882 18776 34888 18828
rect 34940 18776 34946 18828
rect 35158 18776 35164 18828
rect 35216 18776 35222 18828
rect 35452 18816 35480 18847
rect 36081 18819 36139 18825
rect 36081 18816 36093 18819
rect 35452 18788 36093 18816
rect 36081 18785 36093 18788
rect 36127 18785 36139 18819
rect 36924 18816 36952 18912
rect 37737 18887 37795 18893
rect 37737 18853 37749 18887
rect 37783 18884 37795 18887
rect 37783 18856 38424 18884
rect 37783 18853 37795 18856
rect 37737 18847 37795 18853
rect 37093 18819 37151 18825
rect 37093 18816 37105 18819
rect 36924 18788 37105 18816
rect 36081 18779 36139 18785
rect 37093 18785 37105 18788
rect 37139 18785 37151 18819
rect 37093 18779 37151 18785
rect 37277 18819 37335 18825
rect 37277 18785 37289 18819
rect 37323 18816 37335 18819
rect 38010 18816 38016 18828
rect 37323 18788 38016 18816
rect 37323 18785 37335 18788
rect 37277 18779 37335 18785
rect 38010 18776 38016 18788
rect 38068 18776 38074 18828
rect 38396 18825 38424 18856
rect 41156 18825 41184 18924
rect 41414 18912 41420 18924
rect 41472 18912 41478 18964
rect 42242 18912 42248 18964
rect 42300 18952 42306 18964
rect 42613 18955 42671 18961
rect 42613 18952 42625 18955
rect 42300 18924 42625 18952
rect 42300 18912 42306 18924
rect 42613 18921 42625 18924
rect 42659 18921 42671 18955
rect 42613 18915 42671 18921
rect 43622 18912 43628 18964
rect 43680 18952 43686 18964
rect 45557 18955 45615 18961
rect 43680 18924 43944 18952
rect 43680 18912 43686 18924
rect 42521 18887 42579 18893
rect 42521 18853 42533 18887
rect 42567 18884 42579 18887
rect 43916 18884 43944 18924
rect 45557 18921 45569 18955
rect 45603 18952 45615 18955
rect 46014 18952 46020 18964
rect 45603 18924 46020 18952
rect 45603 18921 45615 18924
rect 45557 18915 45615 18921
rect 46014 18912 46020 18924
rect 46072 18912 46078 18964
rect 54294 18952 54300 18964
rect 46124 18924 54300 18952
rect 46124 18884 46152 18924
rect 54294 18912 54300 18924
rect 54352 18912 54358 18964
rect 42567 18856 43852 18884
rect 43916 18856 46152 18884
rect 46860 18856 47532 18884
rect 42567 18853 42579 18856
rect 42521 18847 42579 18853
rect 43824 18828 43852 18856
rect 38381 18819 38439 18825
rect 38381 18785 38393 18819
rect 38427 18785 38439 18819
rect 38381 18779 38439 18785
rect 41141 18819 41199 18825
rect 41141 18785 41153 18819
rect 41187 18785 41199 18819
rect 41141 18779 41199 18785
rect 43070 18776 43076 18828
rect 43128 18816 43134 18828
rect 43165 18819 43223 18825
rect 43165 18816 43177 18819
rect 43128 18788 43177 18816
rect 43128 18776 43134 18788
rect 43165 18785 43177 18788
rect 43211 18785 43223 18819
rect 43165 18779 43223 18785
rect 43806 18776 43812 18828
rect 43864 18816 43870 18828
rect 44729 18819 44787 18825
rect 44729 18816 44741 18819
rect 43864 18788 44741 18816
rect 43864 18776 43870 18788
rect 44729 18785 44741 18788
rect 44775 18785 44787 18819
rect 44729 18779 44787 18785
rect 45465 18819 45523 18825
rect 45465 18785 45477 18819
rect 45511 18816 45523 18819
rect 46201 18819 46259 18825
rect 46201 18816 46213 18819
rect 45511 18788 46213 18816
rect 45511 18785 45523 18788
rect 45465 18779 45523 18785
rect 46201 18785 46213 18788
rect 46247 18816 46259 18819
rect 46750 18816 46756 18828
rect 46247 18788 46756 18816
rect 46247 18785 46259 18788
rect 46201 18779 46259 18785
rect 46750 18776 46756 18788
rect 46808 18776 46814 18828
rect 31113 18751 31171 18757
rect 31113 18717 31125 18751
rect 31159 18748 31171 18751
rect 31938 18748 31944 18760
rect 31159 18720 31944 18748
rect 31159 18717 31171 18720
rect 31113 18711 31171 18717
rect 31938 18708 31944 18720
rect 31996 18708 32002 18760
rect 32030 18708 32036 18760
rect 32088 18708 32094 18760
rect 33229 18751 33287 18757
rect 33229 18748 33241 18751
rect 33060 18720 33241 18748
rect 31205 18683 31263 18689
rect 31205 18649 31217 18683
rect 31251 18680 31263 18683
rect 31478 18680 31484 18692
rect 31251 18652 31484 18680
rect 31251 18649 31263 18652
rect 31205 18643 31263 18649
rect 31478 18640 31484 18652
rect 31536 18680 31542 18692
rect 33060 18680 33088 18720
rect 33229 18717 33241 18720
rect 33275 18748 33287 18751
rect 33594 18748 33600 18760
rect 33275 18720 33600 18748
rect 33275 18717 33287 18720
rect 33229 18711 33287 18717
rect 33594 18708 33600 18720
rect 33652 18748 33658 18760
rect 33652 18720 33824 18748
rect 33652 18708 33658 18720
rect 31536 18652 33088 18680
rect 33137 18683 33195 18689
rect 31536 18640 31542 18652
rect 31110 18612 31116 18624
rect 30699 18584 31116 18612
rect 30699 18581 30711 18584
rect 30653 18575 30711 18581
rect 31110 18572 31116 18584
rect 31168 18572 31174 18624
rect 31570 18572 31576 18624
rect 31628 18572 31634 18624
rect 31956 18621 31984 18652
rect 33137 18649 33149 18683
rect 33183 18680 33195 18683
rect 33689 18683 33747 18689
rect 33689 18680 33701 18683
rect 33183 18652 33701 18680
rect 33183 18649 33195 18652
rect 33137 18643 33195 18649
rect 33689 18649 33701 18652
rect 33735 18649 33747 18683
rect 33796 18680 33824 18720
rect 34238 18708 34244 18760
rect 34296 18708 34302 18760
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18748 35035 18751
rect 35894 18748 35900 18760
rect 35023 18720 35900 18748
rect 35023 18717 35035 18720
rect 34977 18711 35035 18717
rect 34992 18680 35020 18711
rect 35894 18708 35900 18720
rect 35952 18708 35958 18760
rect 36814 18708 36820 18760
rect 36872 18708 36878 18760
rect 37734 18708 37740 18760
rect 37792 18748 37798 18760
rect 38565 18751 38623 18757
rect 38565 18748 38577 18751
rect 37792 18720 38577 18748
rect 37792 18708 37798 18720
rect 38565 18717 38577 18720
rect 38611 18717 38623 18751
rect 43441 18751 43499 18757
rect 43441 18748 43453 18751
rect 38565 18711 38623 18717
rect 41156 18720 43453 18748
rect 41156 18692 41184 18720
rect 43441 18717 43453 18720
rect 43487 18717 43499 18751
rect 43441 18711 43499 18717
rect 43990 18708 43996 18760
rect 44048 18708 44054 18760
rect 45925 18751 45983 18757
rect 45925 18717 45937 18751
rect 45971 18748 45983 18751
rect 46860 18748 46888 18856
rect 47504 18828 47532 18856
rect 47578 18844 47584 18896
rect 47636 18884 47642 18896
rect 48222 18884 48228 18896
rect 47636 18856 48228 18884
rect 47636 18844 47642 18856
rect 48222 18844 48228 18856
rect 48280 18884 48286 18896
rect 52273 18887 52331 18893
rect 48280 18856 48360 18884
rect 48280 18844 48286 18856
rect 47486 18776 47492 18828
rect 47544 18816 47550 18828
rect 48332 18816 48360 18856
rect 52273 18853 52285 18887
rect 52319 18853 52331 18887
rect 52273 18847 52331 18853
rect 56137 18887 56195 18893
rect 56137 18853 56149 18887
rect 56183 18884 56195 18887
rect 58158 18884 58164 18896
rect 56183 18856 58164 18884
rect 56183 18853 56195 18856
rect 56137 18847 56195 18853
rect 48409 18819 48467 18825
rect 48409 18816 48421 18819
rect 47544 18788 48268 18816
rect 48332 18788 48421 18816
rect 47544 18776 47550 18788
rect 45971 18720 46888 18748
rect 45971 18717 45983 18720
rect 45925 18711 45983 18717
rect 47026 18708 47032 18760
rect 47084 18708 47090 18760
rect 48240 18757 48268 18788
rect 48409 18785 48421 18788
rect 48455 18785 48467 18819
rect 48409 18779 48467 18785
rect 48590 18776 48596 18828
rect 48648 18816 48654 18828
rect 48777 18819 48835 18825
rect 48777 18816 48789 18819
rect 48648 18788 48789 18816
rect 48648 18776 48654 18788
rect 48777 18785 48789 18788
rect 48823 18785 48835 18819
rect 48777 18779 48835 18785
rect 52181 18819 52239 18825
rect 52181 18785 52193 18819
rect 52227 18816 52239 18819
rect 52288 18816 52316 18847
rect 58158 18844 58164 18856
rect 58216 18844 58222 18896
rect 52227 18788 52316 18816
rect 52825 18819 52883 18825
rect 52227 18785 52239 18788
rect 52181 18779 52239 18785
rect 52825 18785 52837 18819
rect 52871 18785 52883 18819
rect 52825 18779 52883 18785
rect 55125 18819 55183 18825
rect 55125 18785 55137 18819
rect 55171 18816 55183 18819
rect 55493 18819 55551 18825
rect 55493 18816 55505 18819
rect 55171 18788 55505 18816
rect 55171 18785 55183 18788
rect 55125 18779 55183 18785
rect 55493 18785 55505 18788
rect 55539 18816 55551 18819
rect 56318 18816 56324 18828
rect 55539 18788 56324 18816
rect 55539 18785 55551 18788
rect 55493 18779 55551 18785
rect 47673 18751 47731 18757
rect 47673 18717 47685 18751
rect 47719 18717 47731 18751
rect 47673 18711 47731 18717
rect 48225 18751 48283 18757
rect 48225 18717 48237 18751
rect 48271 18748 48283 18751
rect 48271 18720 49004 18748
rect 48271 18717 48283 18720
rect 48225 18711 48283 18717
rect 33796 18652 35020 18680
rect 35069 18683 35127 18689
rect 33689 18643 33747 18649
rect 35069 18649 35081 18683
rect 35115 18680 35127 18683
rect 36265 18683 36323 18689
rect 36265 18680 36277 18683
rect 35115 18652 36277 18680
rect 35115 18649 35127 18652
rect 35069 18643 35127 18649
rect 36265 18649 36277 18652
rect 36311 18649 36323 18683
rect 36265 18643 36323 18649
rect 41138 18640 41144 18692
rect 41196 18640 41202 18692
rect 41408 18683 41466 18689
rect 41408 18649 41420 18683
rect 41454 18680 41466 18683
rect 41598 18680 41604 18692
rect 41454 18652 41604 18680
rect 41454 18649 41466 18652
rect 41408 18643 41466 18649
rect 41598 18640 41604 18652
rect 41656 18640 41662 18692
rect 43073 18683 43131 18689
rect 43073 18649 43085 18683
rect 43119 18680 43131 18683
rect 44177 18683 44235 18689
rect 44177 18680 44189 18683
rect 43119 18652 44189 18680
rect 43119 18649 43131 18652
rect 43073 18643 43131 18649
rect 44177 18649 44189 18652
rect 44223 18649 44235 18683
rect 47688 18680 47716 18711
rect 48130 18680 48136 18692
rect 44177 18643 44235 18649
rect 46216 18652 48136 18680
rect 46216 18624 46244 18652
rect 48130 18640 48136 18652
rect 48188 18640 48194 18692
rect 48317 18683 48375 18689
rect 48317 18649 48329 18683
rect 48363 18680 48375 18683
rect 48976 18680 49004 18720
rect 49050 18708 49056 18760
rect 49108 18708 49114 18760
rect 49326 18708 49332 18760
rect 49384 18708 49390 18760
rect 50338 18708 50344 18760
rect 50396 18708 50402 18760
rect 52840 18748 52868 18779
rect 56318 18776 56324 18788
rect 56376 18776 56382 18828
rect 52196 18720 52868 18748
rect 49344 18680 49372 18708
rect 52196 18692 52224 18720
rect 53650 18708 53656 18760
rect 53708 18708 53714 18760
rect 55766 18708 55772 18760
rect 55824 18708 55830 18760
rect 56594 18708 56600 18760
rect 56652 18748 56658 18760
rect 56781 18751 56839 18757
rect 56781 18748 56793 18751
rect 56652 18720 56793 18748
rect 56652 18708 56658 18720
rect 56781 18717 56793 18720
rect 56827 18717 56839 18751
rect 56781 18711 56839 18717
rect 57517 18751 57575 18757
rect 57517 18717 57529 18751
rect 57563 18717 57575 18751
rect 57517 18711 57575 18717
rect 48363 18652 48544 18680
rect 48976 18652 49372 18680
rect 48363 18649 48375 18652
rect 48317 18643 48375 18649
rect 31941 18615 31999 18621
rect 31941 18581 31953 18615
rect 31987 18612 31999 18615
rect 32677 18615 32735 18621
rect 31987 18584 32021 18612
rect 31987 18581 31999 18584
rect 31941 18575 31999 18581
rect 32677 18581 32689 18615
rect 32723 18612 32735 18615
rect 32950 18612 32956 18624
rect 32723 18584 32956 18612
rect 32723 18581 32735 18584
rect 32677 18575 32735 18581
rect 32950 18572 32956 18584
rect 33008 18572 33014 18624
rect 33594 18572 33600 18624
rect 33652 18572 33658 18624
rect 35526 18572 35532 18624
rect 35584 18572 35590 18624
rect 37369 18615 37427 18621
rect 37369 18581 37381 18615
rect 37415 18612 37427 18615
rect 37550 18612 37556 18624
rect 37415 18584 37556 18612
rect 37415 18581 37427 18584
rect 37369 18575 37427 18581
rect 37550 18572 37556 18584
rect 37608 18572 37614 18624
rect 37826 18572 37832 18624
rect 37884 18572 37890 18624
rect 39206 18572 39212 18624
rect 39264 18572 39270 18624
rect 39574 18572 39580 18624
rect 39632 18612 39638 18624
rect 42058 18612 42064 18624
rect 39632 18584 42064 18612
rect 39632 18572 39638 18584
rect 42058 18572 42064 18584
rect 42116 18572 42122 18624
rect 42978 18572 42984 18624
rect 43036 18572 43042 18624
rect 46014 18572 46020 18624
rect 46072 18572 46078 18624
rect 46198 18572 46204 18624
rect 46256 18572 46262 18624
rect 46382 18572 46388 18624
rect 46440 18572 46446 18624
rect 46658 18572 46664 18624
rect 46716 18612 46722 18624
rect 47121 18615 47179 18621
rect 47121 18612 47133 18615
rect 46716 18584 47133 18612
rect 46716 18572 46722 18584
rect 47121 18581 47133 18584
rect 47167 18581 47179 18615
rect 47121 18575 47179 18581
rect 47857 18615 47915 18621
rect 47857 18581 47869 18615
rect 47903 18612 47915 18615
rect 48406 18612 48412 18624
rect 47903 18584 48412 18612
rect 47903 18581 47915 18584
rect 47857 18575 47915 18581
rect 48406 18572 48412 18584
rect 48464 18572 48470 18624
rect 48516 18612 48544 18652
rect 52178 18640 52184 18692
rect 52236 18640 52242 18692
rect 52641 18683 52699 18689
rect 52641 18649 52653 18683
rect 52687 18680 52699 18683
rect 53006 18680 53012 18692
rect 52687 18652 53012 18680
rect 52687 18649 52699 18652
rect 52641 18643 52699 18649
rect 53006 18640 53012 18652
rect 53064 18680 53070 18692
rect 53064 18652 55628 18680
rect 53064 18640 53070 18652
rect 55600 18624 55628 18652
rect 48866 18612 48872 18624
rect 48516 18584 48872 18612
rect 48866 18572 48872 18584
rect 48924 18572 48930 18624
rect 48958 18572 48964 18624
rect 49016 18572 49022 18624
rect 49142 18572 49148 18624
rect 49200 18612 49206 18624
rect 49421 18615 49479 18621
rect 49421 18612 49433 18615
rect 49200 18584 49433 18612
rect 49200 18572 49206 18584
rect 49421 18581 49433 18584
rect 49467 18581 49479 18615
rect 49421 18575 49479 18581
rect 50982 18572 50988 18624
rect 51040 18572 51046 18624
rect 51537 18615 51595 18621
rect 51537 18581 51549 18615
rect 51583 18612 51595 18615
rect 51902 18612 51908 18624
rect 51583 18584 51908 18612
rect 51583 18581 51595 18584
rect 51537 18575 51595 18581
rect 51902 18572 51908 18584
rect 51960 18572 51966 18624
rect 52730 18572 52736 18624
rect 52788 18572 52794 18624
rect 52822 18572 52828 18624
rect 52880 18612 52886 18624
rect 53101 18615 53159 18621
rect 53101 18612 53113 18615
rect 52880 18584 53113 18612
rect 52880 18572 52886 18584
rect 53101 18581 53113 18584
rect 53147 18581 53159 18615
rect 53101 18575 53159 18581
rect 54113 18615 54171 18621
rect 54113 18581 54125 18615
rect 54159 18612 54171 18615
rect 54570 18612 54576 18624
rect 54159 18584 54576 18612
rect 54159 18581 54171 18584
rect 54113 18575 54171 18581
rect 54570 18572 54576 18584
rect 54628 18572 54634 18624
rect 55582 18572 55588 18624
rect 55640 18572 55646 18624
rect 55674 18572 55680 18624
rect 55732 18572 55738 18624
rect 56226 18572 56232 18624
rect 56284 18572 56290 18624
rect 56962 18572 56968 18624
rect 57020 18572 57026 18624
rect 57238 18572 57244 18624
rect 57296 18612 57302 18624
rect 57532 18612 57560 18711
rect 57296 18584 57560 18612
rect 57296 18572 57302 18584
rect 1104 18522 59040 18544
rect 1104 18470 15394 18522
rect 15446 18470 15458 18522
rect 15510 18470 15522 18522
rect 15574 18470 15586 18522
rect 15638 18470 15650 18522
rect 15702 18470 29838 18522
rect 29890 18470 29902 18522
rect 29954 18470 29966 18522
rect 30018 18470 30030 18522
rect 30082 18470 30094 18522
rect 30146 18470 44282 18522
rect 44334 18470 44346 18522
rect 44398 18470 44410 18522
rect 44462 18470 44474 18522
rect 44526 18470 44538 18522
rect 44590 18470 58726 18522
rect 58778 18470 58790 18522
rect 58842 18470 58854 18522
rect 58906 18470 58918 18522
rect 58970 18470 58982 18522
rect 59034 18470 59040 18522
rect 1104 18448 59040 18470
rect 8205 18411 8263 18417
rect 6564 18380 8064 18408
rect 4700 18343 4758 18349
rect 2976 18312 4292 18340
rect 2976 18281 3004 18312
rect 4264 18284 4292 18312
rect 4700 18309 4712 18343
rect 4746 18340 4758 18343
rect 5258 18340 5264 18352
rect 4746 18312 5264 18340
rect 4746 18309 4758 18312
rect 4700 18303 4758 18309
rect 5258 18300 5264 18312
rect 5316 18300 5322 18352
rect 2961 18275 3019 18281
rect 2961 18272 2973 18275
rect 2746 18244 2973 18272
rect 2130 18164 2136 18216
rect 2188 18204 2194 18216
rect 2746 18204 2774 18244
rect 2961 18241 2973 18244
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3228 18275 3286 18281
rect 3228 18241 3240 18275
rect 3274 18272 3286 18275
rect 3510 18272 3516 18284
rect 3274 18244 3516 18272
rect 3274 18241 3286 18244
rect 3228 18235 3286 18241
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4304 18244 4445 18272
rect 4304 18232 4310 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 6362 18232 6368 18284
rect 6420 18232 6426 18284
rect 6564 18213 6592 18380
rect 8036 18340 8064 18380
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 9214 18408 9220 18420
rect 8251 18380 9220 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 11112 18380 11529 18408
rect 11112 18368 11118 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 11885 18411 11943 18417
rect 11885 18408 11897 18411
rect 11756 18380 11897 18408
rect 11756 18368 11762 18380
rect 11885 18377 11897 18380
rect 11931 18377 11943 18411
rect 11885 18371 11943 18377
rect 11974 18368 11980 18420
rect 12032 18368 12038 18420
rect 12621 18411 12679 18417
rect 12621 18377 12633 18411
rect 12667 18408 12679 18411
rect 14366 18408 14372 18420
rect 12667 18380 14372 18408
rect 12667 18377 12679 18380
rect 12621 18371 12679 18377
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 18322 18368 18328 18420
rect 18380 18368 18386 18420
rect 18414 18368 18420 18420
rect 18472 18368 18478 18420
rect 18782 18368 18788 18420
rect 18840 18368 18846 18420
rect 19058 18368 19064 18420
rect 19116 18408 19122 18420
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 19116 18380 19165 18408
rect 19116 18368 19122 18380
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 20898 18408 20904 18420
rect 19153 18371 19211 18377
rect 19812 18380 20904 18408
rect 8036 18312 8340 18340
rect 8312 18272 8340 18312
rect 8846 18300 8852 18352
rect 8904 18300 8910 18352
rect 10220 18343 10278 18349
rect 10220 18309 10232 18343
rect 10266 18340 10278 18343
rect 10686 18340 10692 18352
rect 10266 18312 10692 18340
rect 10266 18309 10278 18312
rect 10220 18303 10278 18309
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 15746 18300 15752 18352
rect 15804 18349 15810 18352
rect 15804 18340 15816 18349
rect 17212 18343 17270 18349
rect 15804 18312 15849 18340
rect 15804 18303 15816 18312
rect 17212 18309 17224 18343
rect 17258 18340 17270 18343
rect 18432 18340 18460 18368
rect 17258 18312 18460 18340
rect 17258 18309 17270 18312
rect 17212 18303 17270 18309
rect 15804 18300 15810 18303
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 19812 18340 19840 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 22649 18411 22707 18417
rect 22649 18408 22661 18411
rect 21876 18380 22661 18408
rect 21876 18368 21882 18380
rect 22649 18377 22661 18380
rect 22695 18377 22707 18411
rect 22649 18371 22707 18377
rect 23566 18368 23572 18420
rect 23624 18368 23630 18420
rect 24949 18411 25007 18417
rect 24949 18377 24961 18411
rect 24995 18408 25007 18411
rect 27062 18408 27068 18420
rect 24995 18380 27068 18408
rect 24995 18377 25007 18380
rect 24949 18371 25007 18377
rect 27062 18368 27068 18380
rect 27120 18368 27126 18420
rect 28534 18368 28540 18420
rect 28592 18368 28598 18420
rect 28629 18411 28687 18417
rect 28629 18377 28641 18411
rect 28675 18408 28687 18411
rect 28810 18408 28816 18420
rect 28675 18380 28816 18408
rect 28675 18377 28687 18380
rect 28629 18371 28687 18377
rect 28810 18368 28816 18380
rect 28868 18368 28874 18420
rect 29089 18411 29147 18417
rect 29089 18377 29101 18411
rect 29135 18408 29147 18411
rect 29546 18408 29552 18420
rect 29135 18380 29552 18408
rect 29135 18377 29147 18380
rect 29089 18371 29147 18377
rect 29546 18368 29552 18380
rect 29604 18368 29610 18420
rect 32398 18368 32404 18420
rect 32456 18408 32462 18420
rect 33870 18408 33876 18420
rect 32456 18380 33876 18408
rect 32456 18368 32462 18380
rect 33870 18368 33876 18380
rect 33928 18368 33934 18420
rect 34425 18411 34483 18417
rect 34425 18377 34437 18411
rect 34471 18408 34483 18411
rect 36814 18408 36820 18420
rect 34471 18380 36820 18408
rect 34471 18377 34483 18380
rect 34425 18371 34483 18377
rect 23584 18340 23612 18368
rect 27430 18349 27436 18352
rect 23722 18343 23780 18349
rect 23722 18340 23734 18343
rect 18748 18312 19840 18340
rect 21284 18312 23244 18340
rect 23584 18312 23734 18340
rect 18748 18300 18754 18312
rect 8864 18272 8892 18300
rect 8312 18244 8892 18272
rect 9421 18275 9479 18281
rect 2188 18176 2774 18204
rect 6549 18207 6607 18213
rect 2188 18164 2194 18176
rect 6549 18173 6561 18207
rect 6595 18173 6607 18207
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6549 18167 6607 18173
rect 6656 18176 7297 18204
rect 5810 18096 5816 18148
rect 5868 18136 5874 18148
rect 6656 18136 6684 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 7374 18164 7380 18216
rect 7432 18213 7438 18216
rect 7432 18207 7460 18213
rect 7448 18173 7460 18207
rect 7432 18167 7460 18173
rect 7432 18164 7438 18167
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 7616 18176 8064 18204
rect 7616 18164 7622 18176
rect 5868 18108 6684 18136
rect 7009 18139 7067 18145
rect 5868 18096 5874 18108
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 7098 18136 7104 18148
rect 7055 18108 7104 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 5442 18068 5448 18080
rect 4387 18040 5448 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 5442 18028 5448 18040
rect 5500 18068 5506 18080
rect 7374 18068 7380 18080
rect 5500 18040 7380 18068
rect 5500 18028 5506 18040
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 8036 18068 8064 18176
rect 8312 18145 8340 18244
rect 9421 18241 9433 18275
rect 9467 18272 9479 18275
rect 9766 18272 9772 18284
rect 9467 18244 9772 18272
rect 9467 18241 9479 18244
rect 9421 18235 9479 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16025 18275 16083 18281
rect 16025 18272 16037 18275
rect 15988 18244 16037 18272
rect 15988 18232 15994 18244
rect 16025 18241 16037 18244
rect 16071 18272 16083 18275
rect 16942 18272 16948 18284
rect 16071 18244 16948 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 20346 18232 20352 18284
rect 20404 18281 20410 18284
rect 20404 18275 20453 18281
rect 20404 18241 20407 18275
rect 20441 18241 20453 18275
rect 20404 18235 20453 18241
rect 20404 18232 20410 18235
rect 21284 18216 21312 18312
rect 21358 18232 21364 18284
rect 21416 18272 21422 18284
rect 23216 18281 23244 18312
rect 23722 18309 23734 18312
rect 23768 18309 23780 18343
rect 27424 18340 27436 18349
rect 27391 18312 27436 18340
rect 23722 18303 23780 18309
rect 27424 18303 27436 18312
rect 27430 18300 27436 18303
rect 27488 18300 27494 18352
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 21416 18244 22201 18272
rect 21416 18232 21422 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 23201 18275 23259 18281
rect 23201 18241 23213 18275
rect 23247 18241 23259 18275
rect 23201 18235 23259 18241
rect 26605 18275 26663 18281
rect 26605 18241 26617 18275
rect 26651 18272 26663 18275
rect 28552 18272 28580 18368
rect 28718 18300 28724 18352
rect 28776 18340 28782 18352
rect 28997 18343 29055 18349
rect 28997 18340 29009 18343
rect 28776 18312 29009 18340
rect 28776 18300 28782 18312
rect 28997 18309 29009 18312
rect 29043 18309 29055 18343
rect 28997 18303 29055 18309
rect 30368 18343 30426 18349
rect 30368 18309 30380 18343
rect 30414 18340 30426 18343
rect 30558 18340 30564 18352
rect 30414 18312 30564 18340
rect 30414 18309 30426 18312
rect 30368 18303 30426 18309
rect 30558 18300 30564 18312
rect 30616 18300 30622 18352
rect 26651 18244 28580 18272
rect 26651 18241 26663 18244
rect 26605 18235 26663 18241
rect 29730 18232 29736 18284
rect 29788 18272 29794 18284
rect 30101 18275 30159 18281
rect 30101 18272 30113 18275
rect 29788 18244 30113 18272
rect 29788 18232 29794 18244
rect 30101 18241 30113 18244
rect 30147 18241 30159 18275
rect 30101 18235 30159 18241
rect 33134 18232 33140 18284
rect 33192 18232 33198 18284
rect 34149 18275 34207 18281
rect 34149 18241 34161 18275
rect 34195 18272 34207 18275
rect 34440 18272 34468 18371
rect 36814 18368 36820 18380
rect 36872 18368 36878 18420
rect 37826 18368 37832 18420
rect 37884 18368 37890 18420
rect 38654 18368 38660 18420
rect 38712 18368 38718 18420
rect 39025 18411 39083 18417
rect 39025 18377 39037 18411
rect 39071 18408 39083 18411
rect 39206 18408 39212 18420
rect 39071 18380 39212 18408
rect 39071 18377 39083 18380
rect 39025 18371 39083 18377
rect 39206 18368 39212 18380
rect 39264 18368 39270 18420
rect 43165 18411 43223 18417
rect 43165 18377 43177 18411
rect 43211 18408 43223 18411
rect 43990 18408 43996 18420
rect 43211 18380 43996 18408
rect 43211 18377 43223 18380
rect 43165 18371 43223 18377
rect 43990 18368 43996 18380
rect 44048 18368 44054 18420
rect 44729 18411 44787 18417
rect 44729 18377 44741 18411
rect 44775 18408 44787 18411
rect 45002 18408 45008 18420
rect 44775 18380 45008 18408
rect 44775 18377 44787 18380
rect 44729 18371 44787 18377
rect 35342 18300 35348 18352
rect 35400 18340 35406 18352
rect 37544 18343 37602 18349
rect 35400 18312 35848 18340
rect 35400 18300 35406 18312
rect 34195 18244 34468 18272
rect 34195 18241 34207 18244
rect 34149 18235 34207 18241
rect 35526 18232 35532 18284
rect 35584 18281 35590 18284
rect 35820 18281 35848 18312
rect 37544 18309 37556 18343
rect 37590 18340 37602 18343
rect 37844 18340 37872 18368
rect 41414 18340 41420 18352
rect 37590 18312 37872 18340
rect 40880 18312 41420 18340
rect 37590 18309 37602 18312
rect 37544 18303 37602 18309
rect 40880 18281 40908 18312
rect 41414 18300 41420 18312
rect 41472 18340 41478 18352
rect 42610 18340 42616 18352
rect 41472 18312 42616 18340
rect 41472 18300 41478 18312
rect 42610 18300 42616 18312
rect 42668 18300 42674 18352
rect 42978 18340 42984 18352
rect 42720 18312 42984 18340
rect 41138 18281 41144 18284
rect 35584 18272 35596 18281
rect 35805 18275 35863 18281
rect 35584 18244 35629 18272
rect 35584 18235 35596 18244
rect 35805 18241 35817 18275
rect 35851 18272 35863 18275
rect 37001 18275 37059 18281
rect 37001 18272 37013 18275
rect 35851 18244 37013 18272
rect 35851 18241 35863 18244
rect 35805 18235 35863 18241
rect 37001 18241 37013 18244
rect 37047 18272 37059 18275
rect 37277 18275 37335 18281
rect 37277 18272 37289 18275
rect 37047 18244 37289 18272
rect 37047 18241 37059 18244
rect 37001 18235 37059 18241
rect 37277 18241 37289 18244
rect 37323 18241 37335 18275
rect 39117 18275 39175 18281
rect 39117 18272 39129 18275
rect 37277 18235 37335 18241
rect 38304 18244 39129 18272
rect 35584 18232 35590 18235
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 9953 18207 10011 18213
rect 9953 18204 9965 18207
rect 9723 18176 9965 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 9953 18173 9965 18176
rect 9999 18173 10011 18207
rect 9953 18167 10011 18173
rect 12161 18207 12219 18213
rect 12161 18173 12173 18207
rect 12207 18204 12219 18207
rect 12710 18204 12716 18216
rect 12207 18176 12716 18204
rect 12207 18173 12219 18176
rect 12161 18167 12219 18173
rect 8297 18139 8355 18145
rect 8297 18105 8309 18139
rect 8343 18105 8355 18139
rect 8297 18099 8355 18105
rect 8662 18068 8668 18080
rect 8036 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9968 18068 9996 18167
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 13403 18207 13461 18213
rect 13403 18204 13415 18207
rect 12912 18176 13415 18204
rect 12912 18136 12940 18176
rect 13403 18173 13415 18176
rect 13449 18173 13461 18207
rect 13403 18167 13461 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 14277 18207 14335 18213
rect 13587 18176 13768 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 12406 18108 12940 18136
rect 10226 18068 10232 18080
rect 9968 18040 10232 18068
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 12406 18068 12434 18108
rect 11388 18040 12434 18068
rect 11388 18028 11394 18040
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 13740 18068 13768 18176
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 13814 18096 13820 18148
rect 13872 18096 13878 18148
rect 12584 18040 13768 18068
rect 14292 18068 14320 18167
rect 14458 18164 14464 18216
rect 14516 18164 14522 18216
rect 18322 18164 18328 18216
rect 18380 18204 18386 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18380 18176 18521 18204
rect 18380 18164 18386 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19886 18204 19892 18216
rect 19567 18176 19892 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 19886 18164 19892 18176
rect 19944 18204 19950 18216
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 19944 18176 20269 18204
rect 19944 18164 19950 18176
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 20530 18164 20536 18216
rect 20588 18164 20594 18216
rect 21266 18164 21272 18216
rect 21324 18164 21330 18216
rect 21453 18207 21511 18213
rect 21453 18173 21465 18207
rect 21499 18204 21511 18207
rect 22094 18204 22100 18216
rect 21499 18176 22100 18204
rect 21499 18173 21511 18176
rect 21453 18167 21511 18173
rect 22094 18164 22100 18176
rect 22152 18164 22158 18216
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18105 19671 18139
rect 19613 18099 19671 18105
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14292 18040 14657 18068
rect 12584 18028 12590 18040
rect 14645 18037 14657 18040
rect 14691 18068 14703 18071
rect 16206 18068 16212 18080
rect 14691 18040 16212 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 19628 18068 19656 18099
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 20809 18139 20867 18145
rect 20809 18136 20821 18139
rect 20772 18108 20821 18136
rect 20772 18096 20778 18108
rect 20809 18105 20821 18108
rect 20855 18105 20867 18139
rect 22296 18136 22324 18167
rect 22370 18164 22376 18216
rect 22428 18164 22434 18216
rect 23474 18164 23480 18216
rect 23532 18164 23538 18216
rect 25590 18164 25596 18216
rect 25648 18164 25654 18216
rect 25774 18213 25780 18216
rect 25752 18207 25780 18213
rect 25752 18173 25764 18207
rect 25752 18167 25780 18173
rect 25774 18164 25780 18167
rect 25832 18164 25838 18216
rect 25866 18164 25872 18216
rect 25924 18204 25930 18216
rect 25924 18176 26096 18204
rect 25924 18164 25930 18176
rect 20809 18099 20867 18105
rect 20916 18108 22324 18136
rect 24857 18139 24915 18145
rect 20916 18068 20944 18108
rect 24857 18105 24869 18139
rect 24903 18136 24915 18139
rect 24903 18108 25268 18136
rect 24903 18105 24915 18108
rect 24857 18099 24915 18105
rect 19628 18040 20944 18068
rect 21818 18028 21824 18080
rect 21876 18028 21882 18080
rect 25240 18068 25268 18108
rect 26068 18068 26096 18176
rect 26142 18164 26148 18216
rect 26200 18164 26206 18216
rect 26789 18207 26847 18213
rect 26789 18173 26801 18207
rect 26835 18204 26847 18207
rect 26835 18176 27016 18204
rect 26835 18173 26847 18176
rect 26789 18167 26847 18173
rect 25240 18040 26096 18068
rect 26988 18068 27016 18176
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 27120 18176 27169 18204
rect 27120 18164 27126 18176
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 29178 18164 29184 18216
rect 29236 18164 29242 18216
rect 32766 18204 32772 18216
rect 31726 18176 32772 18204
rect 31481 18139 31539 18145
rect 31481 18105 31493 18139
rect 31527 18136 31539 18139
rect 31726 18136 31754 18176
rect 32766 18164 32772 18176
rect 32824 18204 32830 18216
rect 33275 18207 33333 18213
rect 33275 18204 33287 18207
rect 32824 18176 33287 18204
rect 32824 18164 32830 18176
rect 33275 18173 33287 18176
rect 33321 18173 33333 18207
rect 33275 18167 33333 18173
rect 33410 18164 33416 18216
rect 33468 18164 33474 18216
rect 34238 18164 34244 18216
rect 34296 18204 34302 18216
rect 34333 18207 34391 18213
rect 34333 18204 34345 18207
rect 34296 18176 34345 18204
rect 34296 18164 34302 18176
rect 34333 18173 34345 18176
rect 34379 18173 34391 18207
rect 34333 18167 34391 18173
rect 31527 18108 31754 18136
rect 33689 18139 33747 18145
rect 31527 18105 31539 18108
rect 31481 18099 31539 18105
rect 33689 18105 33701 18139
rect 33735 18136 33747 18139
rect 33870 18136 33876 18148
rect 33735 18108 33876 18136
rect 33735 18105 33747 18108
rect 33689 18099 33747 18105
rect 33870 18096 33876 18108
rect 33928 18136 33934 18148
rect 33928 18108 34468 18136
rect 33928 18096 33934 18108
rect 28902 18068 28908 18080
rect 26988 18040 28908 18068
rect 28902 18028 28908 18040
rect 28960 18028 28966 18080
rect 31849 18071 31907 18077
rect 31849 18037 31861 18071
rect 31895 18068 31907 18071
rect 31938 18068 31944 18080
rect 31895 18040 31944 18068
rect 31895 18037 31907 18040
rect 31849 18031 31907 18037
rect 31938 18028 31944 18040
rect 31996 18068 32002 18080
rect 32122 18068 32128 18080
rect 31996 18040 32128 18068
rect 31996 18028 32002 18040
rect 32122 18028 32128 18040
rect 32180 18028 32186 18080
rect 32493 18071 32551 18077
rect 32493 18037 32505 18071
rect 32539 18068 32551 18071
rect 33778 18068 33784 18080
rect 32539 18040 33784 18068
rect 32539 18037 32551 18040
rect 32493 18031 32551 18037
rect 33778 18028 33784 18040
rect 33836 18028 33842 18080
rect 34440 18068 34468 18108
rect 35986 18068 35992 18080
rect 34440 18040 35992 18068
rect 35986 18028 35992 18040
rect 36044 18028 36050 18080
rect 37550 18028 37556 18080
rect 37608 18068 37614 18080
rect 38304 18068 38332 18244
rect 39117 18241 39129 18244
rect 39163 18241 39175 18275
rect 39117 18235 39175 18241
rect 40865 18275 40923 18281
rect 40865 18241 40877 18275
rect 40911 18241 40923 18275
rect 41132 18272 41144 18281
rect 41099 18244 41144 18272
rect 40865 18235 40923 18241
rect 41132 18235 41144 18244
rect 41138 18232 41144 18235
rect 41196 18232 41202 18284
rect 42242 18232 42248 18284
rect 42300 18272 42306 18284
rect 42720 18281 42748 18312
rect 42978 18300 42984 18312
rect 43036 18300 43042 18352
rect 44836 18281 44864 18380
rect 45002 18368 45008 18380
rect 45060 18368 45066 18420
rect 46198 18368 46204 18420
rect 46256 18368 46262 18420
rect 46382 18368 46388 18420
rect 46440 18368 46446 18420
rect 46658 18368 46664 18420
rect 46716 18368 46722 18420
rect 47026 18368 47032 18420
rect 47084 18368 47090 18420
rect 47486 18368 47492 18420
rect 47544 18368 47550 18420
rect 47581 18411 47639 18417
rect 47581 18377 47593 18411
rect 47627 18408 47639 18411
rect 48958 18408 48964 18420
rect 47627 18380 48964 18408
rect 47627 18377 47639 18380
rect 47581 18371 47639 18377
rect 48958 18368 48964 18380
rect 49016 18368 49022 18420
rect 50982 18368 50988 18420
rect 51040 18368 51046 18420
rect 52546 18368 52552 18420
rect 52604 18368 52610 18420
rect 52822 18368 52828 18420
rect 52880 18368 52886 18420
rect 52914 18368 52920 18420
rect 52972 18408 52978 18420
rect 53101 18411 53159 18417
rect 53101 18408 53113 18411
rect 52972 18380 53113 18408
rect 52972 18368 52978 18380
rect 53101 18377 53113 18380
rect 53147 18377 53159 18411
rect 53101 18371 53159 18377
rect 53469 18411 53527 18417
rect 53469 18377 53481 18411
rect 53515 18408 53527 18411
rect 53650 18408 53656 18420
rect 53515 18380 53656 18408
rect 53515 18377 53527 18380
rect 53469 18371 53527 18377
rect 53650 18368 53656 18380
rect 53708 18368 53714 18420
rect 53929 18411 53987 18417
rect 53929 18377 53941 18411
rect 53975 18408 53987 18411
rect 55674 18408 55680 18420
rect 53975 18380 55680 18408
rect 53975 18377 53987 18380
rect 53929 18371 53987 18377
rect 55674 18368 55680 18380
rect 55732 18368 55738 18420
rect 56686 18408 56692 18420
rect 56060 18380 56692 18408
rect 42705 18275 42763 18281
rect 42705 18272 42717 18275
rect 42300 18244 42717 18272
rect 42300 18232 42306 18244
rect 42705 18241 42717 18244
rect 42751 18241 42763 18275
rect 42705 18235 42763 18241
rect 42797 18275 42855 18281
rect 42797 18241 42809 18275
rect 42843 18272 42855 18275
rect 43257 18275 43315 18281
rect 43257 18272 43269 18275
rect 42843 18244 43269 18272
rect 42843 18241 42855 18244
rect 42797 18235 42855 18241
rect 43257 18241 43269 18244
rect 43303 18241 43315 18275
rect 43257 18235 43315 18241
rect 44821 18275 44879 18281
rect 44821 18241 44833 18275
rect 44867 18241 44879 18275
rect 44821 18235 44879 18241
rect 45088 18275 45146 18281
rect 45088 18241 45100 18275
rect 45134 18272 45146 18275
rect 46400 18272 46428 18368
rect 46569 18343 46627 18349
rect 46569 18309 46581 18343
rect 46615 18340 46627 18343
rect 47504 18340 47532 18368
rect 46615 18312 47532 18340
rect 46615 18309 46627 18312
rect 46569 18303 46627 18309
rect 47670 18300 47676 18352
rect 47728 18300 47734 18352
rect 50648 18343 50706 18349
rect 50648 18309 50660 18343
rect 50694 18340 50706 18343
rect 51000 18340 51028 18368
rect 50694 18312 51028 18340
rect 51436 18343 51494 18349
rect 50694 18309 50706 18312
rect 50648 18303 50706 18309
rect 51436 18309 51448 18343
rect 51482 18340 51494 18343
rect 52840 18340 52868 18368
rect 51482 18312 52868 18340
rect 51482 18309 51494 18312
rect 51436 18303 51494 18309
rect 53006 18300 53012 18352
rect 53064 18300 53070 18352
rect 56060 18340 56088 18380
rect 56686 18368 56692 18380
rect 56744 18368 56750 18420
rect 57238 18408 57244 18420
rect 56888 18380 57244 18408
rect 55600 18312 56088 18340
rect 56128 18343 56186 18349
rect 45134 18244 46428 18272
rect 45134 18241 45146 18244
rect 45088 18235 45146 18241
rect 38746 18164 38752 18216
rect 38804 18204 38810 18216
rect 38933 18207 38991 18213
rect 38933 18204 38945 18207
rect 38804 18176 38945 18204
rect 38804 18164 38810 18176
rect 38933 18173 38945 18176
rect 38979 18204 38991 18207
rect 39574 18204 39580 18216
rect 38979 18176 39580 18204
rect 38979 18173 38991 18176
rect 38933 18167 38991 18173
rect 39574 18164 39580 18176
rect 39632 18164 39638 18216
rect 40129 18207 40187 18213
rect 40129 18173 40141 18207
rect 40175 18173 40187 18207
rect 40129 18167 40187 18173
rect 39485 18139 39543 18145
rect 39485 18105 39497 18139
rect 39531 18136 39543 18139
rect 40144 18136 40172 18167
rect 42518 18164 42524 18216
rect 42576 18164 42582 18216
rect 43809 18207 43867 18213
rect 43809 18173 43821 18207
rect 43855 18173 43867 18207
rect 43809 18167 43867 18173
rect 46477 18207 46535 18213
rect 46477 18173 46489 18207
rect 46523 18204 46535 18207
rect 47688 18204 47716 18300
rect 48314 18232 48320 18284
rect 48372 18281 48378 18284
rect 48372 18275 48421 18281
rect 48372 18241 48375 18275
rect 48409 18241 48421 18275
rect 48372 18235 48421 18241
rect 48372 18232 48378 18235
rect 52546 18232 52552 18284
rect 52604 18272 52610 18284
rect 52604 18244 53604 18272
rect 52604 18232 52610 18244
rect 48227 18207 48285 18213
rect 48227 18204 48239 18207
rect 46523 18176 46612 18204
rect 47688 18176 48239 18204
rect 46523 18173 46535 18176
rect 46477 18167 46535 18173
rect 39531 18108 40172 18136
rect 42245 18139 42303 18145
rect 39531 18105 39543 18108
rect 39485 18099 39543 18105
rect 42245 18105 42257 18139
rect 42291 18136 42303 18139
rect 43254 18136 43260 18148
rect 42291 18108 43260 18136
rect 42291 18105 42303 18108
rect 42245 18099 42303 18105
rect 43254 18096 43260 18108
rect 43312 18136 43318 18148
rect 43824 18136 43852 18167
rect 43312 18108 43852 18136
rect 43312 18096 43318 18108
rect 46584 18080 46612 18176
rect 48227 18173 48239 18176
rect 48273 18173 48285 18207
rect 48227 18167 48285 18173
rect 48498 18164 48504 18216
rect 48556 18164 48562 18216
rect 48774 18164 48780 18216
rect 48832 18164 48838 18216
rect 49237 18207 49295 18213
rect 49237 18173 49249 18207
rect 49283 18173 49295 18207
rect 49237 18167 49295 18173
rect 46750 18096 46756 18148
rect 46808 18136 46814 18148
rect 47118 18136 47124 18148
rect 46808 18108 47124 18136
rect 46808 18096 46814 18108
rect 47118 18096 47124 18108
rect 47176 18096 47182 18148
rect 49252 18136 49280 18167
rect 49418 18164 49424 18216
rect 49476 18164 49482 18216
rect 50893 18207 50951 18213
rect 50893 18173 50905 18207
rect 50939 18204 50951 18207
rect 51166 18204 51172 18216
rect 50939 18176 51172 18204
rect 50939 18173 50951 18176
rect 50893 18167 50951 18173
rect 51166 18164 51172 18176
rect 51224 18164 51230 18216
rect 52822 18164 52828 18216
rect 52880 18164 52886 18216
rect 53576 18204 53604 18244
rect 54570 18232 54576 18284
rect 54628 18232 54634 18284
rect 55600 18281 55628 18312
rect 56128 18309 56140 18343
rect 56174 18340 56186 18343
rect 56226 18340 56232 18352
rect 56174 18312 56232 18340
rect 56174 18309 56186 18312
rect 56128 18303 56186 18309
rect 56226 18300 56232 18312
rect 56284 18300 56290 18352
rect 55585 18275 55643 18281
rect 55585 18241 55597 18275
rect 55631 18241 55643 18275
rect 55585 18235 55643 18241
rect 55769 18275 55827 18281
rect 55769 18241 55781 18275
rect 55815 18272 55827 18275
rect 56888 18272 56916 18380
rect 57238 18368 57244 18380
rect 57296 18368 57302 18420
rect 55815 18244 56916 18272
rect 55815 18241 55827 18244
rect 55769 18235 55827 18241
rect 54711 18207 54769 18213
rect 54711 18204 54723 18207
rect 53576 18176 54723 18204
rect 54711 18173 54723 18176
rect 54757 18173 54769 18207
rect 54711 18167 54769 18173
rect 54846 18164 54852 18216
rect 54904 18164 54910 18216
rect 55861 18207 55919 18213
rect 55861 18173 55873 18207
rect 55907 18173 55919 18207
rect 55861 18167 55919 18173
rect 52840 18136 52868 18164
rect 53745 18139 53803 18145
rect 53745 18136 53757 18139
rect 49252 18108 49556 18136
rect 52840 18108 53757 18136
rect 37608 18040 38332 18068
rect 37608 18028 37614 18040
rect 39574 18028 39580 18080
rect 39632 18028 39638 18080
rect 42518 18028 42524 18080
rect 42576 18068 42582 18080
rect 45830 18068 45836 18080
rect 42576 18040 45836 18068
rect 42576 18028 42582 18040
rect 45830 18028 45836 18040
rect 45888 18028 45894 18080
rect 46566 18028 46572 18080
rect 46624 18068 46630 18080
rect 49528 18077 49556 18108
rect 53745 18105 53757 18108
rect 53791 18105 53803 18139
rect 53745 18099 53803 18105
rect 55125 18139 55183 18145
rect 55125 18105 55137 18139
rect 55171 18105 55183 18139
rect 55125 18099 55183 18105
rect 47305 18071 47363 18077
rect 47305 18068 47317 18071
rect 46624 18040 47317 18068
rect 46624 18028 46630 18040
rect 47305 18037 47317 18040
rect 47351 18037 47363 18071
rect 47305 18031 47363 18037
rect 49513 18071 49571 18077
rect 49513 18037 49525 18071
rect 49559 18068 49571 18071
rect 50706 18068 50712 18080
rect 49559 18040 50712 18068
rect 49559 18037 49571 18040
rect 49513 18031 49571 18037
rect 50706 18028 50712 18040
rect 50764 18028 50770 18080
rect 54386 18028 54392 18080
rect 54444 18068 54450 18080
rect 55140 18068 55168 18099
rect 54444 18040 55168 18068
rect 55876 18068 55904 18167
rect 57698 18164 57704 18216
rect 57756 18204 57762 18216
rect 58437 18207 58495 18213
rect 58437 18204 58449 18207
rect 57756 18176 58449 18204
rect 57756 18164 57762 18176
rect 58437 18173 58449 18176
rect 58483 18173 58495 18207
rect 58437 18167 58495 18173
rect 56134 18068 56140 18080
rect 55876 18040 56140 18068
rect 54444 18028 54450 18040
rect 56134 18028 56140 18040
rect 56192 18028 56198 18080
rect 57330 18028 57336 18080
rect 57388 18068 57394 18080
rect 57885 18071 57943 18077
rect 57885 18068 57897 18071
rect 57388 18040 57897 18068
rect 57388 18028 57394 18040
rect 57885 18037 57897 18040
rect 57931 18037 57943 18071
rect 57885 18031 57943 18037
rect 1104 17978 58880 18000
rect 1104 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 22616 17978
rect 22668 17926 22680 17978
rect 22732 17926 22744 17978
rect 22796 17926 22808 17978
rect 22860 17926 22872 17978
rect 22924 17926 37060 17978
rect 37112 17926 37124 17978
rect 37176 17926 37188 17978
rect 37240 17926 37252 17978
rect 37304 17926 37316 17978
rect 37368 17926 51504 17978
rect 51556 17926 51568 17978
rect 51620 17926 51632 17978
rect 51684 17926 51696 17978
rect 51748 17926 51760 17978
rect 51812 17926 58880 17978
rect 1104 17904 58880 17926
rect 3789 17867 3847 17873
rect 3789 17833 3801 17867
rect 3835 17864 3847 17867
rect 4154 17864 4160 17876
rect 3835 17836 4160 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 5905 17867 5963 17873
rect 5905 17833 5917 17867
rect 5951 17864 5963 17867
rect 6362 17864 6368 17876
rect 5951 17836 6368 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 9582 17864 9588 17876
rect 8720 17836 9588 17864
rect 8720 17824 8726 17836
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 9674 17824 9680 17876
rect 9732 17824 9738 17876
rect 9766 17824 9772 17876
rect 9824 17824 9830 17876
rect 12434 17824 12440 17876
rect 12492 17824 12498 17876
rect 14090 17824 14096 17876
rect 14148 17824 14154 17876
rect 14829 17867 14887 17873
rect 14829 17833 14841 17867
rect 14875 17864 14887 17867
rect 14918 17864 14924 17876
rect 14875 17836 14924 17864
rect 14875 17833 14887 17836
rect 14829 17827 14887 17833
rect 14918 17824 14924 17836
rect 14976 17824 14982 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 18104 17836 18429 17864
rect 18104 17824 18110 17836
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 20165 17867 20223 17873
rect 20165 17833 20177 17867
rect 20211 17864 20223 17867
rect 20254 17864 20260 17876
rect 20211 17836 20260 17864
rect 20211 17833 20223 17836
rect 20165 17827 20223 17833
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 23842 17864 23848 17876
rect 20772 17836 23848 17864
rect 20772 17824 20778 17836
rect 23842 17824 23848 17836
rect 23900 17824 23906 17876
rect 24213 17867 24271 17873
rect 24213 17833 24225 17867
rect 24259 17864 24271 17867
rect 25590 17864 25596 17876
rect 24259 17836 25596 17864
rect 24259 17833 24271 17836
rect 24213 17827 24271 17833
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 25774 17824 25780 17876
rect 25832 17824 25838 17876
rect 28445 17867 28503 17873
rect 28445 17833 28457 17867
rect 28491 17864 28503 17867
rect 28902 17864 28908 17876
rect 28491 17836 28908 17864
rect 28491 17833 28503 17836
rect 28445 17827 28503 17833
rect 28902 17824 28908 17836
rect 28960 17824 28966 17876
rect 33689 17867 33747 17873
rect 33689 17833 33701 17867
rect 33735 17864 33747 17867
rect 34238 17864 34244 17876
rect 33735 17836 34244 17864
rect 33735 17833 33747 17836
rect 33689 17827 33747 17833
rect 34238 17824 34244 17836
rect 34296 17824 34302 17876
rect 38654 17864 38660 17876
rect 38212 17836 38660 17864
rect 7300 17768 10272 17796
rect 7300 17740 7328 17768
rect 10244 17740 10272 17768
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 4212 17700 4353 17728
rect 4212 17688 4218 17700
rect 4341 17697 4353 17700
rect 4387 17728 4399 17731
rect 5261 17731 5319 17737
rect 4387 17700 5212 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 3510 17620 3516 17672
rect 3568 17620 3574 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4430 17660 4436 17672
rect 4295 17632 4436 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 5184 17660 5212 17700
rect 5261 17697 5273 17731
rect 5307 17728 5319 17731
rect 5442 17728 5448 17740
rect 5307 17700 5448 17728
rect 5307 17697 5319 17700
rect 5261 17691 5319 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 9122 17688 9128 17740
rect 9180 17688 9186 17740
rect 9674 17688 9680 17740
rect 9732 17688 9738 17740
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10284 17700 10517 17728
rect 10284 17688 10290 17700
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 12452 17728 12480 17824
rect 13909 17799 13967 17805
rect 13909 17765 13921 17799
rect 13955 17765 13967 17799
rect 13909 17759 13967 17765
rect 18325 17799 18383 17805
rect 18325 17765 18337 17799
rect 18371 17765 18383 17799
rect 18325 17759 18383 17765
rect 23492 17768 24440 17796
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 12452 17700 12541 17728
rect 10505 17691 10563 17697
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 13924 17728 13952 17759
rect 14458 17728 14464 17740
rect 13924 17700 14464 17728
rect 12529 17691 12587 17697
rect 14458 17688 14464 17700
rect 14516 17728 14522 17740
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 14516 17700 14657 17728
rect 14516 17688 14522 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 14792 17700 15393 17728
rect 14792 17688 14798 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 16206 17688 16212 17740
rect 16264 17688 16270 17740
rect 16942 17688 16948 17740
rect 17000 17688 17006 17740
rect 18340 17728 18368 17759
rect 23492 17740 23520 17768
rect 19061 17731 19119 17737
rect 19061 17728 19073 17731
rect 18340 17700 19073 17728
rect 19061 17697 19073 17700
rect 19107 17728 19119 17731
rect 20530 17728 20536 17740
rect 19107 17700 20536 17728
rect 19107 17697 19119 17700
rect 19061 17691 19119 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 23474 17728 23480 17740
rect 21652 17700 23480 17728
rect 5184 17632 5672 17660
rect 5644 17601 5672 17632
rect 7006 17620 7012 17672
rect 7064 17669 7070 17672
rect 7064 17660 7076 17669
rect 9309 17663 9367 17669
rect 7064 17632 7109 17660
rect 7064 17623 7076 17632
rect 9309 17629 9321 17663
rect 9355 17660 9367 17663
rect 9490 17660 9496 17672
rect 9355 17632 9496 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 7064 17620 7070 17623
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 9692 17660 9720 17688
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 9692 17632 10333 17660
rect 10321 17629 10333 17632
rect 10367 17629 10379 17663
rect 10321 17623 10379 17629
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10761 17663 10819 17669
rect 10761 17660 10773 17663
rect 10468 17632 10773 17660
rect 10468 17620 10474 17632
rect 10761 17629 10773 17632
rect 10807 17629 10819 17663
rect 10761 17623 10819 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12618 17660 12624 17672
rect 12483 17632 12624 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12618 17620 12624 17632
rect 12676 17660 12682 17672
rect 13262 17660 13268 17672
rect 12676 17632 13268 17660
rect 12676 17620 12682 17632
rect 13262 17620 13268 17632
rect 13320 17660 13326 17672
rect 13320 17632 13492 17660
rect 13320 17620 13326 17632
rect 13464 17604 13492 17632
rect 15286 17620 15292 17672
rect 15344 17620 15350 17672
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 21652 17669 21680 17700
rect 23474 17688 23480 17700
rect 23532 17688 23538 17740
rect 24412 17737 24440 17768
rect 35986 17756 35992 17808
rect 36044 17796 36050 17808
rect 37185 17799 37243 17805
rect 37185 17796 37197 17799
rect 36044 17768 37197 17796
rect 36044 17756 36050 17768
rect 37185 17765 37197 17768
rect 37231 17796 37243 17799
rect 37918 17796 37924 17808
rect 37231 17768 37924 17796
rect 37231 17765 37243 17768
rect 37185 17759 37243 17765
rect 37918 17756 37924 17768
rect 37976 17796 37982 17808
rect 38105 17799 38163 17805
rect 38105 17796 38117 17799
rect 37976 17768 38117 17796
rect 37976 17756 37982 17768
rect 38105 17765 38117 17768
rect 38151 17765 38163 17799
rect 38105 17759 38163 17765
rect 24397 17731 24455 17737
rect 24397 17697 24409 17731
rect 24443 17697 24455 17731
rect 27062 17728 27068 17740
rect 24397 17691 24455 17697
rect 25700 17700 27068 17728
rect 21637 17663 21695 17669
rect 21637 17660 21649 17663
rect 20864 17632 21649 17660
rect 20864 17620 20870 17632
rect 21637 17629 21649 17632
rect 21683 17629 21695 17663
rect 21637 17623 21695 17629
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22152 17632 22293 17660
rect 22152 17620 22158 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 24412 17660 24440 17691
rect 25700 17660 25728 17700
rect 27062 17688 27068 17700
rect 27120 17688 27126 17740
rect 29730 17688 29736 17740
rect 29788 17728 29794 17740
rect 30193 17731 30251 17737
rect 30193 17728 30205 17731
rect 29788 17700 30205 17728
rect 29788 17688 29794 17700
rect 30193 17697 30205 17700
rect 30239 17697 30251 17731
rect 30193 17691 30251 17697
rect 24412 17632 25728 17660
rect 22281 17623 22339 17629
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 25832 17632 26433 17660
rect 25832 17620 25838 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 27332 17663 27390 17669
rect 27332 17629 27344 17663
rect 27378 17660 27390 17663
rect 28258 17660 28264 17672
rect 27378 17632 28264 17660
rect 27378 17629 27390 17632
rect 27332 17623 27390 17629
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 30208 17660 30236 17691
rect 33778 17688 33784 17740
rect 33836 17688 33842 17740
rect 34422 17688 34428 17740
rect 34480 17728 34486 17740
rect 34793 17731 34851 17737
rect 34793 17728 34805 17731
rect 34480 17700 34805 17728
rect 34480 17688 34486 17700
rect 34793 17697 34805 17700
rect 34839 17697 34851 17731
rect 34793 17691 34851 17697
rect 37461 17731 37519 17737
rect 37461 17697 37473 17731
rect 37507 17728 37519 17731
rect 37734 17728 37740 17740
rect 37507 17700 37740 17728
rect 37507 17697 37519 17700
rect 37461 17691 37519 17697
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 38212 17728 38240 17836
rect 38654 17824 38660 17836
rect 38712 17824 38718 17876
rect 44821 17867 44879 17873
rect 44821 17833 44833 17867
rect 44867 17864 44879 17867
rect 45002 17864 45008 17876
rect 44867 17836 45008 17864
rect 44867 17833 44879 17836
rect 44821 17827 44879 17833
rect 45002 17824 45008 17836
rect 45060 17824 45066 17876
rect 46014 17824 46020 17876
rect 46072 17864 46078 17876
rect 46477 17867 46535 17873
rect 46477 17864 46489 17867
rect 46072 17836 46489 17864
rect 46072 17824 46078 17836
rect 46477 17833 46489 17836
rect 46523 17833 46535 17867
rect 48498 17864 48504 17876
rect 46477 17827 46535 17833
rect 47136 17836 48504 17864
rect 42610 17756 42616 17808
rect 42668 17796 42674 17808
rect 42705 17799 42763 17805
rect 42705 17796 42717 17799
rect 42668 17768 42717 17796
rect 42668 17756 42674 17768
rect 42705 17765 42717 17768
rect 42751 17796 42763 17799
rect 45020 17796 45048 17824
rect 42751 17768 45048 17796
rect 42751 17765 42763 17768
rect 42705 17759 42763 17765
rect 38381 17731 38439 17737
rect 38381 17728 38393 17731
rect 38212 17700 38393 17728
rect 38381 17697 38393 17700
rect 38427 17697 38439 17731
rect 38381 17691 38439 17697
rect 38657 17731 38715 17737
rect 38657 17697 38669 17731
rect 38703 17728 38715 17731
rect 38703 17700 39252 17728
rect 38703 17697 38715 17700
rect 38657 17691 38715 17697
rect 32309 17663 32367 17669
rect 32309 17660 32321 17663
rect 30208 17632 32321 17660
rect 31956 17604 31984 17632
rect 32309 17629 32321 17632
rect 32355 17629 32367 17663
rect 33796 17660 33824 17688
rect 34977 17663 35035 17669
rect 34977 17660 34989 17663
rect 33796 17632 34989 17660
rect 32309 17623 32367 17629
rect 34977 17629 34989 17632
rect 35023 17629 35035 17663
rect 34977 17623 35035 17629
rect 37642 17620 37648 17672
rect 37700 17620 37706 17672
rect 38470 17620 38476 17672
rect 38528 17669 38534 17672
rect 38528 17663 38556 17669
rect 38544 17629 38556 17663
rect 38528 17623 38556 17629
rect 38528 17620 38534 17623
rect 4157 17595 4215 17601
rect 4157 17561 4169 17595
rect 4203 17592 4215 17595
rect 4617 17595 4675 17601
rect 4617 17592 4629 17595
rect 4203 17564 4629 17592
rect 4203 17561 4215 17564
rect 4157 17555 4215 17561
rect 4617 17561 4629 17564
rect 4663 17561 4675 17595
rect 4617 17555 4675 17561
rect 5629 17595 5687 17601
rect 5629 17561 5641 17595
rect 5675 17592 5687 17595
rect 12526 17592 12532 17604
rect 5675 17564 9352 17592
rect 5675 17561 5687 17564
rect 5629 17555 5687 17561
rect 2958 17484 2964 17536
rect 3016 17484 3022 17536
rect 8294 17484 8300 17536
rect 8352 17484 8358 17536
rect 9214 17484 9220 17536
rect 9272 17484 9278 17536
rect 9324 17524 9352 17564
rect 12406 17564 12532 17592
rect 9674 17524 9680 17536
rect 9324 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 11885 17527 11943 17533
rect 11885 17493 11897 17527
rect 11931 17524 11943 17527
rect 12406 17524 12434 17564
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 12796 17595 12854 17601
rect 12796 17561 12808 17595
rect 12842 17592 12854 17595
rect 12986 17592 12992 17604
rect 12842 17564 12992 17592
rect 12842 17561 12854 17564
rect 12796 17555 12854 17561
rect 12986 17552 12992 17564
rect 13044 17552 13050 17604
rect 13446 17552 13452 17604
rect 13504 17552 13510 17604
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17592 15255 17595
rect 15657 17595 15715 17601
rect 15657 17592 15669 17595
rect 15243 17564 15669 17592
rect 15243 17561 15255 17564
rect 15197 17555 15255 17561
rect 15657 17561 15669 17564
rect 15703 17561 15715 17595
rect 15657 17555 15715 17561
rect 17212 17595 17270 17601
rect 17212 17561 17224 17595
rect 17258 17592 17270 17595
rect 17402 17592 17408 17604
rect 17258 17564 17408 17592
rect 17258 17561 17270 17564
rect 17212 17555 17270 17561
rect 17402 17552 17408 17564
rect 17460 17552 17466 17604
rect 21392 17595 21450 17601
rect 21392 17561 21404 17595
rect 21438 17592 21450 17595
rect 22186 17592 22192 17604
rect 21438 17564 22192 17592
rect 21438 17561 21450 17564
rect 21392 17555 21450 17561
rect 22186 17552 22192 17564
rect 22244 17552 22250 17604
rect 24664 17595 24722 17601
rect 24664 17561 24676 17595
rect 24710 17592 24722 17595
rect 25038 17592 25044 17604
rect 24710 17564 25044 17592
rect 24710 17561 24722 17564
rect 24664 17555 24722 17561
rect 25038 17552 25044 17564
rect 25096 17552 25102 17604
rect 26142 17592 26148 17604
rect 25148 17564 26148 17592
rect 11931 17496 12434 17524
rect 20257 17527 20315 17533
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 21266 17524 21272 17536
rect 20303 17496 21272 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 21726 17484 21732 17536
rect 21784 17484 21790 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 24854 17524 24860 17536
rect 23900 17496 24860 17524
rect 23900 17484 23906 17496
rect 24854 17484 24860 17496
rect 24912 17524 24918 17536
rect 25148 17524 25176 17564
rect 26142 17552 26148 17564
rect 26200 17592 26206 17604
rect 26878 17592 26884 17604
rect 26200 17564 26884 17592
rect 26200 17552 26206 17564
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 30460 17595 30518 17601
rect 30460 17561 30472 17595
rect 30506 17592 30518 17595
rect 31018 17592 31024 17604
rect 30506 17564 31024 17592
rect 30506 17561 30518 17564
rect 30460 17555 30518 17561
rect 31018 17552 31024 17564
rect 31076 17552 31082 17604
rect 31849 17595 31907 17601
rect 31849 17561 31861 17595
rect 31895 17592 31907 17595
rect 31938 17592 31944 17604
rect 31895 17564 31944 17592
rect 31895 17561 31907 17564
rect 31849 17555 31907 17561
rect 31938 17552 31944 17564
rect 31996 17552 32002 17604
rect 32576 17595 32634 17601
rect 32576 17561 32588 17595
rect 32622 17592 32634 17595
rect 32858 17592 32864 17604
rect 32622 17564 32864 17592
rect 32622 17561 32634 17564
rect 32576 17555 32634 17561
rect 32858 17552 32864 17564
rect 32916 17552 32922 17604
rect 32950 17552 32956 17604
rect 33008 17592 33014 17604
rect 33008 17564 34652 17592
rect 33008 17552 33014 17564
rect 24912 17496 25176 17524
rect 24912 17484 24918 17496
rect 25866 17484 25872 17536
rect 25924 17484 25930 17536
rect 28718 17484 28724 17536
rect 28776 17524 28782 17536
rect 29178 17524 29184 17536
rect 28776 17496 29184 17524
rect 28776 17484 28782 17496
rect 29178 17484 29184 17496
rect 29236 17484 29242 17536
rect 31573 17527 31631 17533
rect 31573 17493 31585 17527
rect 31619 17524 31631 17527
rect 33410 17524 33416 17536
rect 31619 17496 33416 17524
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 33410 17484 33416 17496
rect 33468 17484 33474 17536
rect 33965 17527 34023 17533
rect 33965 17493 33977 17527
rect 34011 17524 34023 17527
rect 34514 17524 34520 17536
rect 34011 17496 34520 17524
rect 34011 17493 34023 17496
rect 33965 17487 34023 17493
rect 34514 17484 34520 17496
rect 34572 17484 34578 17536
rect 34624 17524 34652 17564
rect 34698 17552 34704 17604
rect 34756 17592 34762 17604
rect 35069 17595 35127 17601
rect 35069 17592 35081 17595
rect 34756 17564 35081 17592
rect 34756 17552 34762 17564
rect 35069 17561 35081 17564
rect 35115 17561 35127 17595
rect 36722 17592 36728 17604
rect 35069 17555 35127 17561
rect 35167 17564 36728 17592
rect 35167 17524 35195 17564
rect 36722 17552 36728 17564
rect 36780 17552 36786 17604
rect 34624 17496 35195 17524
rect 35434 17484 35440 17536
rect 35492 17484 35498 17536
rect 36740 17524 36768 17552
rect 39224 17524 39252 17700
rect 45020 17669 45048 17768
rect 46385 17799 46443 17805
rect 46385 17765 46397 17799
rect 46431 17796 46443 17799
rect 47136 17796 47164 17836
rect 48498 17824 48504 17836
rect 48556 17824 48562 17876
rect 48685 17867 48743 17873
rect 48685 17833 48697 17867
rect 48731 17864 48743 17867
rect 49418 17864 49424 17876
rect 48731 17836 49424 17864
rect 48731 17833 48743 17836
rect 48685 17827 48743 17833
rect 49418 17824 49424 17836
rect 49476 17824 49482 17876
rect 49881 17867 49939 17873
rect 49881 17833 49893 17867
rect 49927 17864 49939 17867
rect 50338 17864 50344 17876
rect 49927 17836 50344 17864
rect 49927 17833 49939 17836
rect 49881 17827 49939 17833
rect 50338 17824 50344 17836
rect 50396 17824 50402 17876
rect 52730 17824 52736 17876
rect 52788 17864 52794 17876
rect 53101 17867 53159 17873
rect 53101 17864 53113 17867
rect 52788 17836 53113 17864
rect 52788 17824 52794 17836
rect 53101 17833 53113 17836
rect 53147 17833 53159 17867
rect 53101 17827 53159 17833
rect 54113 17867 54171 17873
rect 54113 17833 54125 17867
rect 54159 17864 54171 17867
rect 54294 17864 54300 17876
rect 54159 17836 54300 17864
rect 54159 17833 54171 17836
rect 54113 17827 54171 17833
rect 54294 17824 54300 17836
rect 54352 17824 54358 17876
rect 56045 17867 56103 17873
rect 56045 17833 56057 17867
rect 56091 17864 56103 17867
rect 56594 17864 56600 17876
rect 56091 17836 56600 17864
rect 56091 17833 56103 17836
rect 56045 17827 56103 17833
rect 56594 17824 56600 17836
rect 56652 17824 56658 17876
rect 56686 17824 56692 17876
rect 56744 17864 56750 17876
rect 57698 17864 57704 17876
rect 56744 17836 57704 17864
rect 56744 17824 56750 17836
rect 57698 17824 57704 17836
rect 57756 17824 57762 17876
rect 46431 17768 47164 17796
rect 46431 17765 46443 17768
rect 46385 17759 46443 17765
rect 47136 17737 47164 17768
rect 53009 17799 53067 17805
rect 53009 17765 53021 17799
rect 53055 17796 53067 17799
rect 53055 17768 53788 17796
rect 53055 17765 53067 17768
rect 53009 17759 53067 17765
rect 47121 17731 47179 17737
rect 47121 17697 47133 17731
rect 47167 17697 47179 17731
rect 49237 17731 49295 17737
rect 49237 17728 49249 17731
rect 47121 17691 47179 17697
rect 48976 17700 49249 17728
rect 45278 17669 45284 17672
rect 45005 17663 45063 17669
rect 45005 17629 45017 17663
rect 45051 17629 45063 17663
rect 45272 17660 45284 17669
rect 45239 17632 45284 17660
rect 45005 17623 45063 17629
rect 45272 17623 45284 17632
rect 45278 17620 45284 17623
rect 45336 17620 45342 17672
rect 47305 17663 47363 17669
rect 47305 17629 47317 17663
rect 47351 17660 47363 17663
rect 47394 17660 47400 17672
rect 47351 17632 47400 17660
rect 47351 17629 47363 17632
rect 47305 17623 47363 17629
rect 47394 17620 47400 17632
rect 47452 17620 47458 17672
rect 48590 17620 48596 17672
rect 48648 17620 48654 17672
rect 47572 17595 47630 17601
rect 47572 17561 47584 17595
rect 47618 17592 47630 17595
rect 47762 17592 47768 17604
rect 47618 17564 47768 17592
rect 47618 17561 47630 17564
rect 47572 17555 47630 17561
rect 47762 17552 47768 17564
rect 47820 17552 47826 17604
rect 36740 17496 39252 17524
rect 39298 17484 39304 17536
rect 39356 17484 39362 17536
rect 42337 17527 42395 17533
rect 42337 17493 42349 17527
rect 42383 17524 42395 17527
rect 42518 17524 42524 17536
rect 42383 17496 42524 17524
rect 42383 17493 42395 17496
rect 42337 17487 42395 17493
rect 42518 17484 42524 17496
rect 42576 17524 42582 17536
rect 42702 17524 42708 17536
rect 42576 17496 42708 17524
rect 42576 17484 42582 17496
rect 42702 17484 42708 17496
rect 42760 17484 42766 17536
rect 43257 17527 43315 17533
rect 43257 17493 43269 17527
rect 43303 17524 43315 17527
rect 43438 17524 43444 17536
rect 43303 17496 43444 17524
rect 43303 17493 43315 17496
rect 43257 17487 43315 17493
rect 43438 17484 43444 17496
rect 43496 17524 43502 17536
rect 48608 17524 48636 17620
rect 43496 17496 48636 17524
rect 43496 17484 43502 17496
rect 48774 17484 48780 17536
rect 48832 17524 48838 17536
rect 48976 17533 49004 17700
rect 49237 17697 49249 17700
rect 49283 17697 49295 17731
rect 49237 17691 49295 17697
rect 50706 17688 50712 17740
rect 50764 17688 50770 17740
rect 53760 17737 53788 17768
rect 53745 17731 53803 17737
rect 53745 17697 53757 17731
rect 53791 17728 53803 17731
rect 54846 17728 54852 17740
rect 53791 17700 54852 17728
rect 53791 17697 53803 17700
rect 53745 17691 53803 17697
rect 54846 17688 54852 17700
rect 54904 17688 54910 17740
rect 55401 17731 55459 17737
rect 55401 17728 55413 17731
rect 55048 17700 55413 17728
rect 51166 17620 51172 17672
rect 51224 17660 51230 17672
rect 51629 17663 51687 17669
rect 51629 17660 51641 17663
rect 51224 17632 51641 17660
rect 51224 17620 51230 17632
rect 51629 17629 51641 17632
rect 51675 17660 51687 17663
rect 51675 17632 52040 17660
rect 51675 17629 51687 17632
rect 51629 17623 51687 17629
rect 51902 17601 51908 17604
rect 49513 17595 49571 17601
rect 49513 17561 49525 17595
rect 49559 17592 49571 17595
rect 50157 17595 50215 17601
rect 50157 17592 50169 17595
rect 49559 17564 50169 17592
rect 49559 17561 49571 17564
rect 49513 17555 49571 17561
rect 50157 17561 50169 17564
rect 50203 17561 50215 17595
rect 51896 17592 51908 17601
rect 51863 17564 51908 17592
rect 50157 17555 50215 17561
rect 51896 17555 51908 17564
rect 51902 17552 51908 17555
rect 51960 17552 51966 17604
rect 52012 17536 52040 17632
rect 48961 17527 49019 17533
rect 48961 17524 48973 17527
rect 48832 17496 48973 17524
rect 48832 17484 48838 17496
rect 48961 17493 48973 17496
rect 49007 17493 49019 17527
rect 48961 17487 49019 17493
rect 49326 17484 49332 17536
rect 49384 17524 49390 17536
rect 49421 17527 49479 17533
rect 49421 17524 49433 17527
rect 49384 17496 49433 17524
rect 49384 17484 49390 17496
rect 49421 17493 49433 17496
rect 49467 17524 49479 17527
rect 49878 17524 49884 17536
rect 49467 17496 49884 17524
rect 49467 17493 49479 17496
rect 49421 17487 49479 17493
rect 49878 17484 49884 17496
rect 49936 17484 49942 17536
rect 51994 17484 52000 17536
rect 52052 17484 52058 17536
rect 54294 17484 54300 17536
rect 54352 17524 54358 17536
rect 55048 17533 55076 17700
rect 55401 17697 55413 17700
rect 55447 17697 55459 17731
rect 55401 17691 55459 17697
rect 55585 17731 55643 17737
rect 55585 17697 55597 17731
rect 55631 17728 55643 17731
rect 55631 17700 56456 17728
rect 55631 17697 55643 17700
rect 55585 17691 55643 17697
rect 56134 17620 56140 17672
rect 56192 17660 56198 17672
rect 56321 17663 56379 17669
rect 56321 17660 56333 17663
rect 56192 17632 56333 17660
rect 56192 17620 56198 17632
rect 56321 17629 56333 17632
rect 56367 17629 56379 17663
rect 56428 17660 56456 17700
rect 56962 17660 56968 17672
rect 56428 17632 56968 17660
rect 56321 17623 56379 17629
rect 56962 17620 56968 17632
rect 57020 17620 57026 17672
rect 58342 17620 58348 17672
rect 58400 17620 58406 17672
rect 56588 17595 56646 17601
rect 56588 17561 56600 17595
rect 56634 17592 56646 17595
rect 57793 17595 57851 17601
rect 57793 17592 57805 17595
rect 56634 17564 57805 17592
rect 56634 17561 56646 17564
rect 56588 17555 56646 17561
rect 57793 17561 57805 17564
rect 57839 17561 57851 17595
rect 57793 17555 57851 17561
rect 55033 17527 55091 17533
rect 55033 17524 55045 17527
rect 54352 17496 55045 17524
rect 54352 17484 54358 17496
rect 55033 17493 55045 17496
rect 55079 17493 55091 17527
rect 55033 17487 55091 17493
rect 55674 17484 55680 17536
rect 55732 17484 55738 17536
rect 1104 17434 59040 17456
rect 1104 17382 15394 17434
rect 15446 17382 15458 17434
rect 15510 17382 15522 17434
rect 15574 17382 15586 17434
rect 15638 17382 15650 17434
rect 15702 17382 29838 17434
rect 29890 17382 29902 17434
rect 29954 17382 29966 17434
rect 30018 17382 30030 17434
rect 30082 17382 30094 17434
rect 30146 17382 44282 17434
rect 44334 17382 44346 17434
rect 44398 17382 44410 17434
rect 44462 17382 44474 17434
rect 44526 17382 44538 17434
rect 44590 17382 58726 17434
rect 58778 17382 58790 17434
rect 58842 17382 58854 17434
rect 58906 17382 58918 17434
rect 58970 17382 58982 17434
rect 59034 17382 59040 17434
rect 1104 17360 59040 17382
rect 3329 17323 3387 17329
rect 3329 17289 3341 17323
rect 3375 17320 3387 17323
rect 3510 17320 3516 17332
rect 3375 17292 3516 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 7282 17320 7288 17332
rect 6871 17292 7288 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9398 17320 9404 17332
rect 9263 17292 9404 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 12986 17280 12992 17332
rect 13044 17280 13050 17332
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 17402 17280 17408 17332
rect 17460 17280 17466 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 19668 17292 20545 17320
rect 19668 17280 19674 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20533 17283 20591 17289
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21726 17320 21732 17332
rect 21039 17292 21732 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21726 17280 21732 17292
rect 21784 17280 21790 17332
rect 22097 17323 22155 17329
rect 22097 17289 22109 17323
rect 22143 17320 22155 17323
rect 22370 17320 22376 17332
rect 22143 17292 22376 17320
rect 22143 17289 22155 17292
rect 22097 17283 22155 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 25038 17280 25044 17332
rect 25096 17280 25102 17332
rect 25866 17280 25872 17332
rect 25924 17280 25930 17332
rect 26053 17323 26111 17329
rect 26053 17289 26065 17323
rect 26099 17320 26111 17323
rect 26602 17320 26608 17332
rect 26099 17292 26608 17320
rect 26099 17289 26111 17292
rect 26053 17283 26111 17289
rect 26602 17280 26608 17292
rect 26660 17320 26666 17332
rect 28166 17320 28172 17332
rect 26660 17292 28172 17320
rect 26660 17280 26666 17292
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 31018 17280 31024 17332
rect 31076 17280 31082 17332
rect 32030 17280 32036 17332
rect 32088 17320 32094 17332
rect 32125 17323 32183 17329
rect 32125 17320 32137 17323
rect 32088 17292 32137 17320
rect 32088 17280 32094 17292
rect 32125 17289 32137 17292
rect 32171 17289 32183 17323
rect 32125 17283 32183 17289
rect 32858 17280 32864 17332
rect 32916 17280 32922 17332
rect 37734 17280 37740 17332
rect 37792 17320 37798 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 37792 17292 37841 17320
rect 37792 17280 37798 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 37829 17283 37887 17289
rect 38838 17280 38844 17332
rect 38896 17280 38902 17332
rect 39298 17280 39304 17332
rect 39356 17320 39362 17332
rect 39761 17323 39819 17329
rect 39761 17320 39773 17323
rect 39356 17292 39773 17320
rect 39356 17280 39362 17292
rect 39761 17289 39773 17292
rect 39807 17289 39819 17323
rect 39761 17283 39819 17289
rect 43714 17280 43720 17332
rect 43772 17280 43778 17332
rect 47213 17323 47271 17329
rect 47213 17289 47225 17323
rect 47259 17320 47271 17323
rect 47394 17320 47400 17332
rect 47259 17292 47400 17320
rect 47259 17289 47271 17292
rect 47213 17283 47271 17289
rect 47394 17280 47400 17292
rect 47452 17280 47458 17332
rect 47762 17280 47768 17332
rect 47820 17280 47826 17332
rect 48501 17323 48559 17329
rect 48501 17289 48513 17323
rect 48547 17320 48559 17323
rect 48866 17320 48872 17332
rect 48547 17292 48872 17320
rect 48547 17289 48559 17292
rect 48501 17283 48559 17289
rect 48866 17280 48872 17292
rect 48924 17280 48930 17332
rect 57057 17323 57115 17329
rect 57057 17289 57069 17323
rect 57103 17320 57115 17323
rect 57330 17320 57336 17332
rect 57103 17292 57336 17320
rect 57103 17289 57115 17292
rect 57057 17283 57115 17289
rect 57330 17280 57336 17292
rect 57388 17280 57394 17332
rect 57425 17323 57483 17329
rect 57425 17289 57437 17323
rect 57471 17320 57483 17323
rect 58342 17320 58348 17332
rect 57471 17292 58348 17320
rect 57471 17289 57483 17292
rect 57425 17283 57483 17289
rect 58342 17280 58348 17292
rect 58400 17280 58406 17332
rect 3697 17255 3755 17261
rect 3697 17221 3709 17255
rect 3743 17252 3755 17255
rect 3970 17252 3976 17264
rect 3743 17224 3976 17252
rect 3743 17221 3755 17224
rect 3697 17215 3755 17221
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 9122 17212 9128 17264
rect 9180 17252 9186 17264
rect 9861 17255 9919 17261
rect 9861 17252 9873 17255
rect 9180 17224 9873 17252
rect 9180 17212 9186 17224
rect 9861 17221 9873 17224
rect 9907 17252 9919 17255
rect 14752 17252 14780 17280
rect 9907 17224 14780 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 19886 17212 19892 17264
rect 19944 17252 19950 17264
rect 24581 17255 24639 17261
rect 19944 17224 22094 17252
rect 19944 17212 19950 17224
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 3835 17156 4169 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8294 17184 8300 17196
rect 8159 17156 8300 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8294 17144 8300 17156
rect 8352 17184 8358 17196
rect 9766 17184 9772 17196
rect 8352 17156 9772 17184
rect 8352 17144 8358 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13228 17156 13553 17184
rect 13228 17144 13234 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 17954 17144 17960 17196
rect 18012 17144 18018 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 22066 17184 22094 17224
rect 24581 17221 24593 17255
rect 24627 17252 24639 17255
rect 25884 17252 25912 17280
rect 24627 17224 25912 17252
rect 24627 17221 24639 17224
rect 24581 17215 24639 17221
rect 25498 17184 25504 17196
rect 22066 17156 25504 17184
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 31570 17144 31576 17196
rect 31628 17144 31634 17196
rect 32769 17187 32827 17193
rect 32769 17153 32781 17187
rect 32815 17184 32827 17187
rect 33410 17184 33416 17196
rect 32815 17156 33416 17184
rect 32815 17153 32827 17156
rect 32769 17147 32827 17153
rect 33410 17144 33416 17156
rect 33468 17144 33474 17196
rect 33505 17187 33563 17193
rect 33505 17153 33517 17187
rect 33551 17184 33563 17187
rect 33594 17184 33600 17196
rect 33551 17156 33600 17184
rect 33551 17153 33563 17156
rect 33505 17147 33563 17153
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 38856 17184 38884 17280
rect 38964 17255 39022 17261
rect 38964 17221 38976 17255
rect 39010 17252 39022 17255
rect 39574 17252 39580 17264
rect 39010 17224 39580 17252
rect 39010 17221 39022 17224
rect 38964 17215 39022 17221
rect 39574 17212 39580 17224
rect 39632 17212 39638 17264
rect 39669 17187 39727 17193
rect 39669 17184 39681 17187
rect 38856 17156 39681 17184
rect 39669 17153 39681 17156
rect 39715 17153 39727 17187
rect 39669 17147 39727 17153
rect 39868 17156 43484 17184
rect 3234 17076 3240 17128
rect 3292 17076 3298 17128
rect 3973 17119 4031 17125
rect 3973 17085 3985 17119
rect 4019 17085 4031 17119
rect 3973 17079 4031 17085
rect 2590 16940 2596 16992
rect 2648 16940 2654 16992
rect 3988 16980 4016 17079
rect 4614 17076 4620 17128
rect 4672 17116 4678 17128
rect 4709 17119 4767 17125
rect 4709 17116 4721 17119
rect 4672 17088 4721 17116
rect 4672 17076 4678 17088
rect 4709 17085 4721 17088
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5316 17088 6193 17116
rect 5316 17076 5322 17088
rect 6181 17085 6193 17088
rect 6227 17116 6239 17119
rect 8662 17116 8668 17128
rect 6227 17088 8668 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8754 17076 8760 17128
rect 8812 17076 8818 17128
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20364 17088 21097 17116
rect 9214 17008 9220 17060
rect 9272 17048 9278 17060
rect 9950 17048 9956 17060
rect 9272 17020 9956 17048
rect 9272 17008 9278 17020
rect 9950 17008 9956 17020
rect 10008 17008 10014 17060
rect 20364 16992 20392 17088
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 21085 17079 21143 17085
rect 24136 17088 24317 17116
rect 24136 16992 24164 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 24305 17079 24363 17085
rect 24489 17119 24547 17125
rect 24489 17085 24501 17119
rect 24535 17116 24547 17119
rect 24762 17116 24768 17128
rect 24535 17088 24768 17116
rect 24535 17085 24547 17088
rect 24489 17079 24547 17085
rect 24762 17076 24768 17088
rect 24820 17116 24826 17128
rect 25130 17116 25136 17128
rect 24820 17088 25136 17116
rect 24820 17076 24826 17088
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 39868 17125 39896 17156
rect 43456 17128 43484 17156
rect 48406 17144 48412 17196
rect 48464 17144 48470 17196
rect 49145 17187 49203 17193
rect 49145 17153 49157 17187
rect 49191 17184 49203 17187
rect 49418 17184 49424 17196
rect 49191 17156 49424 17184
rect 49191 17153 49203 17156
rect 49145 17147 49203 17153
rect 49418 17144 49424 17156
rect 49476 17144 49482 17196
rect 25593 17119 25651 17125
rect 25593 17085 25605 17119
rect 25639 17085 25651 17119
rect 25593 17079 25651 17085
rect 39209 17119 39267 17125
rect 39209 17085 39221 17119
rect 39255 17085 39267 17119
rect 39209 17079 39267 17085
rect 39853 17119 39911 17125
rect 39853 17085 39865 17119
rect 39899 17085 39911 17119
rect 39853 17079 39911 17085
rect 24949 17051 25007 17057
rect 24949 17017 24961 17051
rect 24995 17048 25007 17051
rect 25608 17048 25636 17079
rect 24995 17020 25636 17048
rect 24995 17017 25007 17020
rect 24949 17011 25007 17017
rect 5166 16980 5172 16992
rect 3988 16952 5172 16980
rect 5166 16940 5172 16952
rect 5224 16980 5230 16992
rect 5994 16980 6000 16992
rect 5224 16952 6000 16980
rect 5224 16940 5230 16952
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 7098 16980 7104 16992
rect 6328 16952 7104 16980
rect 6328 16940 6334 16952
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7926 16940 7932 16992
rect 7984 16980 7990 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7984 16952 8217 16980
rect 7984 16940 7990 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12710 16980 12716 16992
rect 12483 16952 12716 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12710 16940 12716 16952
rect 12768 16980 12774 16992
rect 12986 16980 12992 16992
rect 12768 16952 12992 16980
rect 12768 16940 12774 16952
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 17586 16940 17592 16992
rect 17644 16980 17650 16992
rect 18322 16980 18328 16992
rect 17644 16952 18328 16980
rect 17644 16940 17650 16952
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 19337 16983 19395 16989
rect 19337 16949 19349 16983
rect 19383 16980 19395 16983
rect 19702 16980 19708 16992
rect 19383 16952 19708 16980
rect 19383 16949 19395 16952
rect 19337 16943 19395 16949
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 20346 16940 20352 16992
rect 20404 16940 20410 16992
rect 24118 16940 24124 16992
rect 24176 16940 24182 16992
rect 34333 16983 34391 16989
rect 34333 16949 34345 16983
rect 34379 16980 34391 16983
rect 34514 16980 34520 16992
rect 34379 16952 34520 16980
rect 34379 16949 34391 16952
rect 34333 16943 34391 16949
rect 34514 16940 34520 16952
rect 34572 16980 34578 16992
rect 35342 16980 35348 16992
rect 34572 16952 35348 16980
rect 34572 16940 34578 16952
rect 35342 16940 35348 16952
rect 35400 16980 35406 16992
rect 35529 16983 35587 16989
rect 35529 16980 35541 16983
rect 35400 16952 35541 16980
rect 35400 16940 35406 16952
rect 35529 16949 35541 16952
rect 35575 16980 35587 16983
rect 37001 16983 37059 16989
rect 37001 16980 37013 16983
rect 35575 16952 37013 16980
rect 35575 16949 35587 16952
rect 35529 16943 35587 16949
rect 37001 16949 37013 16952
rect 37047 16980 37059 16983
rect 37461 16983 37519 16989
rect 37461 16980 37473 16983
rect 37047 16952 37473 16980
rect 37047 16949 37059 16952
rect 37001 16943 37059 16949
rect 37461 16949 37473 16952
rect 37507 16980 37519 16983
rect 38838 16980 38844 16992
rect 37507 16952 38844 16980
rect 37507 16949 37519 16952
rect 37461 16943 37519 16949
rect 38838 16940 38844 16952
rect 38896 16980 38902 16992
rect 39224 16980 39252 17079
rect 39868 16992 39896 17079
rect 42978 17076 42984 17128
rect 43036 17076 43042 17128
rect 43438 17076 43444 17128
rect 43496 17076 43502 17128
rect 43622 17076 43628 17128
rect 43680 17076 43686 17128
rect 44266 17076 44272 17128
rect 44324 17076 44330 17128
rect 45557 17119 45615 17125
rect 45557 17085 45569 17119
rect 45603 17116 45615 17119
rect 45646 17116 45652 17128
rect 45603 17088 45652 17116
rect 45603 17085 45615 17088
rect 45557 17079 45615 17085
rect 45646 17076 45652 17088
rect 45704 17076 45710 17128
rect 56597 17119 56655 17125
rect 56597 17085 56609 17119
rect 56643 17116 56655 17119
rect 56870 17116 56876 17128
rect 56643 17088 56876 17116
rect 56643 17085 56655 17088
rect 56597 17079 56655 17085
rect 56870 17076 56876 17088
rect 56928 17076 56934 17128
rect 56965 17119 57023 17125
rect 56965 17085 56977 17119
rect 57011 17085 57023 17119
rect 56965 17079 57023 17085
rect 43990 17008 43996 17060
rect 44048 17048 44054 17060
rect 44913 17051 44971 17057
rect 44913 17048 44925 17051
rect 44048 17020 44925 17048
rect 44048 17008 44054 17020
rect 44913 17017 44925 17020
rect 44959 17017 44971 17051
rect 44913 17011 44971 17017
rect 55674 17008 55680 17060
rect 55732 17048 55738 17060
rect 56980 17048 57008 17079
rect 57698 17076 57704 17128
rect 57756 17116 57762 17128
rect 58437 17119 58495 17125
rect 58437 17116 58449 17119
rect 57756 17088 58449 17116
rect 57756 17076 57762 17088
rect 58437 17085 58449 17088
rect 58483 17085 58495 17119
rect 58437 17079 58495 17085
rect 58250 17048 58256 17060
rect 55732 17020 58256 17048
rect 55732 17008 55738 17020
rect 58250 17008 58256 17020
rect 58308 17008 58314 17060
rect 38896 16952 39252 16980
rect 38896 16940 38902 16952
rect 39298 16940 39304 16992
rect 39356 16940 39362 16992
rect 39850 16940 39856 16992
rect 39908 16940 39914 16992
rect 41598 16940 41604 16992
rect 41656 16980 41662 16992
rect 42334 16980 42340 16992
rect 41656 16952 42340 16980
rect 41656 16940 41662 16952
rect 42334 16940 42340 16952
rect 42392 16940 42398 16992
rect 42426 16940 42432 16992
rect 42484 16940 42490 16992
rect 44082 16940 44088 16992
rect 44140 16940 44146 16992
rect 44818 16940 44824 16992
rect 44876 16940 44882 16992
rect 53190 16940 53196 16992
rect 53248 16980 53254 16992
rect 53561 16983 53619 16989
rect 53561 16980 53573 16983
rect 53248 16952 53573 16980
rect 53248 16940 53254 16952
rect 53561 16949 53573 16952
rect 53607 16980 53619 16983
rect 55769 16983 55827 16989
rect 55769 16980 55781 16983
rect 53607 16952 55781 16980
rect 53607 16949 53619 16952
rect 53561 16943 53619 16949
rect 55769 16949 55781 16952
rect 55815 16980 55827 16983
rect 56134 16980 56140 16992
rect 55815 16952 56140 16980
rect 55815 16949 55827 16952
rect 55769 16943 55827 16949
rect 56134 16940 56140 16952
rect 56192 16940 56198 16992
rect 57882 16940 57888 16992
rect 57940 16940 57946 16992
rect 1104 16890 58880 16912
rect 1104 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 22616 16890
rect 22668 16838 22680 16890
rect 22732 16838 22744 16890
rect 22796 16838 22808 16890
rect 22860 16838 22872 16890
rect 22924 16838 37060 16890
rect 37112 16838 37124 16890
rect 37176 16838 37188 16890
rect 37240 16838 37252 16890
rect 37304 16838 37316 16890
rect 37368 16838 51504 16890
rect 51556 16838 51568 16890
rect 51620 16838 51632 16890
rect 51684 16838 51696 16890
rect 51748 16838 51760 16890
rect 51812 16838 58880 16890
rect 1104 16816 58880 16838
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 6362 16776 6368 16788
rect 4571 16748 6368 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 6362 16736 6368 16748
rect 6420 16736 6426 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 23477 16779 23535 16785
rect 6503 16748 9536 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 5721 16711 5779 16717
rect 5721 16677 5733 16711
rect 5767 16708 5779 16711
rect 6270 16708 6276 16720
rect 5767 16680 6276 16708
rect 5767 16677 5779 16680
rect 5721 16671 5779 16677
rect 6270 16668 6276 16680
rect 6328 16668 6334 16720
rect 5328 16643 5386 16649
rect 5328 16640 5340 16643
rect 4356 16612 5340 16640
rect 4356 16584 4384 16612
rect 5328 16609 5340 16612
rect 5374 16609 5386 16643
rect 5328 16603 5386 16609
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6365 16643 6423 16649
rect 6227 16612 6316 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 2188 16544 2237 16572
rect 2188 16532 2194 16544
rect 2225 16541 2237 16544
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2492 16575 2550 16581
rect 2492 16541 2504 16575
rect 2538 16572 2550 16575
rect 2958 16572 2964 16584
rect 2538 16544 2964 16572
rect 2538 16541 2550 16544
rect 2492 16535 2550 16541
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 4338 16532 4344 16584
rect 4396 16532 4402 16584
rect 5166 16532 5172 16584
rect 5224 16532 5230 16584
rect 5442 16532 5448 16584
rect 5500 16532 5506 16584
rect 6288 16572 6316 16612
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 6472 16640 6500 16739
rect 6411 16612 6500 16640
rect 8573 16643 8631 16649
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9398 16640 9404 16652
rect 8619 16612 9404 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9508 16649 9536 16748
rect 23477 16745 23489 16779
rect 23523 16776 23535 16779
rect 23750 16776 23756 16788
rect 23523 16748 23756 16776
rect 23523 16745 23535 16748
rect 23477 16739 23535 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 26602 16736 26608 16788
rect 26660 16736 26666 16788
rect 31665 16779 31723 16785
rect 31665 16745 31677 16779
rect 31711 16776 31723 16779
rect 31938 16776 31944 16788
rect 31711 16748 31944 16776
rect 31711 16745 31723 16748
rect 31665 16739 31723 16745
rect 31938 16736 31944 16748
rect 31996 16776 32002 16788
rect 32858 16776 32864 16788
rect 31996 16748 32864 16776
rect 31996 16736 32002 16748
rect 32858 16736 32864 16748
rect 32916 16776 32922 16788
rect 33781 16779 33839 16785
rect 33781 16776 33793 16779
rect 32916 16748 33793 16776
rect 32916 16736 32922 16748
rect 33781 16745 33793 16748
rect 33827 16776 33839 16779
rect 34514 16776 34520 16788
rect 33827 16748 34520 16776
rect 33827 16745 33839 16748
rect 33781 16739 33839 16745
rect 34514 16736 34520 16748
rect 34572 16736 34578 16788
rect 38286 16736 38292 16788
rect 38344 16776 38350 16788
rect 39117 16779 39175 16785
rect 39117 16776 39129 16779
rect 38344 16748 39129 16776
rect 38344 16736 38350 16748
rect 39117 16745 39129 16748
rect 39163 16776 39175 16779
rect 39850 16776 39856 16788
rect 39163 16748 39856 16776
rect 39163 16745 39175 16748
rect 39117 16739 39175 16745
rect 39850 16736 39856 16748
rect 39908 16736 39914 16788
rect 42426 16776 42432 16788
rect 42260 16748 42432 16776
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 12158 16708 12164 16720
rect 9732 16680 12164 16708
rect 9732 16668 9738 16680
rect 12158 16668 12164 16680
rect 12216 16708 12222 16720
rect 12894 16708 12900 16720
rect 12216 16680 12900 16708
rect 12216 16668 12222 16680
rect 12894 16668 12900 16680
rect 12952 16708 12958 16720
rect 13173 16711 13231 16717
rect 13173 16708 13185 16711
rect 12952 16680 13185 16708
rect 12952 16668 12958 16680
rect 13173 16677 13185 16680
rect 13219 16708 13231 16711
rect 17586 16708 17592 16720
rect 13219 16680 17592 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 17586 16668 17592 16680
rect 17644 16668 17650 16720
rect 23382 16668 23388 16720
rect 23440 16708 23446 16720
rect 26620 16708 26648 16736
rect 23440 16680 26648 16708
rect 32033 16711 32091 16717
rect 23440 16668 23446 16680
rect 32033 16677 32045 16711
rect 32079 16708 32091 16711
rect 32398 16708 32404 16720
rect 32079 16680 32404 16708
rect 32079 16677 32091 16680
rect 32033 16671 32091 16677
rect 32398 16668 32404 16680
rect 32456 16668 32462 16720
rect 41693 16711 41751 16717
rect 41693 16677 41705 16711
rect 41739 16677 41751 16711
rect 41693 16671 41751 16677
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 17678 16600 17684 16652
rect 17736 16600 17742 16652
rect 18782 16600 18788 16652
rect 18840 16600 18846 16652
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16640 23719 16643
rect 23707 16612 24348 16640
rect 23707 16609 23719 16612
rect 23661 16603 23719 16609
rect 24320 16584 24348 16612
rect 25590 16600 25596 16652
rect 25648 16640 25654 16652
rect 26234 16640 26240 16652
rect 25648 16612 26240 16640
rect 25648 16600 25654 16612
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 32416 16640 32444 16668
rect 32416 16612 33180 16640
rect 6288 16544 7236 16572
rect 4614 16504 4620 16516
rect 3620 16476 4620 16504
rect 3620 16445 3648 16476
rect 4614 16464 4620 16476
rect 4672 16464 4678 16516
rect 7208 16504 7236 16544
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7837 16575 7895 16581
rect 7837 16572 7849 16575
rect 7340 16544 7849 16572
rect 7340 16532 7346 16544
rect 7837 16541 7849 16544
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 7926 16532 7932 16584
rect 7984 16532 7990 16584
rect 8754 16572 8760 16584
rect 8036 16544 8760 16572
rect 7466 16504 7472 16516
rect 7208 16476 7472 16504
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 7592 16507 7650 16513
rect 7592 16473 7604 16507
rect 7638 16504 7650 16507
rect 7944 16504 7972 16532
rect 7638 16476 7972 16504
rect 7638 16473 7650 16476
rect 7592 16467 7650 16473
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16405 3663 16439
rect 3605 16399 3663 16405
rect 3786 16396 3792 16448
rect 3844 16396 3850 16448
rect 4632 16436 4660 16464
rect 5442 16436 5448 16448
rect 4632 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8036 16436 8064 16544
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 11514 16532 11520 16584
rect 11572 16532 11578 16584
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 13814 16532 13820 16584
rect 13872 16532 13878 16584
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13964 16544 14105 16572
rect 13964 16532 13970 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 15252 16544 15393 16572
rect 15252 16532 15258 16544
rect 15381 16541 15393 16544
rect 15427 16541 15439 16575
rect 15381 16535 15439 16541
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18104 16544 18337 16572
rect 18104 16532 18110 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 21358 16532 21364 16584
rect 21416 16532 21422 16584
rect 24302 16532 24308 16584
rect 24360 16532 24366 16584
rect 25038 16532 25044 16584
rect 25096 16532 25102 16584
rect 26326 16532 26332 16584
rect 26384 16532 26390 16584
rect 30834 16532 30840 16584
rect 30892 16532 30898 16584
rect 33152 16572 33180 16612
rect 35618 16600 35624 16652
rect 35676 16640 35682 16652
rect 35989 16643 36047 16649
rect 35989 16640 36001 16643
rect 35676 16612 36001 16640
rect 35676 16600 35682 16612
rect 35989 16609 36001 16612
rect 36035 16609 36047 16643
rect 35989 16603 36047 16609
rect 37826 16600 37832 16652
rect 37884 16640 37890 16652
rect 38470 16640 38476 16652
rect 37884 16612 38476 16640
rect 37884 16600 37890 16612
rect 38470 16600 38476 16612
rect 38528 16600 38534 16652
rect 33502 16572 33508 16584
rect 33152 16544 33508 16572
rect 33502 16532 33508 16544
rect 33560 16532 33566 16584
rect 35250 16532 35256 16584
rect 35308 16532 35314 16584
rect 36814 16532 36820 16584
rect 36872 16572 36878 16584
rect 37001 16575 37059 16581
rect 37001 16572 37013 16575
rect 36872 16544 37013 16572
rect 36872 16532 36878 16544
rect 37001 16541 37013 16544
rect 37047 16541 37059 16575
rect 37001 16535 37059 16541
rect 37918 16532 37924 16584
rect 37976 16532 37982 16584
rect 38838 16532 38844 16584
rect 38896 16572 38902 16584
rect 40129 16575 40187 16581
rect 40129 16572 40141 16575
rect 38896 16544 40141 16572
rect 38896 16532 38902 16544
rect 40129 16541 40141 16544
rect 40175 16572 40187 16575
rect 40313 16575 40371 16581
rect 40313 16572 40325 16575
rect 40175 16544 40325 16572
rect 40175 16541 40187 16544
rect 40129 16535 40187 16541
rect 40313 16541 40325 16544
rect 40359 16541 40371 16575
rect 41708 16572 41736 16671
rect 42260 16649 42288 16748
rect 42426 16736 42432 16748
rect 42484 16736 42490 16788
rect 44545 16779 44603 16785
rect 44545 16776 44557 16779
rect 42904 16748 44557 16776
rect 42245 16643 42303 16649
rect 42245 16609 42257 16643
rect 42291 16609 42303 16643
rect 42245 16603 42303 16609
rect 42334 16600 42340 16652
rect 42392 16600 42398 16652
rect 42904 16649 42932 16748
rect 44545 16745 44557 16748
rect 44591 16776 44603 16779
rect 45554 16776 45560 16788
rect 44591 16748 45560 16776
rect 44591 16745 44603 16748
rect 44545 16739 44603 16745
rect 45554 16736 45560 16748
rect 45612 16736 45618 16788
rect 49694 16736 49700 16788
rect 49752 16776 49758 16788
rect 51077 16779 51135 16785
rect 51077 16776 51089 16779
rect 49752 16748 51089 16776
rect 49752 16736 49758 16748
rect 51077 16745 51089 16748
rect 51123 16745 51135 16779
rect 51077 16739 51135 16745
rect 44266 16668 44272 16720
rect 44324 16708 44330 16720
rect 44634 16708 44640 16720
rect 44324 16680 44640 16708
rect 44324 16668 44330 16680
rect 44634 16668 44640 16680
rect 44692 16668 44698 16720
rect 50522 16708 50528 16720
rect 48792 16680 50528 16708
rect 48792 16652 48820 16680
rect 50522 16668 50528 16680
rect 50580 16668 50586 16720
rect 57333 16711 57391 16717
rect 57333 16677 57345 16711
rect 57379 16708 57391 16711
rect 57379 16680 58020 16708
rect 57379 16677 57391 16680
rect 57333 16671 57391 16677
rect 42889 16643 42947 16649
rect 42889 16609 42901 16643
rect 42935 16609 42947 16643
rect 42889 16603 42947 16609
rect 45094 16600 45100 16652
rect 45152 16640 45158 16652
rect 45557 16643 45615 16649
rect 45557 16640 45569 16643
rect 45152 16612 45569 16640
rect 45152 16600 45158 16612
rect 45557 16609 45569 16612
rect 45603 16640 45615 16643
rect 48774 16640 48780 16652
rect 45603 16612 48780 16640
rect 45603 16609 45615 16612
rect 45557 16603 45615 16609
rect 48774 16600 48780 16612
rect 48832 16600 48838 16652
rect 49418 16600 49424 16652
rect 49476 16640 49482 16652
rect 54570 16640 54576 16652
rect 49476 16612 54576 16640
rect 49476 16600 49482 16612
rect 54570 16600 54576 16612
rect 54628 16600 54634 16652
rect 56505 16643 56563 16649
rect 56505 16609 56517 16643
rect 56551 16640 56563 16643
rect 56781 16643 56839 16649
rect 56781 16640 56793 16643
rect 56551 16612 56793 16640
rect 56551 16609 56563 16612
rect 56505 16603 56563 16609
rect 56781 16609 56793 16612
rect 56827 16640 56839 16643
rect 57054 16640 57060 16652
rect 56827 16612 57060 16640
rect 56827 16609 56839 16612
rect 56781 16603 56839 16609
rect 57054 16600 57060 16612
rect 57112 16600 57118 16652
rect 57992 16649 58020 16680
rect 57977 16643 58035 16649
rect 57977 16609 57989 16643
rect 58023 16609 58035 16643
rect 57977 16603 58035 16609
rect 42978 16572 42984 16584
rect 41708 16544 42984 16572
rect 40313 16535 40371 16541
rect 42978 16532 42984 16544
rect 43036 16532 43042 16584
rect 43156 16575 43214 16581
rect 43156 16541 43168 16575
rect 43202 16572 43214 16575
rect 43990 16572 43996 16584
rect 43202 16544 43996 16572
rect 43202 16541 43214 16544
rect 43156 16535 43214 16541
rect 43990 16532 43996 16544
rect 44048 16532 44054 16584
rect 44818 16532 44824 16584
rect 44876 16572 44882 16584
rect 45373 16575 45431 16581
rect 45373 16572 45385 16575
rect 44876 16544 45385 16572
rect 44876 16532 44882 16544
rect 45373 16541 45385 16544
rect 45419 16541 45431 16575
rect 45373 16535 45431 16541
rect 45646 16532 45652 16584
rect 45704 16532 45710 16584
rect 47762 16532 47768 16584
rect 47820 16532 47826 16584
rect 49142 16532 49148 16584
rect 49200 16532 49206 16584
rect 49970 16532 49976 16584
rect 50028 16572 50034 16584
rect 50709 16575 50767 16581
rect 50709 16572 50721 16575
rect 50028 16544 50721 16572
rect 50028 16532 50034 16544
rect 50709 16541 50721 16544
rect 50755 16541 50767 16575
rect 50709 16535 50767 16541
rect 53834 16532 53840 16584
rect 53892 16532 53898 16584
rect 56965 16575 57023 16581
rect 56965 16541 56977 16575
rect 57011 16572 57023 16575
rect 57882 16572 57888 16584
rect 57011 16544 57888 16572
rect 57011 16541 57023 16544
rect 56965 16535 57023 16541
rect 57882 16532 57888 16544
rect 57940 16532 57946 16584
rect 34238 16464 34244 16516
rect 34296 16504 34302 16516
rect 40580 16507 40638 16513
rect 34296 16476 40264 16504
rect 34296 16464 34302 16476
rect 7975 16408 8064 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 8168 16408 8309 16436
rect 8168 16396 8174 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 8297 16399 8355 16405
rect 8389 16439 8447 16445
rect 8389 16405 8401 16439
rect 8435 16436 8447 16439
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8435 16408 8953 16436
rect 8435 16405 8447 16408
rect 8389 16399 8447 16405
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 10870 16396 10876 16448
rect 10928 16396 10934 16448
rect 11698 16396 11704 16448
rect 11756 16396 11762 16448
rect 12710 16396 12716 16448
rect 12768 16396 12774 16448
rect 13262 16396 13268 16448
rect 13320 16396 13326 16448
rect 14734 16396 14740 16448
rect 14792 16396 14798 16448
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17037 16439 17095 16445
rect 17037 16436 17049 16439
rect 16908 16408 17049 16436
rect 16908 16396 16914 16408
rect 17037 16405 17049 16408
rect 17083 16405 17095 16439
rect 17037 16399 17095 16405
rect 17770 16396 17776 16448
rect 17828 16396 17834 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20809 16439 20867 16445
rect 20809 16436 20821 16439
rect 20772 16408 20821 16436
rect 20772 16396 20778 16408
rect 20809 16405 20821 16408
rect 20855 16405 20867 16439
rect 20809 16399 20867 16405
rect 24210 16396 24216 16448
rect 24268 16396 24274 16448
rect 24394 16396 24400 16448
rect 24452 16396 24458 16448
rect 25590 16396 25596 16448
rect 25648 16436 25654 16448
rect 25777 16439 25835 16445
rect 25777 16436 25789 16439
rect 25648 16408 25789 16436
rect 25648 16396 25654 16408
rect 25777 16405 25789 16408
rect 25823 16405 25835 16439
rect 25777 16399 25835 16405
rect 30282 16396 30288 16448
rect 30340 16396 30346 16448
rect 31202 16396 31208 16448
rect 31260 16396 31266 16448
rect 34698 16396 34704 16448
rect 34756 16396 34762 16448
rect 35434 16396 35440 16448
rect 35492 16396 35498 16448
rect 36446 16396 36452 16448
rect 36504 16396 36510 16448
rect 36906 16396 36912 16448
rect 36964 16436 36970 16448
rect 37185 16439 37243 16445
rect 37185 16436 37197 16439
rect 36964 16408 37197 16436
rect 36964 16396 36970 16408
rect 37185 16405 37197 16408
rect 37231 16405 37243 16439
rect 37185 16399 37243 16405
rect 38562 16396 38568 16448
rect 38620 16396 38626 16448
rect 40236 16436 40264 16476
rect 40580 16473 40592 16507
rect 40626 16504 40638 16507
rect 41230 16504 41236 16516
rect 40626 16476 41236 16504
rect 40626 16473 40638 16476
rect 40580 16467 40638 16473
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 42996 16504 43024 16532
rect 43346 16504 43352 16516
rect 41386 16476 42840 16504
rect 42996 16476 43352 16504
rect 41386 16436 41414 16476
rect 40236 16408 41414 16436
rect 41782 16396 41788 16448
rect 41840 16396 41846 16448
rect 42153 16439 42211 16445
rect 42153 16405 42165 16439
rect 42199 16436 42211 16439
rect 42242 16436 42248 16448
rect 42199 16408 42248 16436
rect 42199 16405 42211 16408
rect 42153 16399 42211 16405
rect 42242 16396 42248 16408
rect 42300 16396 42306 16448
rect 42812 16436 42840 16476
rect 43346 16464 43352 16476
rect 43404 16464 43410 16516
rect 45664 16504 45692 16532
rect 45020 16476 45692 16504
rect 44174 16436 44180 16448
rect 42812 16408 44180 16436
rect 44174 16396 44180 16408
rect 44232 16396 44238 16448
rect 45020 16445 45048 16476
rect 45738 16464 45744 16516
rect 45796 16504 45802 16516
rect 55766 16504 55772 16516
rect 45796 16476 55772 16504
rect 45796 16464 45802 16476
rect 55766 16464 55772 16476
rect 55824 16464 55830 16516
rect 45005 16439 45063 16445
rect 45005 16405 45017 16439
rect 45051 16405 45063 16439
rect 45005 16399 45063 16405
rect 45370 16396 45376 16448
rect 45428 16436 45434 16448
rect 45465 16439 45523 16445
rect 45465 16436 45477 16439
rect 45428 16408 45477 16436
rect 45428 16396 45434 16408
rect 45465 16405 45477 16408
rect 45511 16405 45523 16439
rect 45465 16399 45523 16405
rect 48222 16396 48228 16448
rect 48280 16436 48286 16448
rect 48409 16439 48467 16445
rect 48409 16436 48421 16439
rect 48280 16408 48421 16436
rect 48280 16396 48286 16408
rect 48409 16405 48421 16408
rect 48455 16405 48467 16439
rect 48409 16399 48467 16405
rect 48590 16396 48596 16448
rect 48648 16396 48654 16448
rect 50154 16396 50160 16448
rect 50212 16396 50218 16448
rect 53098 16396 53104 16448
rect 53156 16436 53162 16448
rect 53193 16439 53251 16445
rect 53193 16436 53205 16439
rect 53156 16408 53205 16436
rect 53156 16396 53162 16408
rect 53193 16405 53205 16408
rect 53239 16405 53251 16439
rect 53193 16399 53251 16405
rect 56778 16396 56784 16448
rect 56836 16436 56842 16448
rect 56873 16439 56931 16445
rect 56873 16436 56885 16439
rect 56836 16408 56885 16436
rect 56836 16396 56842 16408
rect 56873 16405 56885 16408
rect 56919 16405 56931 16439
rect 56873 16399 56931 16405
rect 57422 16396 57428 16448
rect 57480 16396 57486 16448
rect 1104 16346 59040 16368
rect 1104 16294 15394 16346
rect 15446 16294 15458 16346
rect 15510 16294 15522 16346
rect 15574 16294 15586 16346
rect 15638 16294 15650 16346
rect 15702 16294 29838 16346
rect 29890 16294 29902 16346
rect 29954 16294 29966 16346
rect 30018 16294 30030 16346
rect 30082 16294 30094 16346
rect 30146 16294 44282 16346
rect 44334 16294 44346 16346
rect 44398 16294 44410 16346
rect 44462 16294 44474 16346
rect 44526 16294 44538 16346
rect 44590 16294 58726 16346
rect 58778 16294 58790 16346
rect 58842 16294 58854 16346
rect 58906 16294 58918 16346
rect 58970 16294 58982 16346
rect 59034 16294 59040 16346
rect 1104 16272 59040 16294
rect 3234 16192 3240 16244
rect 3292 16232 3298 16244
rect 3513 16235 3571 16241
rect 3513 16232 3525 16235
rect 3292 16204 3525 16232
rect 3292 16192 3298 16204
rect 3513 16201 3525 16204
rect 3559 16201 3571 16235
rect 3513 16195 3571 16201
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3844 16204 3893 16232
rect 3844 16192 3850 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 3970 16192 3976 16244
rect 4028 16192 4034 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6270 16232 6276 16244
rect 6227 16204 6276 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 2308 16167 2366 16173
rect 2308 16133 2320 16167
rect 2354 16164 2366 16167
rect 2590 16164 2596 16176
rect 2354 16136 2596 16164
rect 2354 16133 2366 16136
rect 2308 16127 2366 16133
rect 2590 16124 2596 16136
rect 2648 16124 2654 16176
rect 7300 16164 7328 16195
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 7524 16204 8769 16232
rect 7524 16192 7530 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 7622 16167 7680 16173
rect 7622 16164 7634 16167
rect 7300 16136 7634 16164
rect 7622 16133 7634 16136
rect 7668 16133 7680 16167
rect 7622 16127 7680 16133
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7340 16068 7389 16096
rect 7340 16056 7346 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 8772 16096 8800 16195
rect 11514 16192 11520 16244
rect 11572 16192 11578 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11756 16204 11897 16232
rect 11756 16192 11762 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 13173 16235 13231 16241
rect 13173 16201 13185 16235
rect 13219 16232 13231 16235
rect 13262 16232 13268 16244
rect 13219 16204 13268 16232
rect 13219 16201 13231 16204
rect 13173 16195 13231 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13633 16235 13691 16241
rect 13633 16201 13645 16235
rect 13679 16232 13691 16235
rect 13906 16232 13912 16244
rect 13679 16204 13912 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16232 14151 16235
rect 14826 16232 14832 16244
rect 14139 16204 14832 16232
rect 14139 16201 14151 16204
rect 14093 16195 14151 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 17770 16192 17776 16244
rect 17828 16192 17834 16244
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20622 16232 20628 16244
rect 19760 16204 20628 16232
rect 19760 16192 19766 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 24029 16235 24087 16241
rect 24029 16201 24041 16235
rect 24075 16232 24087 16235
rect 24210 16232 24216 16244
rect 24075 16204 24216 16232
rect 24075 16201 24087 16204
rect 24029 16195 24087 16201
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 24854 16192 24860 16244
rect 24912 16192 24918 16244
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 26326 16232 26332 16244
rect 25915 16204 26332 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 30469 16235 30527 16241
rect 30469 16201 30481 16235
rect 30515 16232 30527 16235
rect 30834 16232 30840 16244
rect 30515 16204 30840 16232
rect 30515 16201 30527 16204
rect 30469 16195 30527 16201
rect 30834 16192 30840 16204
rect 30892 16192 30898 16244
rect 33965 16235 34023 16241
rect 33965 16201 33977 16235
rect 34011 16232 34023 16235
rect 34514 16232 34520 16244
rect 34011 16204 34520 16232
rect 34011 16201 34023 16204
rect 33965 16195 34023 16201
rect 34514 16192 34520 16204
rect 34572 16232 34578 16244
rect 35250 16232 35256 16244
rect 34572 16204 35256 16232
rect 34572 16192 34578 16204
rect 35250 16192 35256 16204
rect 35308 16192 35314 16244
rect 35434 16192 35440 16244
rect 35492 16192 35498 16244
rect 36446 16192 36452 16244
rect 36504 16192 36510 16244
rect 37093 16235 37151 16241
rect 37093 16201 37105 16235
rect 37139 16232 37151 16235
rect 37826 16232 37832 16244
rect 37139 16204 37832 16232
rect 37139 16201 37151 16204
rect 37093 16195 37151 16201
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 38562 16192 38568 16244
rect 38620 16192 38626 16244
rect 41230 16192 41236 16244
rect 41288 16192 41294 16244
rect 41782 16192 41788 16244
rect 41840 16192 41846 16244
rect 42429 16235 42487 16241
rect 42429 16201 42441 16235
rect 42475 16232 42487 16235
rect 43622 16232 43628 16244
rect 42475 16204 43628 16232
rect 42475 16201 42487 16204
rect 42429 16195 42487 16201
rect 43622 16192 43628 16204
rect 43680 16192 43686 16244
rect 47581 16235 47639 16241
rect 47581 16201 47593 16235
rect 47627 16232 47639 16235
rect 47762 16232 47768 16244
rect 47627 16204 47768 16232
rect 47627 16201 47639 16204
rect 47581 16195 47639 16201
rect 47762 16192 47768 16204
rect 47820 16192 47826 16244
rect 48041 16235 48099 16241
rect 48041 16201 48053 16235
rect 48087 16232 48099 16235
rect 48590 16232 48596 16244
rect 48087 16204 48596 16232
rect 48087 16201 48099 16204
rect 48041 16195 48099 16201
rect 48590 16192 48596 16204
rect 48648 16192 48654 16244
rect 51721 16235 51779 16241
rect 51721 16232 51733 16235
rect 49252 16204 51733 16232
rect 16936 16167 16994 16173
rect 16936 16133 16948 16167
rect 16982 16164 16994 16167
rect 17788 16164 17816 16192
rect 16982 16136 17816 16164
rect 20824 16164 20852 16192
rect 33873 16167 33931 16173
rect 20824 16136 21220 16164
rect 16982 16133 16994 16136
rect 16936 16127 16994 16133
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 8772 16068 9413 16096
rect 7377 16059 7435 16065
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 11606 16096 11612 16108
rect 10836 16068 11612 16096
rect 10836 16056 10842 16068
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 11882 16056 11888 16108
rect 11940 16096 11946 16108
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11940 16068 11989 16096
rect 11940 16056 11946 16068
rect 11977 16065 11989 16068
rect 12023 16096 12035 16099
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 12023 16068 13277 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 13265 16065 13277 16068
rect 13311 16096 13323 16099
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13311 16068 14013 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16096 19395 16099
rect 19886 16096 19892 16108
rect 19383 16068 19892 16096
rect 19383 16065 19395 16068
rect 19337 16059 19395 16065
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 20921 16099 20979 16105
rect 20921 16065 20933 16099
rect 20967 16096 20979 16099
rect 21082 16096 21088 16108
rect 20967 16068 21088 16096
rect 20967 16065 20979 16068
rect 20921 16059 20979 16065
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 21192 16105 21220 16136
rect 33873 16133 33885 16167
rect 33919 16164 33931 16167
rect 34238 16164 34244 16176
rect 33919 16136 34244 16164
rect 33919 16133 33931 16136
rect 33873 16127 33931 16133
rect 34238 16124 34244 16136
rect 34296 16124 34302 16176
rect 35100 16167 35158 16173
rect 35100 16133 35112 16167
rect 35146 16164 35158 16167
rect 35452 16164 35480 16192
rect 35146 16136 35480 16164
rect 35980 16167 36038 16173
rect 35146 16133 35158 16136
rect 35100 16127 35158 16133
rect 35980 16133 35992 16167
rect 36026 16164 36038 16167
rect 36464 16164 36492 16192
rect 36026 16136 36492 16164
rect 38412 16167 38470 16173
rect 36026 16133 36038 16136
rect 35980 16127 36038 16133
rect 38412 16133 38424 16167
rect 38458 16164 38470 16167
rect 38580 16164 38608 16192
rect 38458 16136 38608 16164
rect 38458 16133 38470 16136
rect 38412 16127 38470 16133
rect 21177 16099 21235 16105
rect 21177 16065 21189 16099
rect 21223 16065 21235 16099
rect 23937 16099 23995 16105
rect 21177 16059 21235 16065
rect 22066 16068 23796 16096
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 4203 16000 4660 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 4338 15960 4344 15972
rect 3467 15932 4344 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 4338 15920 4344 15932
rect 4396 15920 4402 15972
rect 4632 15901 4660 16000
rect 6730 15988 6736 16040
rect 6788 15988 6794 16040
rect 10796 15960 10824 16056
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 11790 15988 11796 16040
rect 11848 15988 11854 16040
rect 12158 15988 12164 16040
rect 12216 15988 12222 16040
rect 12710 16028 12716 16040
rect 12406 16000 12716 16028
rect 8680 15932 10824 15960
rect 11808 15960 11836 15988
rect 12406 15960 12434 16000
rect 12710 15988 12716 16000
rect 12768 16028 12774 16040
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12768 16000 13001 16028
rect 12768 15988 12774 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14642 16028 14648 16040
rect 13955 16000 14648 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 11808 15932 12434 15960
rect 12805 15963 12863 15969
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 8680 15892 8708 15932
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13924 15960 13952 15991
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 12851 15932 13952 15960
rect 14461 15963 14519 15969
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 14461 15929 14473 15963
rect 14507 15960 14519 15963
rect 14936 15960 14964 15991
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16540 16000 16681 16028
rect 16540 15988 16546 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 20162 16028 20168 16040
rect 19015 16000 20168 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 14507 15932 14964 15960
rect 18049 15963 18107 15969
rect 14507 15929 14519 15932
rect 14461 15923 14519 15929
rect 18049 15929 18061 15963
rect 18095 15960 18107 15963
rect 18984 15960 19012 15991
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 22066 15972 22094 16068
rect 23768 16040 23796 16068
rect 23937 16065 23949 16099
rect 23983 16096 23995 16099
rect 24670 16096 24676 16108
rect 23983 16068 24676 16096
rect 23983 16065 23995 16068
rect 23937 16059 23995 16065
rect 24670 16056 24676 16068
rect 24728 16096 24734 16108
rect 25774 16096 25780 16108
rect 24728 16068 25780 16096
rect 24728 16056 24734 16068
rect 25774 16056 25780 16068
rect 25832 16096 25838 16108
rect 26237 16099 26295 16105
rect 26237 16096 26249 16099
rect 25832 16068 26249 16096
rect 25832 16056 25838 16068
rect 26237 16065 26249 16068
rect 26283 16065 26295 16099
rect 26237 16059 26295 16065
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16096 26387 16099
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26375 16068 26985 16096
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 30834 16056 30840 16108
rect 30892 16056 30898 16108
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16096 30987 16099
rect 31297 16099 31355 16105
rect 31297 16096 31309 16099
rect 30975 16068 31309 16096
rect 30975 16065 30987 16068
rect 30929 16059 30987 16065
rect 31297 16065 31309 16068
rect 31343 16065 31355 16099
rect 31297 16059 31355 16065
rect 35342 16056 35348 16108
rect 35400 16096 35406 16108
rect 35713 16099 35771 16105
rect 35713 16096 35725 16099
rect 35400 16068 35725 16096
rect 35400 16056 35406 16068
rect 35713 16065 35725 16068
rect 35759 16065 35771 16099
rect 35713 16059 35771 16065
rect 38657 16099 38715 16105
rect 38657 16065 38669 16099
rect 38703 16096 38715 16099
rect 38838 16096 38844 16108
rect 38703 16068 38844 16096
rect 38703 16065 38715 16068
rect 38657 16059 38715 16065
rect 38838 16056 38844 16068
rect 38896 16056 38902 16108
rect 41800 16105 41828 16192
rect 41785 16099 41843 16105
rect 41785 16065 41797 16099
rect 41831 16065 41843 16099
rect 41785 16059 41843 16065
rect 43346 16056 43352 16108
rect 43404 16056 43410 16108
rect 44085 16099 44143 16105
rect 44085 16065 44097 16099
rect 44131 16096 44143 16099
rect 44634 16096 44640 16108
rect 44131 16068 44640 16096
rect 44131 16065 44143 16068
rect 44085 16059 44143 16065
rect 44634 16056 44640 16068
rect 44692 16056 44698 16108
rect 47578 16096 47584 16108
rect 45020 16068 47584 16096
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 18095 15932 19012 15960
rect 18095 15929 18107 15932
rect 18049 15923 18107 15929
rect 19058 15920 19064 15972
rect 19116 15960 19122 15972
rect 22002 15960 22008 15972
rect 19116 15932 19932 15960
rect 19116 15920 19122 15932
rect 4663 15864 8708 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 8846 15852 8852 15904
rect 8904 15852 8910 15904
rect 10686 15852 10692 15904
rect 10744 15852 10750 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 12894 15892 12900 15904
rect 11572 15864 12900 15892
rect 11572 15852 11578 15864
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 15562 15852 15568 15904
rect 15620 15852 15626 15904
rect 18322 15852 18328 15904
rect 18380 15852 18386 15904
rect 19794 15852 19800 15904
rect 19852 15852 19858 15904
rect 19904 15892 19932 15932
rect 21192 15932 22008 15960
rect 21192 15892 21220 15932
rect 22002 15920 22008 15932
rect 22060 15932 22094 15972
rect 22940 15960 22968 15991
rect 23750 15988 23756 16040
rect 23808 16028 23814 16040
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 23808 16000 24133 16028
rect 23808 15988 23814 16000
rect 24121 15997 24133 16000
rect 24167 15997 24179 16031
rect 24121 15991 24179 15997
rect 25498 15988 25504 16040
rect 25556 15988 25562 16040
rect 26513 16031 26571 16037
rect 26513 15997 26525 16031
rect 26559 16028 26571 16031
rect 26602 16028 26608 16040
rect 26559 16000 26608 16028
rect 26559 15997 26571 16000
rect 26513 15991 26571 15997
rect 26602 15988 26608 16000
rect 26660 15988 26666 16040
rect 27522 15988 27528 16040
rect 27580 15988 27586 16040
rect 28350 15988 28356 16040
rect 28408 15988 28414 16040
rect 30377 16031 30435 16037
rect 30377 15997 30389 16031
rect 30423 16028 30435 16031
rect 31018 16028 31024 16040
rect 30423 16000 31024 16028
rect 30423 15997 30435 16000
rect 30377 15991 30435 15997
rect 31018 15988 31024 16000
rect 31076 15988 31082 16040
rect 31846 15988 31852 16040
rect 31904 15988 31910 16040
rect 39301 16031 39359 16037
rect 39301 15997 39313 16031
rect 39347 15997 39359 16031
rect 39301 15991 39359 15997
rect 23569 15963 23627 15969
rect 23569 15960 23581 15963
rect 22940 15932 23581 15960
rect 22060 15920 22066 15932
rect 23569 15929 23581 15932
rect 23615 15929 23627 15963
rect 23569 15923 23627 15929
rect 24302 15920 24308 15972
rect 24360 15960 24366 15972
rect 39316 15960 39344 15991
rect 41322 15988 41328 16040
rect 41380 16028 41386 16040
rect 42886 16028 42892 16040
rect 41380 16000 42892 16028
rect 41380 15988 41386 16000
rect 42886 15988 42892 16000
rect 42944 16028 42950 16040
rect 43070 16028 43076 16040
rect 42944 16000 43076 16028
rect 42944 15988 42950 16000
rect 43070 15988 43076 16000
rect 43128 15988 43134 16040
rect 43254 16037 43260 16040
rect 43232 16031 43260 16037
rect 43232 15997 43244 16031
rect 43232 15991 43260 15997
rect 43254 15988 43260 15991
rect 43312 15988 43318 16040
rect 43530 15988 43536 16040
rect 43588 16028 43594 16040
rect 43625 16031 43683 16037
rect 43625 16028 43637 16031
rect 43588 16000 43637 16028
rect 43588 15988 43594 16000
rect 43625 15997 43637 16000
rect 43671 15997 43683 16031
rect 43625 15991 43683 15997
rect 44269 16031 44327 16037
rect 44269 15997 44281 16031
rect 44315 16028 44327 16031
rect 44726 16028 44732 16040
rect 44315 16000 44732 16028
rect 44315 15997 44327 16000
rect 44269 15991 44327 15997
rect 44726 15988 44732 16000
rect 44784 16028 44790 16040
rect 44913 16031 44971 16037
rect 44913 16028 44925 16031
rect 44784 16000 44925 16028
rect 44784 15988 44790 16000
rect 44913 15997 44925 16000
rect 44959 15997 44971 16031
rect 44913 15991 44971 15997
rect 24360 15932 26648 15960
rect 24360 15920 24366 15932
rect 26620 15904 26648 15932
rect 38672 15932 39344 15960
rect 42153 15963 42211 15969
rect 19904 15864 21220 15892
rect 21545 15895 21603 15901
rect 21545 15861 21557 15895
rect 21591 15892 21603 15895
rect 22094 15892 22100 15904
rect 21591 15864 22100 15892
rect 21591 15861 21603 15864
rect 21545 15855 21603 15861
rect 22094 15852 22100 15864
rect 22152 15892 22158 15904
rect 23382 15892 23388 15904
rect 22152 15864 23388 15892
rect 22152 15852 22158 15864
rect 23382 15852 23388 15864
rect 23440 15852 23446 15904
rect 23474 15852 23480 15904
rect 23532 15852 23538 15904
rect 24946 15852 24952 15904
rect 25004 15852 25010 15904
rect 26602 15852 26608 15904
rect 26660 15852 26666 15904
rect 27798 15852 27804 15904
rect 27856 15852 27862 15904
rect 32585 15895 32643 15901
rect 32585 15861 32597 15895
rect 32631 15892 32643 15895
rect 32858 15892 32864 15904
rect 32631 15864 32864 15892
rect 32631 15861 32643 15864
rect 32585 15855 32643 15861
rect 32858 15852 32864 15864
rect 32916 15852 32922 15904
rect 37277 15895 37335 15901
rect 37277 15861 37289 15895
rect 37323 15892 37335 15895
rect 37642 15892 37648 15904
rect 37323 15864 37648 15892
rect 37323 15861 37335 15864
rect 37277 15855 37335 15861
rect 37642 15852 37648 15864
rect 37700 15892 37706 15904
rect 38672 15892 38700 15932
rect 42153 15929 42165 15963
rect 42199 15960 42211 15963
rect 42610 15960 42616 15972
rect 42199 15932 42616 15960
rect 42199 15929 42211 15932
rect 42153 15923 42211 15929
rect 42610 15920 42616 15932
rect 42668 15920 42674 15972
rect 45020 15960 45048 16068
rect 47578 16056 47584 16068
rect 47636 16056 47642 16108
rect 47949 16099 48007 16105
rect 47949 16065 47961 16099
rect 47995 16096 48007 16099
rect 48038 16096 48044 16108
rect 47995 16068 48044 16096
rect 47995 16065 48007 16068
rect 47949 16059 48007 16065
rect 48038 16056 48044 16068
rect 48096 16056 48102 16108
rect 49252 16105 49280 16204
rect 51721 16201 51733 16204
rect 51767 16232 51779 16235
rect 51994 16232 52000 16244
rect 51767 16204 52000 16232
rect 51767 16201 51779 16204
rect 51721 16195 51779 16201
rect 51994 16192 52000 16204
rect 52052 16232 52058 16244
rect 53009 16235 53067 16241
rect 53009 16232 53021 16235
rect 52052 16204 53021 16232
rect 52052 16192 52058 16204
rect 53009 16201 53021 16204
rect 53055 16232 53067 16235
rect 53190 16232 53196 16244
rect 53055 16204 53196 16232
rect 53055 16201 53067 16204
rect 53009 16195 53067 16201
rect 53190 16192 53196 16204
rect 53248 16192 53254 16244
rect 53285 16235 53343 16241
rect 53285 16201 53297 16235
rect 53331 16232 53343 16235
rect 53834 16232 53840 16244
rect 53331 16204 53840 16232
rect 53331 16201 53343 16204
rect 53285 16195 53343 16201
rect 53834 16192 53840 16204
rect 53892 16192 53898 16244
rect 55766 16192 55772 16244
rect 55824 16192 55830 16244
rect 57422 16192 57428 16244
rect 57480 16192 57486 16244
rect 57698 16192 57704 16244
rect 57756 16192 57762 16244
rect 49504 16167 49562 16173
rect 49504 16133 49516 16167
rect 49550 16164 49562 16167
rect 50154 16164 50160 16176
rect 49550 16136 50160 16164
rect 49550 16133 49562 16136
rect 49504 16127 49562 16133
rect 50154 16124 50160 16136
rect 50212 16124 50218 16176
rect 56588 16167 56646 16173
rect 56588 16133 56600 16167
rect 56634 16164 56646 16167
rect 57440 16164 57468 16192
rect 56634 16136 57468 16164
rect 56634 16133 56646 16136
rect 56588 16127 56646 16133
rect 49237 16099 49295 16105
rect 49237 16096 49249 16099
rect 48286 16068 49249 16096
rect 47118 15988 47124 16040
rect 47176 16028 47182 16040
rect 48133 16031 48191 16037
rect 48133 16028 48145 16031
rect 47176 16000 48145 16028
rect 47176 15988 47182 16000
rect 48133 15997 48145 16000
rect 48179 15997 48191 16031
rect 48133 15991 48191 15997
rect 47305 15963 47363 15969
rect 47305 15960 47317 15963
rect 43640 15932 45048 15960
rect 46860 15932 47317 15960
rect 37700 15864 38700 15892
rect 37700 15852 37706 15864
rect 38746 15852 38752 15904
rect 38804 15852 38810 15904
rect 41046 15852 41052 15904
rect 41104 15852 41110 15904
rect 42058 15852 42064 15904
rect 42116 15892 42122 15904
rect 43530 15892 43536 15904
rect 42116 15864 43536 15892
rect 42116 15852 42122 15864
rect 43530 15852 43536 15864
rect 43588 15892 43594 15904
rect 43640 15892 43668 15932
rect 46860 15904 46888 15932
rect 47305 15929 47317 15932
rect 47351 15960 47363 15963
rect 48286 15960 48314 16068
rect 49237 16065 49249 16068
rect 49283 16065 49295 16099
rect 49237 16059 49295 16065
rect 53653 16099 53711 16105
rect 53653 16065 53665 16099
rect 53699 16096 53711 16099
rect 54849 16099 54907 16105
rect 54849 16096 54861 16099
rect 53699 16068 54861 16096
rect 53699 16065 53711 16068
rect 53653 16059 53711 16065
rect 54849 16065 54861 16068
rect 54895 16065 54907 16099
rect 54849 16059 54907 16065
rect 57146 16056 57152 16108
rect 57204 16096 57210 16108
rect 58437 16099 58495 16105
rect 58437 16096 58449 16099
rect 57204 16068 58449 16096
rect 57204 16056 57210 16068
rect 58437 16065 58449 16068
rect 58483 16065 58495 16099
rect 58437 16059 58495 16065
rect 49050 15988 49056 16040
rect 49108 15988 49114 16040
rect 51261 16031 51319 16037
rect 51261 16028 51273 16031
rect 50632 16000 51273 16028
rect 47351 15932 48314 15960
rect 47351 15929 47363 15932
rect 47305 15923 47363 15929
rect 50632 15904 50660 16000
rect 51261 15997 51273 16000
rect 51307 15997 51319 16031
rect 51261 15991 51319 15997
rect 53742 15988 53748 16040
rect 53800 15988 53806 16040
rect 53837 16031 53895 16037
rect 53837 15997 53849 16031
rect 53883 15997 53895 16031
rect 53837 15991 53895 15997
rect 53852 15960 53880 15991
rect 54662 15988 54668 16040
rect 54720 15988 54726 16040
rect 55401 16031 55459 16037
rect 55401 15997 55413 16031
rect 55447 15997 55459 16031
rect 56321 16031 56379 16037
rect 56321 16028 56333 16031
rect 55401 15991 55459 15997
rect 56152 16000 56333 16028
rect 55416 15960 55444 15991
rect 56042 15960 56048 15972
rect 52564 15932 53880 15960
rect 54220 15932 56048 15960
rect 52564 15904 52592 15932
rect 54220 15904 54248 15932
rect 56042 15920 56048 15932
rect 56100 15920 56106 15972
rect 56152 15904 56180 16000
rect 56321 15997 56333 16000
rect 56367 15997 56379 16031
rect 56321 15991 56379 15997
rect 43588 15864 43668 15892
rect 43588 15852 43594 15864
rect 44358 15852 44364 15904
rect 44416 15852 44422 15904
rect 45094 15852 45100 15904
rect 45152 15892 45158 15904
rect 45281 15895 45339 15901
rect 45281 15892 45293 15895
rect 45152 15864 45293 15892
rect 45152 15852 45158 15864
rect 45281 15861 45293 15864
rect 45327 15861 45339 15895
rect 45281 15855 45339 15861
rect 46842 15852 46848 15904
rect 46900 15852 46906 15904
rect 47029 15895 47087 15901
rect 47029 15861 47041 15895
rect 47075 15892 47087 15895
rect 47118 15892 47124 15904
rect 47075 15864 47124 15892
rect 47075 15861 47087 15864
rect 47029 15855 47087 15861
rect 47118 15852 47124 15864
rect 47176 15852 47182 15904
rect 48406 15852 48412 15904
rect 48464 15852 48470 15904
rect 49050 15852 49056 15904
rect 49108 15892 49114 15904
rect 49510 15892 49516 15904
rect 49108 15864 49516 15892
rect 49108 15852 49114 15864
rect 49510 15852 49516 15864
rect 49568 15852 49574 15904
rect 50614 15852 50620 15904
rect 50672 15852 50678 15904
rect 50706 15852 50712 15904
rect 50764 15852 50770 15904
rect 52546 15852 52552 15904
rect 52604 15852 52610 15904
rect 54110 15852 54116 15904
rect 54168 15852 54174 15904
rect 54202 15852 54208 15904
rect 54260 15852 54266 15904
rect 56134 15852 56140 15904
rect 56192 15852 56198 15904
rect 57882 15852 57888 15904
rect 57940 15852 57946 15904
rect 1104 15802 58880 15824
rect 1104 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 22616 15802
rect 22668 15750 22680 15802
rect 22732 15750 22744 15802
rect 22796 15750 22808 15802
rect 22860 15750 22872 15802
rect 22924 15750 37060 15802
rect 37112 15750 37124 15802
rect 37176 15750 37188 15802
rect 37240 15750 37252 15802
rect 37304 15750 37316 15802
rect 37368 15750 51504 15802
rect 51556 15750 51568 15802
rect 51620 15750 51632 15802
rect 51684 15750 51696 15802
rect 51748 15750 51760 15802
rect 51812 15750 58880 15802
rect 1104 15728 58880 15750
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 6788 15660 7757 15688
rect 6788 15648 6794 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 8938 15688 8944 15700
rect 7745 15651 7803 15657
rect 8404 15660 8944 15688
rect 8404 15561 8432 15660
rect 8938 15648 8944 15660
rect 8996 15688 9002 15700
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 8996 15660 9229 15688
rect 8996 15648 9002 15660
rect 9217 15657 9229 15660
rect 9263 15688 9275 15691
rect 9858 15688 9864 15700
rect 9263 15660 9864 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 11514 15648 11520 15700
rect 11572 15648 11578 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13740 15660 14105 15688
rect 8846 15580 8852 15632
rect 8904 15580 8910 15632
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 3234 15444 3240 15496
rect 3292 15444 3298 15496
rect 4338 15444 4344 15496
rect 4396 15444 4402 15496
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15484 5963 15487
rect 6178 15484 6184 15496
rect 5951 15456 6184 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8864 15484 8892 15580
rect 12894 15561 12900 15564
rect 12851 15555 12900 15561
rect 12851 15521 12863 15555
rect 12897 15521 12900 15555
rect 12851 15515 12900 15521
rect 12894 15512 12900 15515
rect 12952 15512 12958 15564
rect 12986 15512 12992 15564
rect 13044 15512 13050 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 13228 15524 13277 15552
rect 13228 15512 13234 15524
rect 13265 15521 13277 15524
rect 13311 15552 13323 15555
rect 13630 15552 13636 15564
rect 13311 15524 13636 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 13740 15561 13768 15660
rect 14093 15657 14105 15660
rect 14139 15688 14151 15691
rect 15194 15688 15200 15700
rect 14139 15660 15200 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15562 15648 15568 15700
rect 15620 15648 15626 15700
rect 18046 15648 18052 15700
rect 18104 15648 18110 15700
rect 18322 15648 18328 15700
rect 18380 15648 18386 15700
rect 21177 15691 21235 15697
rect 21177 15657 21189 15691
rect 21223 15688 21235 15691
rect 21358 15688 21364 15700
rect 21223 15660 21364 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 22741 15691 22799 15697
rect 22741 15657 22753 15691
rect 22787 15688 22799 15691
rect 24302 15688 24308 15700
rect 22787 15660 24308 15688
rect 22787 15657 22799 15660
rect 22741 15651 22799 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 25038 15648 25044 15700
rect 25096 15688 25102 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 25096 15660 25145 15688
rect 25096 15648 25102 15660
rect 25133 15657 25145 15660
rect 25179 15657 25191 15691
rect 25133 15651 25191 15657
rect 25498 15648 25504 15700
rect 25556 15688 25562 15700
rect 27617 15691 27675 15697
rect 25556 15660 26832 15688
rect 25556 15648 25562 15660
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 13909 15555 13967 15561
rect 13909 15552 13921 15555
rect 13872 15524 13921 15552
rect 13872 15512 13878 15524
rect 13909 15521 13921 15524
rect 13955 15521 13967 15555
rect 15580 15552 15608 15648
rect 13909 15515 13967 15521
rect 15396 15524 15608 15552
rect 18340 15552 18368 15648
rect 19058 15620 19064 15632
rect 18708 15592 19064 15620
rect 18708 15564 18736 15592
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 20441 15623 20499 15629
rect 20441 15589 20453 15623
rect 20487 15620 20499 15623
rect 20622 15620 20628 15632
rect 20487 15592 20628 15620
rect 20487 15589 20499 15592
rect 20441 15583 20499 15589
rect 20622 15580 20628 15592
rect 20680 15580 20686 15632
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 18340 15524 18521 15552
rect 8159 15456 8892 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9916 15456 10149 15484
rect 9916 15444 9922 15456
rect 10137 15453 10149 15456
rect 10183 15484 10195 15487
rect 10226 15484 10232 15496
rect 10183 15456 10232 15484
rect 10183 15453 10195 15456
rect 10137 15447 10195 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10404 15487 10462 15493
rect 10404 15453 10416 15487
rect 10450 15484 10462 15487
rect 10686 15484 10692 15496
rect 10450 15456 10692 15484
rect 10450 15453 10462 15456
rect 10404 15447 10462 15453
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 15217 15487 15275 15493
rect 15217 15453 15229 15487
rect 15263 15484 15275 15487
rect 15396 15484 15424 15524
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 18509 15515 18567 15521
rect 18690 15512 18696 15564
rect 18748 15512 18754 15564
rect 18874 15512 18880 15564
rect 18932 15552 18938 15564
rect 20027 15555 20085 15561
rect 20027 15552 20039 15555
rect 18932 15524 20039 15552
rect 18932 15512 18938 15524
rect 20027 15521 20039 15524
rect 20073 15521 20085 15555
rect 20027 15515 20085 15521
rect 20162 15512 20168 15564
rect 20220 15512 20226 15564
rect 21821 15555 21879 15561
rect 21821 15521 21833 15555
rect 21867 15552 21879 15555
rect 22094 15552 22100 15564
rect 21867 15524 22100 15552
rect 21867 15521 21879 15524
rect 21821 15515 21879 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 24670 15512 24676 15564
rect 24728 15512 24734 15564
rect 25501 15555 25559 15561
rect 25501 15521 25513 15555
rect 25547 15552 25559 15555
rect 25958 15552 25964 15564
rect 25547 15524 25964 15552
rect 25547 15521 25559 15524
rect 25501 15515 25559 15521
rect 15263 15456 15424 15484
rect 15473 15487 15531 15493
rect 15263 15453 15275 15456
rect 15217 15447 15275 15453
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 16482 15484 16488 15496
rect 15519 15456 15792 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 6454 15416 6460 15428
rect 5736 15388 6460 15416
rect 5736 15360 5764 15388
rect 6454 15376 6460 15388
rect 6512 15416 6518 15428
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 6512 15388 7021 15416
rect 6512 15376 6518 15388
rect 7009 15385 7021 15388
rect 7055 15416 7067 15419
rect 11790 15416 11796 15428
rect 7055 15388 11796 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 15764 15360 15792 15456
rect 16408 15456 16488 15484
rect 2682 15308 2688 15360
rect 2740 15308 2746 15360
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 5258 15308 5264 15360
rect 5316 15308 5322 15360
rect 5718 15308 5724 15360
rect 5776 15308 5782 15360
rect 6086 15308 6092 15360
rect 6144 15308 6150 15360
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7984 15320 8217 15348
rect 7984 15308 7990 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 9582 15308 9588 15360
rect 9640 15348 9646 15360
rect 11974 15348 11980 15360
rect 9640 15320 11980 15348
rect 9640 15308 9646 15320
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 13354 15348 13360 15360
rect 12115 15320 13360 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16408 15357 16436 15456
rect 16482 15444 16488 15456
rect 16540 15484 16546 15496
rect 16850 15493 16856 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16540 15456 16589 15484
rect 16540 15444 16546 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16844 15484 16856 15493
rect 16811 15456 16856 15484
rect 16577 15447 16635 15453
rect 16844 15447 16856 15456
rect 16850 15444 16856 15447
rect 16908 15444 16914 15496
rect 18892 15416 18920 15512
rect 19886 15444 19892 15496
rect 19944 15444 19950 15496
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21450 15484 21456 15496
rect 21131 15456 21456 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 17972 15388 18920 15416
rect 17972 15357 18000 15388
rect 16393 15351 16451 15357
rect 16393 15348 16405 15351
rect 15804 15320 16405 15348
rect 15804 15308 15810 15320
rect 16393 15317 16405 15320
rect 16439 15317 16451 15351
rect 16393 15311 16451 15317
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 18414 15308 18420 15360
rect 18472 15308 18478 15360
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15348 19303 15351
rect 19610 15348 19616 15360
rect 19291 15320 19616 15348
rect 19291 15317 19303 15320
rect 19245 15311 19303 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20916 15348 20944 15447
rect 21450 15444 21456 15456
rect 21508 15484 21514 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 21508 15456 22569 15484
rect 21508 15444 21514 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 23854 15487 23912 15493
rect 23854 15484 23866 15487
rect 23532 15456 23866 15484
rect 23532 15444 23538 15456
rect 23854 15453 23866 15456
rect 23900 15453 23912 15487
rect 23854 15447 23912 15453
rect 24121 15487 24179 15493
rect 24121 15453 24133 15487
rect 24167 15484 24179 15487
rect 25516 15484 25544 15515
rect 25958 15512 25964 15524
rect 26016 15512 26022 15564
rect 26326 15512 26332 15564
rect 26384 15512 26390 15564
rect 26488 15555 26546 15561
rect 26488 15521 26500 15555
rect 26534 15552 26546 15555
rect 26804 15552 26832 15660
rect 27617 15657 27629 15691
rect 27663 15688 27675 15691
rect 28350 15688 28356 15700
rect 27663 15660 28356 15688
rect 27663 15657 27675 15660
rect 27617 15651 27675 15657
rect 26878 15580 26884 15632
rect 26936 15580 26942 15632
rect 26534 15524 26832 15552
rect 27341 15555 27399 15561
rect 26534 15521 26546 15524
rect 26488 15515 26546 15521
rect 27341 15521 27353 15555
rect 27387 15552 27399 15555
rect 27632 15552 27660 15651
rect 28350 15648 28356 15660
rect 28408 15648 28414 15700
rect 31864 15660 33456 15688
rect 31864 15632 31892 15660
rect 31205 15623 31263 15629
rect 31205 15589 31217 15623
rect 31251 15620 31263 15623
rect 31754 15620 31760 15632
rect 31251 15592 31760 15620
rect 31251 15589 31263 15592
rect 31205 15583 31263 15589
rect 31754 15580 31760 15592
rect 31812 15580 31818 15632
rect 31846 15580 31852 15632
rect 31904 15580 31910 15632
rect 27387 15524 27660 15552
rect 31389 15555 31447 15561
rect 27387 15521 27399 15524
rect 27341 15515 27399 15521
rect 31389 15521 31401 15555
rect 31435 15521 31447 15555
rect 32950 15552 32956 15564
rect 31389 15515 31447 15521
rect 32232 15524 32956 15552
rect 24167 15456 25544 15484
rect 24167 15453 24179 15456
rect 24121 15447 24179 15453
rect 26602 15444 26608 15496
rect 26660 15444 26666 15496
rect 27522 15444 27528 15496
rect 27580 15444 27586 15496
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15484 29055 15487
rect 29825 15487 29883 15493
rect 29825 15484 29837 15487
rect 29043 15456 29837 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 24946 15416 24952 15428
rect 24811 15388 24952 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 19852 15320 20944 15348
rect 19852 15308 19858 15320
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21545 15351 21603 15357
rect 21545 15348 21557 15351
rect 21048 15320 21557 15348
rect 21048 15308 21054 15320
rect 21545 15317 21557 15320
rect 21591 15317 21603 15351
rect 21545 15311 21603 15317
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21683 15320 22017 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 26602 15348 26608 15360
rect 25731 15320 26608 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 26602 15308 26608 15320
rect 26660 15308 26666 15360
rect 26694 15308 26700 15360
rect 26752 15348 26758 15360
rect 27540 15348 27568 15444
rect 28752 15419 28810 15425
rect 28752 15385 28764 15419
rect 28798 15416 28810 15419
rect 29178 15416 29184 15428
rect 28798 15388 29184 15416
rect 28798 15385 28810 15388
rect 28752 15379 28810 15385
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 29748 15360 29776 15456
rect 29825 15453 29837 15456
rect 29871 15453 29883 15487
rect 29825 15447 29883 15453
rect 30558 15444 30564 15496
rect 30616 15484 30622 15496
rect 31202 15484 31208 15496
rect 30616 15456 31208 15484
rect 30616 15444 30622 15456
rect 31202 15444 31208 15456
rect 31260 15484 31266 15496
rect 31404 15484 31432 15515
rect 32232 15496 32260 15524
rect 32950 15512 32956 15524
rect 33008 15512 33014 15564
rect 33229 15555 33287 15561
rect 33229 15521 33241 15555
rect 33275 15552 33287 15555
rect 33428 15552 33456 15660
rect 36814 15648 36820 15700
rect 36872 15648 36878 15700
rect 37645 15691 37703 15697
rect 37645 15657 37657 15691
rect 37691 15688 37703 15691
rect 37918 15688 37924 15700
rect 37691 15660 37924 15688
rect 37691 15657 37703 15660
rect 37645 15651 37703 15657
rect 37918 15648 37924 15660
rect 37976 15648 37982 15700
rect 38746 15648 38752 15700
rect 38804 15648 38810 15700
rect 38838 15648 38844 15700
rect 38896 15688 38902 15700
rect 40129 15691 40187 15697
rect 40129 15688 40141 15691
rect 38896 15660 40141 15688
rect 38896 15648 38902 15660
rect 40129 15657 40141 15660
rect 40175 15657 40187 15691
rect 40129 15651 40187 15657
rect 33502 15580 33508 15632
rect 33560 15580 33566 15632
rect 35437 15623 35495 15629
rect 35437 15589 35449 15623
rect 35483 15589 35495 15623
rect 38654 15620 38660 15632
rect 35437 15583 35495 15589
rect 36464 15592 38660 15620
rect 33275 15524 33456 15552
rect 33965 15555 34023 15561
rect 33275 15521 33287 15524
rect 33229 15515 33287 15521
rect 33965 15521 33977 15555
rect 34011 15552 34023 15555
rect 34514 15552 34520 15564
rect 34011 15524 34520 15552
rect 34011 15521 34023 15524
rect 33965 15515 34023 15521
rect 34514 15512 34520 15524
rect 34572 15512 34578 15564
rect 34885 15555 34943 15561
rect 34885 15521 34897 15555
rect 34931 15552 34943 15555
rect 35158 15552 35164 15564
rect 34931 15524 35164 15552
rect 34931 15521 34943 15524
rect 34885 15515 34943 15521
rect 35158 15512 35164 15524
rect 35216 15512 35222 15564
rect 35452 15552 35480 15583
rect 36081 15555 36139 15561
rect 36081 15552 36093 15555
rect 35452 15524 36093 15552
rect 36081 15521 36093 15524
rect 36127 15521 36139 15555
rect 36081 15515 36139 15521
rect 31260 15456 31432 15484
rect 31260 15444 31266 15456
rect 32214 15444 32220 15496
rect 32272 15444 32278 15496
rect 33134 15493 33140 15496
rect 33112 15487 33140 15493
rect 33112 15453 33124 15487
rect 33112 15447 33140 15453
rect 33134 15444 33140 15447
rect 33192 15444 33198 15496
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15484 34207 15487
rect 34330 15484 34336 15496
rect 34195 15456 34336 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 34330 15444 34336 15456
rect 34388 15444 34394 15496
rect 35176 15484 35204 15512
rect 36464 15493 36492 15592
rect 38654 15580 38660 15592
rect 38712 15580 38718 15632
rect 36906 15512 36912 15564
rect 36964 15512 36970 15564
rect 37369 15555 37427 15561
rect 37369 15521 37381 15555
rect 37415 15521 37427 15555
rect 37369 15515 37427 15521
rect 36449 15487 36507 15493
rect 36449 15484 36461 15487
rect 35176 15456 36461 15484
rect 36449 15453 36461 15456
rect 36495 15453 36507 15487
rect 36924 15484 36952 15512
rect 37185 15487 37243 15493
rect 37185 15484 37197 15487
rect 36924 15456 37197 15484
rect 36449 15447 36507 15453
rect 37185 15453 37197 15456
rect 37231 15453 37243 15487
rect 37185 15447 37243 15453
rect 30092 15419 30150 15425
rect 30092 15385 30104 15419
rect 30138 15416 30150 15419
rect 31294 15416 31300 15428
rect 30138 15388 31300 15416
rect 30138 15385 30150 15388
rect 30092 15379 30150 15385
rect 31294 15376 31300 15388
rect 31352 15376 31358 15428
rect 34790 15416 34796 15428
rect 34440 15388 34796 15416
rect 26752 15320 27568 15348
rect 29365 15351 29423 15357
rect 26752 15308 26758 15320
rect 29365 15317 29377 15351
rect 29411 15348 29423 15351
rect 29730 15348 29736 15360
rect 29411 15320 29736 15348
rect 29411 15317 29423 15320
rect 29365 15311 29423 15317
rect 29730 15308 29736 15320
rect 29788 15308 29794 15360
rect 30834 15308 30840 15360
rect 30892 15348 30898 15360
rect 31573 15351 31631 15357
rect 31573 15348 31585 15351
rect 30892 15320 31585 15348
rect 30892 15308 30898 15320
rect 31573 15317 31585 15320
rect 31619 15317 31631 15351
rect 31573 15311 31631 15317
rect 31665 15351 31723 15357
rect 31665 15317 31677 15351
rect 31711 15348 31723 15351
rect 31938 15348 31944 15360
rect 31711 15320 31944 15348
rect 31711 15317 31723 15320
rect 31665 15311 31723 15317
rect 31938 15308 31944 15320
rect 31996 15308 32002 15360
rect 32030 15308 32036 15360
rect 32088 15308 32094 15360
rect 32309 15351 32367 15357
rect 32309 15317 32321 15351
rect 32355 15348 32367 15351
rect 34440 15348 34468 15388
rect 34790 15376 34796 15388
rect 34848 15376 34854 15428
rect 37384 15416 37412 15515
rect 37458 15512 37464 15564
rect 37516 15552 37522 15564
rect 38197 15555 38255 15561
rect 38197 15552 38209 15555
rect 37516 15524 38209 15552
rect 37516 15512 37522 15524
rect 38197 15521 38209 15524
rect 38243 15521 38255 15555
rect 38197 15515 38255 15521
rect 38013 15487 38071 15493
rect 38013 15453 38025 15487
rect 38059 15484 38071 15487
rect 38764 15484 38792 15648
rect 40144 15552 40172 15651
rect 42610 15648 42616 15700
rect 42668 15688 42674 15700
rect 43438 15688 43444 15700
rect 42668 15660 43444 15688
rect 42668 15648 42674 15660
rect 43438 15648 43444 15660
rect 43496 15648 43502 15700
rect 44358 15688 44364 15700
rect 43640 15660 44364 15688
rect 41693 15623 41751 15629
rect 41693 15589 41705 15623
rect 41739 15620 41751 15623
rect 43254 15620 43260 15632
rect 41739 15592 43260 15620
rect 41739 15589 41751 15592
rect 41693 15583 41751 15589
rect 40313 15555 40371 15561
rect 40313 15552 40325 15555
rect 40144 15524 40325 15552
rect 40313 15521 40325 15524
rect 40359 15521 40371 15555
rect 40313 15515 40371 15521
rect 42150 15512 42156 15564
rect 42208 15552 42214 15564
rect 43180 15561 43208 15592
rect 43254 15580 43260 15592
rect 43312 15580 43318 15632
rect 42337 15555 42395 15561
rect 42337 15552 42349 15555
rect 42208 15524 42349 15552
rect 42208 15512 42214 15524
rect 42337 15521 42349 15524
rect 42383 15521 42395 15555
rect 42337 15515 42395 15521
rect 43165 15555 43223 15561
rect 43165 15521 43177 15555
rect 43211 15521 43223 15555
rect 43165 15515 43223 15521
rect 43530 15512 43536 15564
rect 43588 15512 43594 15564
rect 43640 15561 43668 15660
rect 44358 15648 44364 15660
rect 44416 15648 44422 15700
rect 49053 15691 49111 15697
rect 49053 15657 49065 15691
rect 49099 15688 49111 15691
rect 49142 15688 49148 15700
rect 49099 15660 49148 15688
rect 49099 15657 49111 15660
rect 49053 15651 49111 15657
rect 49142 15648 49148 15660
rect 49200 15688 49206 15700
rect 49602 15688 49608 15700
rect 49200 15660 49608 15688
rect 49200 15648 49206 15660
rect 49602 15648 49608 15660
rect 49660 15648 49666 15700
rect 49970 15648 49976 15700
rect 50028 15648 50034 15700
rect 54202 15648 54208 15700
rect 54260 15648 54266 15700
rect 54297 15691 54355 15697
rect 54297 15657 54309 15691
rect 54343 15688 54355 15691
rect 54662 15688 54668 15700
rect 54343 15660 54668 15688
rect 54343 15657 54355 15660
rect 54297 15651 54355 15657
rect 54662 15648 54668 15660
rect 54720 15648 54726 15700
rect 55416 15660 56824 15688
rect 44085 15623 44143 15629
rect 44085 15589 44097 15623
rect 44131 15620 44143 15623
rect 44131 15592 44772 15620
rect 44131 15589 44143 15592
rect 44085 15583 44143 15589
rect 44744 15561 44772 15592
rect 43625 15555 43683 15561
rect 43625 15521 43637 15555
rect 43671 15521 43683 15555
rect 43625 15515 43683 15521
rect 44729 15555 44787 15561
rect 44729 15521 44741 15555
rect 44775 15521 44787 15555
rect 44729 15515 44787 15521
rect 49421 15555 49479 15561
rect 49421 15521 49433 15555
rect 49467 15552 49479 15555
rect 50341 15555 50399 15561
rect 50341 15552 50353 15555
rect 49467 15524 50353 15552
rect 49467 15521 49479 15524
rect 49421 15515 49479 15521
rect 50341 15521 50353 15524
rect 50387 15552 50399 15555
rect 50387 15524 51074 15552
rect 50387 15521 50399 15524
rect 50341 15515 50399 15521
rect 38059 15456 38792 15484
rect 38059 15453 38071 15456
rect 38013 15447 38071 15453
rect 42242 15444 42248 15496
rect 42300 15484 42306 15496
rect 43717 15487 43775 15493
rect 43717 15484 43729 15487
rect 42300 15456 43729 15484
rect 42300 15444 42306 15456
rect 43717 15453 43729 15456
rect 43763 15484 43775 15487
rect 45370 15484 45376 15496
rect 43763 15456 45376 15484
rect 43763 15453 43775 15456
rect 43717 15447 43775 15453
rect 45370 15444 45376 15456
rect 45428 15444 45434 15496
rect 45554 15444 45560 15496
rect 45612 15484 45618 15496
rect 46201 15487 46259 15493
rect 46201 15484 46213 15487
rect 45612 15456 46213 15484
rect 45612 15444 45618 15456
rect 46201 15453 46213 15456
rect 46247 15484 46259 15487
rect 46290 15484 46296 15496
rect 46247 15456 46296 15484
rect 46247 15453 46259 15456
rect 46201 15447 46259 15453
rect 46290 15444 46296 15456
rect 46348 15484 46354 15496
rect 46842 15484 46848 15496
rect 46348 15456 46848 15484
rect 46348 15444 46354 15456
rect 46842 15444 46848 15456
rect 46900 15484 46906 15496
rect 47673 15487 47731 15493
rect 47673 15484 47685 15487
rect 46900 15456 47685 15484
rect 46900 15444 46906 15456
rect 47673 15453 47685 15456
rect 47719 15453 47731 15487
rect 47673 15447 47731 15453
rect 47940 15487 47998 15493
rect 47940 15453 47952 15487
rect 47986 15484 47998 15487
rect 48222 15484 48228 15496
rect 47986 15456 48228 15484
rect 47986 15453 47998 15456
rect 47940 15447 47998 15453
rect 48222 15444 48228 15456
rect 48280 15444 48286 15496
rect 49694 15444 49700 15496
rect 49752 15484 49758 15496
rect 50617 15487 50675 15493
rect 50617 15484 50629 15487
rect 49752 15456 50629 15484
rect 49752 15444 49758 15456
rect 50617 15453 50629 15456
rect 50663 15453 50675 15487
rect 50617 15447 50675 15453
rect 50706 15444 50712 15496
rect 50764 15444 50770 15496
rect 36556 15388 37412 15416
rect 40580 15419 40638 15425
rect 36556 15360 36584 15388
rect 40580 15385 40592 15419
rect 40626 15416 40638 15419
rect 41230 15416 41236 15428
rect 40626 15388 41236 15416
rect 40626 15385 40638 15388
rect 40580 15379 40638 15385
rect 41230 15376 41236 15388
rect 41288 15376 41294 15428
rect 42153 15419 42211 15425
rect 42153 15385 42165 15419
rect 42199 15416 42211 15419
rect 42613 15419 42671 15425
rect 42613 15416 42625 15419
rect 42199 15388 42625 15416
rect 42199 15385 42211 15388
rect 42153 15379 42211 15385
rect 42613 15385 42625 15388
rect 42659 15385 42671 15419
rect 42613 15379 42671 15385
rect 43070 15376 43076 15428
rect 43128 15416 43134 15428
rect 45738 15416 45744 15428
rect 43128 15388 45744 15416
rect 43128 15376 43134 15388
rect 45738 15376 45744 15388
rect 45796 15376 45802 15428
rect 46468 15419 46526 15425
rect 46468 15385 46480 15419
rect 46514 15416 46526 15419
rect 46750 15416 46756 15428
rect 46514 15388 46756 15416
rect 46514 15385 46526 15388
rect 46468 15379 46526 15385
rect 46750 15376 46756 15388
rect 46808 15376 46814 15428
rect 48038 15376 48044 15428
rect 48096 15416 48102 15428
rect 49513 15419 49571 15425
rect 48096 15388 49464 15416
rect 48096 15376 48102 15388
rect 32355 15320 34468 15348
rect 34517 15351 34575 15357
rect 32355 15317 32367 15320
rect 32309 15311 32367 15317
rect 34517 15317 34529 15351
rect 34563 15348 34575 15351
rect 34882 15348 34888 15360
rect 34563 15320 34888 15348
rect 34563 15317 34575 15320
rect 34517 15311 34575 15317
rect 34882 15308 34888 15320
rect 34940 15308 34946 15360
rect 34974 15308 34980 15360
rect 35032 15308 35038 15360
rect 35066 15308 35072 15360
rect 35124 15308 35130 15360
rect 35526 15308 35532 15360
rect 35584 15308 35590 15360
rect 36538 15308 36544 15360
rect 36596 15308 36602 15360
rect 37277 15351 37335 15357
rect 37277 15317 37289 15351
rect 37323 15348 37335 15351
rect 37550 15348 37556 15360
rect 37323 15320 37556 15348
rect 37323 15317 37335 15320
rect 37277 15311 37335 15317
rect 37550 15308 37556 15320
rect 37608 15348 37614 15360
rect 38105 15351 38163 15357
rect 38105 15348 38117 15351
rect 37608 15320 38117 15348
rect 37608 15308 37614 15320
rect 38105 15317 38117 15320
rect 38151 15348 38163 15351
rect 38654 15348 38660 15360
rect 38151 15320 38660 15348
rect 38151 15317 38163 15320
rect 38105 15311 38163 15317
rect 38654 15308 38660 15320
rect 38712 15308 38718 15360
rect 41782 15308 41788 15360
rect 41840 15308 41846 15360
rect 44177 15351 44235 15357
rect 44177 15317 44189 15351
rect 44223 15348 44235 15351
rect 44634 15348 44640 15360
rect 44223 15320 44640 15348
rect 44223 15317 44235 15320
rect 44177 15311 44235 15317
rect 44634 15308 44640 15320
rect 44692 15308 44698 15360
rect 45756 15348 45784 15376
rect 46198 15348 46204 15360
rect 45756 15320 46204 15348
rect 46198 15308 46204 15320
rect 46256 15308 46262 15360
rect 47581 15351 47639 15357
rect 47581 15317 47593 15351
rect 47627 15348 47639 15351
rect 49050 15348 49056 15360
rect 47627 15320 49056 15348
rect 47627 15317 47639 15320
rect 47581 15311 47639 15317
rect 49050 15308 49056 15320
rect 49108 15308 49114 15360
rect 49436 15348 49464 15388
rect 49513 15385 49525 15419
rect 49559 15416 49571 15419
rect 50724 15416 50752 15444
rect 49559 15388 50752 15416
rect 49559 15385 49571 15388
rect 49513 15379 49571 15385
rect 49605 15351 49663 15357
rect 49605 15348 49617 15351
rect 49436 15320 49617 15348
rect 49605 15317 49617 15320
rect 49651 15348 49663 15351
rect 50430 15348 50436 15360
rect 49651 15320 50436 15348
rect 49651 15317 49663 15320
rect 49605 15311 49663 15317
rect 50430 15308 50436 15320
rect 50488 15308 50494 15360
rect 51046 15348 51074 15524
rect 54846 15512 54852 15564
rect 54904 15512 54910 15564
rect 52365 15487 52423 15493
rect 52365 15453 52377 15487
rect 52411 15484 52423 15487
rect 52733 15487 52791 15493
rect 52733 15484 52745 15487
rect 52411 15456 52745 15484
rect 52411 15453 52423 15456
rect 52365 15447 52423 15453
rect 52733 15453 52745 15456
rect 52779 15484 52791 15487
rect 52825 15487 52883 15493
rect 52825 15484 52837 15487
rect 52779 15456 52837 15484
rect 52779 15453 52791 15456
rect 52733 15447 52791 15453
rect 52825 15453 52837 15456
rect 52871 15484 52883 15487
rect 54665 15487 54723 15493
rect 52871 15456 53236 15484
rect 52871 15453 52883 15456
rect 52825 15447 52883 15453
rect 53208 15428 53236 15456
rect 54665 15453 54677 15487
rect 54711 15484 54723 15487
rect 55416 15484 55444 15660
rect 56796 15632 56824 15660
rect 57238 15648 57244 15700
rect 57296 15688 57302 15700
rect 57698 15688 57704 15700
rect 57296 15660 57704 15688
rect 57296 15648 57302 15660
rect 57698 15648 57704 15660
rect 57756 15648 57762 15700
rect 57882 15648 57888 15700
rect 57940 15648 57946 15700
rect 56778 15580 56784 15632
rect 56836 15580 56842 15632
rect 56888 15592 57468 15620
rect 55766 15512 55772 15564
rect 55824 15552 55830 15564
rect 55824 15524 55996 15552
rect 55824 15512 55830 15524
rect 55968 15493 55996 15524
rect 56042 15512 56048 15564
rect 56100 15561 56106 15564
rect 56100 15555 56149 15561
rect 56100 15521 56103 15555
rect 56137 15521 56149 15555
rect 56100 15515 56149 15521
rect 56100 15512 56106 15515
rect 56502 15512 56508 15564
rect 56560 15512 56566 15564
rect 56594 15512 56600 15564
rect 56652 15552 56658 15564
rect 56888 15552 56916 15592
rect 56652 15524 56916 15552
rect 56652 15512 56658 15524
rect 57146 15512 57152 15564
rect 57204 15512 57210 15564
rect 57238 15512 57244 15564
rect 57296 15512 57302 15564
rect 57440 15561 57468 15592
rect 57425 15555 57483 15561
rect 57425 15521 57437 15555
rect 57471 15521 57483 15555
rect 57425 15515 57483 15521
rect 57517 15555 57575 15561
rect 57517 15521 57529 15555
rect 57563 15552 57575 15555
rect 57900 15552 57928 15648
rect 57563 15524 57928 15552
rect 57563 15521 57575 15524
rect 57517 15515 57575 15521
rect 54711 15456 55444 15484
rect 55953 15487 56011 15493
rect 54711 15453 54723 15456
rect 54665 15447 54723 15453
rect 55953 15453 55965 15487
rect 55999 15453 56011 15487
rect 55953 15447 56011 15453
rect 53098 15425 53104 15428
rect 53092 15416 53104 15425
rect 53059 15388 53104 15416
rect 53092 15379 53104 15388
rect 53098 15376 53104 15379
rect 53156 15376 53162 15428
rect 53190 15376 53196 15428
rect 53248 15376 53254 15428
rect 53742 15376 53748 15428
rect 53800 15416 53806 15428
rect 54680 15416 54708 15447
rect 56226 15444 56232 15496
rect 56284 15444 56290 15496
rect 56965 15487 57023 15493
rect 56965 15453 56977 15487
rect 57011 15484 57023 15487
rect 57256 15484 57284 15512
rect 57011 15456 57284 15484
rect 57011 15453 57023 15456
rect 56965 15447 57023 15453
rect 53800 15388 54708 15416
rect 57440 15416 57468 15515
rect 58253 15419 58311 15425
rect 58253 15416 58265 15419
rect 57440 15388 58265 15416
rect 53800 15376 53806 15388
rect 58253 15385 58265 15388
rect 58299 15385 58311 15419
rect 58253 15379 58311 15385
rect 54478 15348 54484 15360
rect 51046 15320 54484 15348
rect 54478 15308 54484 15320
rect 54536 15308 54542 15360
rect 54754 15308 54760 15360
rect 54812 15308 54818 15360
rect 55309 15351 55367 15357
rect 55309 15317 55321 15351
rect 55355 15348 55367 15351
rect 56318 15348 56324 15360
rect 55355 15320 56324 15348
rect 55355 15317 55367 15320
rect 55309 15311 55367 15317
rect 56318 15308 56324 15320
rect 56376 15308 56382 15360
rect 56778 15308 56784 15360
rect 56836 15348 56842 15360
rect 57609 15351 57667 15357
rect 57609 15348 57621 15351
rect 56836 15320 57621 15348
rect 56836 15308 56842 15320
rect 57609 15317 57621 15320
rect 57655 15317 57667 15351
rect 57609 15311 57667 15317
rect 57974 15308 57980 15360
rect 58032 15308 58038 15360
rect 1104 15258 59040 15280
rect 1104 15206 15394 15258
rect 15446 15206 15458 15258
rect 15510 15206 15522 15258
rect 15574 15206 15586 15258
rect 15638 15206 15650 15258
rect 15702 15206 29838 15258
rect 29890 15206 29902 15258
rect 29954 15206 29966 15258
rect 30018 15206 30030 15258
rect 30082 15206 30094 15258
rect 30146 15206 44282 15258
rect 44334 15206 44346 15258
rect 44398 15206 44410 15258
rect 44462 15206 44474 15258
rect 44526 15206 44538 15258
rect 44590 15206 58726 15258
rect 58778 15206 58790 15258
rect 58842 15206 58854 15258
rect 58906 15206 58918 15258
rect 58970 15206 58982 15258
rect 59034 15206 59040 15258
rect 1104 15184 59040 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3234 15144 3240 15156
rect 3007 15116 3240 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3329 15147 3387 15153
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3786 15144 3792 15156
rect 3375 15116 3792 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 3970 15104 3976 15156
rect 4028 15104 4034 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 6086 15144 6092 15156
rect 5767 15116 6092 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 6178 15104 6184 15156
rect 6236 15104 6242 15156
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 6420 15116 6745 15144
rect 6420 15104 6426 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 7742 15144 7748 15156
rect 7515 15116 7748 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 3421 15079 3479 15085
rect 3421 15045 3433 15079
rect 3467 15076 3479 15079
rect 3988 15076 4016 15104
rect 3467 15048 5856 15076
rect 3467 15045 3479 15048
rect 3421 15039 3479 15045
rect 5828 15020 5856 15048
rect 5810 14968 5816 15020
rect 5868 14968 5874 15020
rect 7484 15008 7512 15107
rect 7742 15104 7748 15116
rect 7800 15144 7806 15156
rect 10042 15144 10048 15156
rect 7800 15116 10048 15144
rect 7800 15104 7806 15116
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11388 15116 11529 15144
rect 11388 15104 11394 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11882 15104 11888 15156
rect 11940 15104 11946 15156
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12710 15144 12716 15156
rect 12032 15116 12716 15144
rect 12032 15104 12038 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15144 13231 15147
rect 13814 15144 13820 15156
rect 13219 15116 13820 15144
rect 13219 15113 13231 15116
rect 13173 15107 13231 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14200 15116 17080 15144
rect 10220 15079 10278 15085
rect 10220 15045 10232 15079
rect 10266 15076 10278 15079
rect 10870 15076 10876 15088
rect 10266 15048 10876 15076
rect 10266 15045 10278 15048
rect 10220 15039 10278 15045
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 12250 15076 12256 15088
rect 11112 15048 12256 15076
rect 11112 15036 11118 15048
rect 12250 15036 12256 15048
rect 12308 15076 12314 15088
rect 14200 15076 14228 15116
rect 12308 15048 14228 15076
rect 14308 15079 14366 15085
rect 12308 15036 12314 15048
rect 14308 15045 14320 15079
rect 14354 15076 14366 15079
rect 14734 15076 14740 15088
rect 14354 15048 14740 15076
rect 14354 15045 14366 15048
rect 14308 15039 14366 15045
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 17052 15085 17080 15116
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 17865 15147 17923 15153
rect 17865 15144 17877 15147
rect 17736 15116 17877 15144
rect 17736 15104 17742 15116
rect 17865 15113 17877 15116
rect 17911 15113 17923 15147
rect 17865 15107 17923 15113
rect 18690 15104 18696 15156
rect 18748 15104 18754 15156
rect 18782 15104 18788 15156
rect 18840 15144 18846 15156
rect 19153 15147 19211 15153
rect 19153 15144 19165 15147
rect 18840 15116 19165 15144
rect 18840 15104 18846 15116
rect 19153 15113 19165 15116
rect 19199 15113 19211 15147
rect 19153 15107 19211 15113
rect 17037 15079 17095 15085
rect 17037 15045 17049 15079
rect 17083 15076 17095 15079
rect 18708 15076 18736 15104
rect 17083 15048 18736 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 6472 14980 7512 15008
rect 11977 15011 12035 15017
rect 2866 14900 2872 14952
rect 2924 14900 2930 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 4154 14940 4160 14952
rect 3651 14912 4160 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 4356 14872 4384 14903
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 5629 14943 5687 14949
rect 4764 14912 5580 14940
rect 4764 14900 4770 14912
rect 5350 14872 5356 14884
rect 3528 14844 5356 14872
rect 3528 14816 3556 14844
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 5552 14872 5580 14912
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 5718 14940 5724 14952
rect 5675 14912 5724 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6472 14949 6500 14980
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 12023 14980 12357 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 13722 15008 13728 15020
rect 13136 14980 13728 15008
rect 13136 14968 13142 14980
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 17957 15011 18015 15017
rect 17957 15008 17969 15011
rect 17543 14980 17969 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 17957 14977 17969 14980
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 15008 18659 15011
rect 18874 15008 18880 15020
rect 18647 14980 18880 15008
rect 18647 14977 18659 14980
rect 18601 14971 18659 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 19168 15008 19196 15107
rect 21082 15104 21088 15156
rect 21140 15104 21146 15156
rect 21450 15104 21456 15156
rect 21508 15104 21514 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15144 23535 15147
rect 23750 15144 23756 15156
rect 23523 15116 23756 15144
rect 23523 15113 23535 15116
rect 23477 15107 23535 15113
rect 23750 15104 23756 15116
rect 23808 15144 23814 15156
rect 24578 15144 24584 15156
rect 23808 15116 24584 15144
rect 23808 15104 23814 15116
rect 24578 15104 24584 15116
rect 24636 15104 24642 15156
rect 24949 15147 25007 15153
rect 24949 15113 24961 15147
rect 24995 15144 25007 15147
rect 25498 15144 25504 15156
rect 24995 15116 25504 15144
rect 24995 15113 25007 15116
rect 24949 15107 25007 15113
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 25774 15104 25780 15156
rect 25832 15144 25838 15156
rect 25832 15116 26280 15144
rect 25832 15104 25838 15116
rect 20340 15079 20398 15085
rect 20340 15045 20352 15079
rect 20386 15076 20398 15079
rect 20714 15076 20720 15088
rect 20386 15048 20720 15076
rect 20386 15045 20398 15048
rect 20340 15039 20398 15045
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 21100 15076 21128 15104
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21100 15048 21833 15076
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 23836 15079 23894 15085
rect 23836 15045 23848 15079
rect 23882 15076 23894 15079
rect 24394 15076 24400 15088
rect 23882 15048 24400 15076
rect 23882 15045 23894 15048
rect 23836 15039 23894 15045
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 25332 15048 26096 15076
rect 20070 15008 20076 15020
rect 19168 14980 20076 15008
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 25332 15017 25360 15048
rect 26068 15020 26096 15048
rect 25590 15017 25596 15020
rect 25317 15011 25375 15017
rect 22520 14980 24716 15008
rect 22520 14968 22526 14980
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 6546 14900 6552 14952
rect 6604 14940 6610 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 6604 14912 6653 14940
rect 6604 14900 6610 14912
rect 6641 14909 6653 14912
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 8570 14900 8576 14952
rect 8628 14900 8634 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9916 14912 9965 14940
rect 9916 14900 9922 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 11698 14940 11704 14952
rect 9953 14903 10011 14909
rect 10980 14912 11704 14940
rect 5552 14844 9996 14872
rect 2222 14764 2228 14816
rect 2280 14764 2286 14816
rect 3510 14764 3516 14816
rect 3568 14764 3574 14816
rect 3786 14764 3792 14816
rect 3844 14764 3850 14816
rect 7098 14764 7104 14816
rect 7156 14764 7162 14816
rect 8018 14764 8024 14816
rect 8076 14764 8082 14816
rect 9968 14804 9996 14844
rect 10980 14804 11008 14912
rect 11698 14900 11704 14912
rect 11756 14940 11762 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11756 14912 12081 14940
rect 11756 14900 11762 14912
rect 12069 14909 12081 14912
rect 12115 14940 12127 14943
rect 12250 14940 12256 14952
rect 12115 14912 12256 14940
rect 12115 14909 12127 14912
rect 12069 14903 12127 14909
rect 12250 14900 12256 14912
rect 12308 14940 12314 14952
rect 13096 14940 13124 14968
rect 12308 14912 13124 14940
rect 14553 14943 14611 14949
rect 12308 14900 12314 14912
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 15746 14940 15752 14952
rect 14599 14912 15752 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 11333 14875 11391 14881
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 12342 14872 12348 14884
rect 11379 14844 12348 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 14936 14816 14964 14912
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17405 14943 17463 14949
rect 17267 14912 17301 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17405 14909 17417 14943
rect 17451 14940 17463 14943
rect 18414 14940 18420 14952
rect 17451 14912 18420 14940
rect 17451 14909 17463 14912
rect 17405 14903 17463 14909
rect 16485 14875 16543 14881
rect 16485 14841 16497 14875
rect 16531 14872 16543 14875
rect 17126 14872 17132 14884
rect 16531 14844 17132 14872
rect 16531 14841 16543 14844
rect 16485 14835 16543 14841
rect 17126 14832 17132 14844
rect 17184 14872 17190 14884
rect 17236 14872 17264 14903
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 19150 14900 19156 14952
rect 19208 14900 19214 14952
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14940 19487 14943
rect 19794 14940 19800 14952
rect 19475 14912 19800 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 22370 14900 22376 14952
rect 22428 14900 22434 14952
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 19168 14872 19196 14900
rect 17184 14844 19196 14872
rect 17184 14832 17190 14844
rect 9968 14776 11008 14804
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 19978 14764 19984 14816
rect 20036 14764 20042 14816
rect 23584 14804 23612 14903
rect 23934 14804 23940 14816
rect 23584 14776 23940 14804
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 24688 14804 24716 14980
rect 25317 14977 25329 15011
rect 25363 14977 25375 15011
rect 25584 15008 25596 15017
rect 25551 14980 25596 15008
rect 25317 14971 25375 14977
rect 25584 14971 25596 14980
rect 25590 14968 25596 14971
rect 25648 14968 25654 15020
rect 26050 14968 26056 15020
rect 26108 14968 26114 15020
rect 26252 15008 26280 15116
rect 26694 15104 26700 15156
rect 26752 15104 26758 15156
rect 27798 15104 27804 15156
rect 27856 15144 27862 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 27856 15116 27905 15144
rect 27856 15104 27862 15116
rect 27893 15113 27905 15116
rect 27939 15113 27951 15147
rect 27893 15107 27951 15113
rect 29178 15104 29184 15156
rect 29236 15104 29242 15156
rect 31294 15104 31300 15156
rect 31352 15104 31358 15156
rect 31938 15104 31944 15156
rect 31996 15144 32002 15156
rect 32125 15147 32183 15153
rect 32125 15144 32137 15147
rect 31996 15116 32137 15144
rect 31996 15104 32002 15116
rect 32125 15113 32137 15116
rect 32171 15113 32183 15147
rect 32125 15107 32183 15113
rect 34698 15104 34704 15156
rect 34756 15144 34762 15156
rect 34793 15147 34851 15153
rect 34793 15144 34805 15147
rect 34756 15116 34805 15144
rect 34756 15104 34762 15116
rect 34793 15113 34805 15116
rect 34839 15113 34851 15147
rect 34793 15107 34851 15113
rect 34974 15104 34980 15156
rect 35032 15144 35038 15156
rect 35253 15147 35311 15153
rect 35253 15144 35265 15147
rect 35032 15116 35265 15144
rect 35032 15104 35038 15116
rect 35253 15113 35265 15116
rect 35299 15113 35311 15147
rect 35253 15107 35311 15113
rect 36722 15104 36728 15156
rect 36780 15144 36786 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 36780 15116 37841 15144
rect 36780 15104 36786 15116
rect 37829 15113 37841 15116
rect 37875 15144 37887 15147
rect 38010 15144 38016 15156
rect 37875 15116 38016 15144
rect 37875 15113 37887 15116
rect 37829 15107 37887 15113
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 41230 15104 41236 15156
rect 41288 15104 41294 15156
rect 42889 15147 42947 15153
rect 42889 15113 42901 15147
rect 42935 15144 42947 15147
rect 43530 15144 43536 15156
rect 42935 15116 43536 15144
rect 42935 15113 42947 15116
rect 42889 15107 42947 15113
rect 43530 15104 43536 15116
rect 43588 15104 43594 15156
rect 44729 15147 44787 15153
rect 44729 15113 44741 15147
rect 44775 15144 44787 15147
rect 45554 15144 45560 15156
rect 44775 15116 45560 15144
rect 44775 15113 44787 15116
rect 44729 15107 44787 15113
rect 30092 15079 30150 15085
rect 30092 15045 30104 15079
rect 30138 15076 30150 15079
rect 30282 15076 30288 15088
rect 30138 15048 30288 15076
rect 30138 15045 30150 15048
rect 30092 15039 30150 15045
rect 30282 15036 30288 15048
rect 30340 15036 30346 15088
rect 33220 15079 33278 15085
rect 33220 15045 33232 15079
rect 33266 15076 33278 15079
rect 35526 15076 35532 15088
rect 33266 15048 35532 15076
rect 33266 15045 33278 15048
rect 33220 15039 33278 15045
rect 35526 15036 35532 15048
rect 35584 15036 35590 15088
rect 41386 15048 44404 15076
rect 27801 15011 27859 15017
rect 27801 15008 27813 15011
rect 26252 14980 27813 15008
rect 27801 14977 27813 14980
rect 27847 15008 27859 15011
rect 27890 15008 27896 15020
rect 27847 14980 27896 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 27890 14968 27896 14980
rect 27948 14968 27954 15020
rect 31941 15011 31999 15017
rect 31941 14977 31953 15011
rect 31987 15008 31999 15011
rect 32030 15008 32036 15020
rect 31987 14980 32036 15008
rect 31987 14977 31999 14980
rect 31941 14971 31999 14977
rect 32030 14968 32036 14980
rect 32088 14968 32094 15020
rect 33042 15008 33048 15020
rect 32692 14980 33048 15008
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27356 14912 27629 14940
rect 26694 14804 26700 14816
rect 24688 14776 26700 14804
rect 26694 14764 26700 14776
rect 26752 14804 26758 14816
rect 27356 14813 27384 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 28537 14943 28595 14949
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 28537 14903 28595 14909
rect 28261 14875 28319 14881
rect 28261 14841 28273 14875
rect 28307 14872 28319 14875
rect 28552 14872 28580 14903
rect 29730 14900 29736 14952
rect 29788 14940 29794 14952
rect 29825 14943 29883 14949
rect 29825 14940 29837 14943
rect 29788 14912 29837 14940
rect 29788 14900 29794 14912
rect 29825 14909 29837 14912
rect 29871 14909 29883 14943
rect 29825 14903 29883 14909
rect 31754 14900 31760 14952
rect 31812 14940 31818 14952
rect 32692 14949 32720 14980
rect 33042 14968 33048 14980
rect 33100 14968 33106 15020
rect 37458 15008 37464 15020
rect 34624 14980 37464 15008
rect 32677 14943 32735 14949
rect 32677 14940 32689 14943
rect 31812 14912 32689 14940
rect 31812 14900 31818 14912
rect 32677 14909 32689 14912
rect 32723 14909 32735 14943
rect 32677 14903 32735 14909
rect 32858 14900 32864 14952
rect 32916 14940 32922 14952
rect 34624 14949 34652 14980
rect 37458 14968 37464 14980
rect 37516 14968 37522 15020
rect 32953 14943 33011 14949
rect 32953 14940 32965 14943
rect 32916 14912 32965 14940
rect 32916 14900 32922 14912
rect 32953 14909 32965 14912
rect 32999 14909 33011 14943
rect 32953 14903 33011 14909
rect 34609 14943 34667 14949
rect 34609 14909 34621 14943
rect 34655 14909 34667 14943
rect 34609 14903 34667 14909
rect 34701 14943 34759 14949
rect 34701 14909 34713 14943
rect 34747 14940 34759 14943
rect 35066 14940 35072 14952
rect 34747 14912 35072 14940
rect 34747 14909 34759 14912
rect 34701 14903 34759 14909
rect 28307 14844 28580 14872
rect 31205 14875 31263 14881
rect 28307 14841 28319 14844
rect 28261 14835 28319 14841
rect 31205 14841 31217 14875
rect 31251 14872 31263 14875
rect 31846 14872 31852 14884
rect 31251 14844 31852 14872
rect 31251 14841 31263 14844
rect 31205 14835 31263 14841
rect 31846 14832 31852 14844
rect 31904 14832 31910 14884
rect 34624 14872 34652 14903
rect 35066 14900 35072 14912
rect 35124 14900 35130 14952
rect 35618 14900 35624 14952
rect 35676 14900 35682 14952
rect 35805 14943 35863 14949
rect 35805 14909 35817 14943
rect 35851 14909 35863 14943
rect 35805 14903 35863 14909
rect 34882 14872 34888 14884
rect 34624 14844 34888 14872
rect 34882 14832 34888 14844
rect 34940 14832 34946 14884
rect 35161 14875 35219 14881
rect 35161 14841 35173 14875
rect 35207 14872 35219 14875
rect 35636 14872 35664 14900
rect 35207 14844 35664 14872
rect 35207 14841 35219 14844
rect 35161 14835 35219 14841
rect 27341 14807 27399 14813
rect 27341 14804 27353 14807
rect 26752 14776 27353 14804
rect 26752 14764 26758 14776
rect 27341 14773 27353 14776
rect 27387 14773 27399 14807
rect 27341 14767 27399 14773
rect 34330 14764 34336 14816
rect 34388 14804 34394 14816
rect 35820 14804 35848 14903
rect 38194 14900 38200 14952
rect 38252 14940 38258 14952
rect 38657 14943 38715 14949
rect 38657 14940 38669 14943
rect 38252 14912 38669 14940
rect 38252 14900 38258 14912
rect 38657 14909 38669 14912
rect 38703 14909 38715 14943
rect 38657 14903 38715 14909
rect 39758 14832 39764 14884
rect 39816 14872 39822 14884
rect 41386 14872 41414 15048
rect 41782 14968 41788 15020
rect 41840 14968 41846 15020
rect 44376 15017 44404 15048
rect 44105 15011 44163 15017
rect 44105 14977 44117 15011
rect 44151 15008 44163 15011
rect 44361 15011 44419 15017
rect 44151 14980 44312 15008
rect 44151 14977 44163 14980
rect 44105 14971 44163 14977
rect 44284 14940 44312 14980
rect 44361 14977 44373 15011
rect 44407 15008 44419 15011
rect 44744 15008 44772 15107
rect 45554 15104 45560 15116
rect 45612 15104 45618 15156
rect 46750 15104 46756 15156
rect 46808 15104 46814 15156
rect 47949 15147 48007 15153
rect 47949 15113 47961 15147
rect 47995 15144 48007 15147
rect 48406 15144 48412 15156
rect 47995 15116 48412 15144
rect 47995 15113 48007 15116
rect 47949 15107 48007 15113
rect 48406 15104 48412 15116
rect 48464 15104 48470 15156
rect 52638 15144 52644 15156
rect 48516 15116 52644 15144
rect 48516 15076 48544 15116
rect 52638 15104 52644 15116
rect 52696 15104 52702 15156
rect 53190 15104 53196 15156
rect 53248 15104 53254 15156
rect 54573 15147 54631 15153
rect 54573 15113 54585 15147
rect 54619 15144 54631 15147
rect 54754 15144 54760 15156
rect 54619 15116 54760 15144
rect 54619 15113 54631 15116
rect 54573 15107 54631 15113
rect 54754 15104 54760 15116
rect 54812 15104 54818 15156
rect 57146 15104 57152 15156
rect 57204 15144 57210 15156
rect 57517 15147 57575 15153
rect 57517 15144 57529 15147
rect 57204 15116 57529 15144
rect 57204 15104 57210 15116
rect 57517 15113 57529 15116
rect 57563 15113 57575 15147
rect 57517 15107 57575 15113
rect 44407 14980 44772 15008
rect 48148 15048 48544 15076
rect 44407 14977 44419 14980
rect 44361 14971 44419 14977
rect 44634 14940 44640 14952
rect 44284 14912 44640 14940
rect 44634 14900 44640 14912
rect 44692 14900 44698 14952
rect 47397 14943 47455 14949
rect 47397 14909 47409 14943
rect 47443 14909 47455 14943
rect 47397 14903 47455 14909
rect 39816 14844 41414 14872
rect 47412 14872 47440 14903
rect 48038 14900 48044 14952
rect 48096 14900 48102 14952
rect 48148 14949 48176 15048
rect 48682 15036 48688 15088
rect 48740 15036 48746 15088
rect 50890 15036 50896 15088
rect 50948 15076 50954 15088
rect 52457 15079 52515 15085
rect 52457 15076 52469 15079
rect 50948 15048 52469 15076
rect 50948 15036 50954 15048
rect 48133 14943 48191 14949
rect 48133 14909 48145 14943
rect 48179 14909 48191 14943
rect 48700 14940 48728 15036
rect 49418 14968 49424 15020
rect 49476 14968 49482 15020
rect 49510 14968 49516 15020
rect 49568 15017 49574 15020
rect 49568 15011 49617 15017
rect 49568 14977 49571 15011
rect 49605 14977 49617 15011
rect 49568 14971 49617 14977
rect 49568 14968 49574 14971
rect 49694 14968 49700 15020
rect 49752 14968 49758 15020
rect 50614 14968 50620 15020
rect 50672 14968 50678 15020
rect 51833 15011 51891 15017
rect 51833 14977 51845 15011
rect 51879 15008 51891 15011
rect 51994 15008 52000 15020
rect 51879 14980 52000 15008
rect 51879 14977 51891 14980
rect 51833 14971 51891 14977
rect 51994 14968 52000 14980
rect 52052 14968 52058 15020
rect 52104 15017 52132 15048
rect 52457 15045 52469 15048
rect 52503 15076 52515 15079
rect 53208 15076 53236 15104
rect 52503 15048 53236 15076
rect 52503 15045 52515 15048
rect 52457 15039 52515 15045
rect 52932 15017 52960 15048
rect 54110 15036 54116 15088
rect 54168 15036 54174 15088
rect 52089 15011 52147 15017
rect 52089 14977 52101 15011
rect 52135 14977 52147 15011
rect 52089 14971 52147 14977
rect 52917 15011 52975 15017
rect 52917 14977 52929 15011
rect 52963 14977 52975 15011
rect 52917 14971 52975 14977
rect 53184 15011 53242 15017
rect 53184 14977 53196 15011
rect 53230 15008 53242 15011
rect 54128 15008 54156 15036
rect 53230 14980 54156 15008
rect 55217 15011 55275 15017
rect 53230 14977 53242 14980
rect 53184 14971 53242 14977
rect 55217 14977 55229 15011
rect 55263 15008 55275 15011
rect 56226 15008 56232 15020
rect 55263 14980 56232 15008
rect 55263 14977 55275 14980
rect 55217 14971 55275 14977
rect 49970 14940 49976 14952
rect 48700 14912 49976 14940
rect 48133 14903 48191 14909
rect 47581 14875 47639 14881
rect 47581 14872 47593 14875
rect 47412 14844 47593 14872
rect 39816 14832 39822 14844
rect 47581 14841 47593 14844
rect 47627 14841 47639 14875
rect 47581 14835 47639 14841
rect 34388 14776 35848 14804
rect 34388 14764 34394 14776
rect 36538 14764 36544 14816
rect 36596 14804 36602 14816
rect 36633 14807 36691 14813
rect 36633 14804 36645 14807
rect 36596 14776 36645 14804
rect 36596 14764 36602 14776
rect 36633 14773 36645 14776
rect 36679 14773 36691 14807
rect 36633 14767 36691 14773
rect 39298 14764 39304 14816
rect 39356 14764 39362 14816
rect 42150 14764 42156 14816
rect 42208 14764 42214 14816
rect 42981 14807 43039 14813
rect 42981 14773 42993 14807
rect 43027 14804 43039 14807
rect 44726 14804 44732 14816
rect 43027 14776 44732 14804
rect 43027 14773 43039 14776
rect 42981 14767 43039 14773
rect 44726 14764 44732 14776
rect 44784 14764 44790 14816
rect 46566 14764 46572 14816
rect 46624 14804 46630 14816
rect 48148 14804 48176 14903
rect 49970 14900 49976 14912
rect 50028 14900 50034 14952
rect 50433 14943 50491 14949
rect 50433 14909 50445 14943
rect 50479 14909 50491 14943
rect 50433 14903 50491 14909
rect 50448 14872 50476 14903
rect 50709 14875 50767 14881
rect 50709 14872 50721 14875
rect 50448 14844 50721 14872
rect 50709 14841 50721 14844
rect 50755 14872 50767 14875
rect 54297 14875 54355 14881
rect 50755 14844 51074 14872
rect 50755 14841 50767 14844
rect 50709 14835 50767 14841
rect 46624 14776 48176 14804
rect 48777 14807 48835 14813
rect 46624 14764 46630 14776
rect 48777 14773 48789 14807
rect 48823 14804 48835 14807
rect 50798 14804 50804 14816
rect 48823 14776 50804 14804
rect 48823 14773 48835 14776
rect 48777 14767 48835 14773
rect 50798 14764 50804 14776
rect 50856 14764 50862 14816
rect 51046 14804 51074 14844
rect 54297 14841 54309 14875
rect 54343 14872 54355 14875
rect 55232 14872 55260 14971
rect 56226 14968 56232 14980
rect 56284 14968 56290 15020
rect 56404 15011 56462 15017
rect 56404 14977 56416 15011
rect 56450 15008 56462 15011
rect 57885 15011 57943 15017
rect 57885 15008 57897 15011
rect 56450 14980 57897 15008
rect 56450 14977 56462 14980
rect 56404 14971 56462 14977
rect 57885 14977 57897 14980
rect 57931 14977 57943 15011
rect 57885 14971 57943 14977
rect 57974 14968 57980 15020
rect 58032 15008 58038 15020
rect 58437 15011 58495 15017
rect 58437 15008 58449 15011
rect 58032 14980 58449 15008
rect 58032 14968 58038 14980
rect 58437 14977 58449 14980
rect 58483 14977 58495 15011
rect 58437 14971 58495 14977
rect 56137 14943 56195 14949
rect 56137 14909 56149 14943
rect 56183 14909 56195 14943
rect 56137 14903 56195 14909
rect 54343 14844 55260 14872
rect 54343 14841 54355 14844
rect 54297 14835 54355 14841
rect 56152 14816 56180 14903
rect 52086 14804 52092 14816
rect 51046 14776 52092 14804
rect 52086 14764 52092 14776
rect 52144 14764 52150 14816
rect 55214 14764 55220 14816
rect 55272 14804 55278 14816
rect 55493 14807 55551 14813
rect 55493 14804 55505 14807
rect 55272 14776 55505 14804
rect 55272 14764 55278 14776
rect 55493 14773 55505 14776
rect 55539 14773 55551 14807
rect 55493 14767 55551 14773
rect 56045 14807 56103 14813
rect 56045 14773 56057 14807
rect 56091 14804 56103 14807
rect 56134 14804 56140 14816
rect 56091 14776 56140 14804
rect 56091 14773 56103 14776
rect 56045 14767 56103 14773
rect 56134 14764 56140 14776
rect 56192 14764 56198 14816
rect 1104 14714 58880 14736
rect 1104 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 22616 14714
rect 22668 14662 22680 14714
rect 22732 14662 22744 14714
rect 22796 14662 22808 14714
rect 22860 14662 22872 14714
rect 22924 14662 37060 14714
rect 37112 14662 37124 14714
rect 37176 14662 37188 14714
rect 37240 14662 37252 14714
rect 37304 14662 37316 14714
rect 37368 14662 51504 14714
rect 51556 14662 51568 14714
rect 51620 14662 51632 14714
rect 51684 14662 51696 14714
rect 51748 14662 51760 14714
rect 51812 14662 58880 14714
rect 1104 14640 58880 14662
rect 4065 14603 4123 14609
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4154 14600 4160 14612
rect 4111 14572 4160 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 6546 14600 6552 14612
rect 4479 14572 6552 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 8662 14600 8668 14612
rect 7055 14572 8668 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 8662 14560 8668 14572
rect 8720 14600 8726 14612
rect 9582 14600 9588 14612
rect 8720 14572 9588 14600
rect 8720 14560 8726 14572
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12342 14600 12348 14612
rect 11839 14572 12348 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 12342 14560 12348 14572
rect 12400 14600 12406 14612
rect 13170 14600 13176 14612
rect 12400 14572 13176 14600
rect 12400 14560 12406 14572
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13909 14603 13967 14609
rect 13909 14569 13921 14603
rect 13955 14600 13967 14603
rect 14182 14600 14188 14612
rect 13955 14572 14188 14600
rect 13955 14569 13967 14572
rect 13909 14563 13967 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20993 14603 21051 14609
rect 20036 14572 20668 14600
rect 20036 14560 20042 14572
rect 3513 14535 3571 14541
rect 3513 14501 3525 14535
rect 3559 14501 3571 14535
rect 3513 14495 3571 14501
rect 5629 14535 5687 14541
rect 5629 14501 5641 14535
rect 5675 14532 5687 14535
rect 6178 14532 6184 14544
rect 5675 14504 6184 14532
rect 5675 14501 5687 14504
rect 5629 14495 5687 14501
rect 3528 14464 3556 14495
rect 6178 14492 6184 14504
rect 6236 14492 6242 14544
rect 12250 14492 12256 14544
rect 12308 14492 12314 14544
rect 4338 14464 4344 14476
rect 3528 14436 4344 14464
rect 4338 14424 4344 14436
rect 4396 14464 4402 14476
rect 5215 14467 5273 14473
rect 5215 14464 5227 14467
rect 4396 14436 5227 14464
rect 4396 14424 4402 14436
rect 5215 14433 5227 14436
rect 5261 14433 5273 14467
rect 5215 14427 5273 14433
rect 5350 14424 5356 14476
rect 5408 14424 5414 14476
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6638 14464 6644 14476
rect 6319 14436 6644 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9858 14464 9864 14476
rect 8619 14436 9864 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 12268 14464 12296 14492
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12268 14436 12357 14464
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14433 20499 14467
rect 20441 14427 20499 14433
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 2400 14399 2458 14405
rect 2400 14365 2412 14399
rect 2446 14396 2458 14399
rect 2682 14396 2688 14408
rect 2446 14368 2688 14396
rect 2446 14365 2458 14368
rect 2400 14359 2458 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 5074 14356 5080 14408
rect 5132 14356 5138 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 2148 14328 2176 14356
rect 6104 14328 6132 14359
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8306 14399 8364 14405
rect 8306 14396 8318 14399
rect 8076 14368 8318 14396
rect 8076 14356 8082 14368
rect 8306 14365 8318 14368
rect 8352 14365 8364 14399
rect 8306 14359 8364 14365
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9508 14328 9536 14359
rect 10594 14356 10600 14408
rect 10652 14356 10658 14408
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13538 14396 13544 14408
rect 13044 14368 13544 14396
rect 13044 14356 13050 14368
rect 13538 14356 13544 14368
rect 13596 14396 13602 14408
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 13596 14368 14197 14396
rect 13596 14356 13602 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 17218 14356 17224 14408
rect 17276 14396 17282 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17276 14368 17509 14396
rect 17276 14356 17282 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 18322 14356 18328 14408
rect 18380 14356 18386 14408
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20456 14396 20484 14427
rect 20640 14405 20668 14572
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 22370 14600 22376 14612
rect 21039 14572 22376 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 31389 14603 31447 14609
rect 31389 14569 31401 14603
rect 31435 14600 31447 14603
rect 32306 14600 32312 14612
rect 31435 14572 32312 14600
rect 31435 14569 31447 14572
rect 31389 14563 31447 14569
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 32398 14560 32404 14612
rect 32456 14560 32462 14612
rect 38194 14560 38200 14612
rect 38252 14560 38258 14612
rect 39758 14560 39764 14612
rect 39816 14560 39822 14612
rect 51994 14560 52000 14612
rect 52052 14600 52058 14612
rect 52273 14603 52331 14609
rect 52273 14600 52285 14603
rect 52052 14572 52285 14600
rect 52052 14560 52058 14572
rect 52273 14569 52285 14572
rect 52319 14569 52331 14603
rect 52273 14563 52331 14569
rect 54205 14603 54263 14609
rect 54205 14569 54217 14603
rect 54251 14600 54263 14603
rect 54294 14600 54300 14612
rect 54251 14572 54300 14600
rect 54251 14569 54263 14572
rect 54205 14563 54263 14569
rect 54294 14560 54300 14572
rect 54352 14600 54358 14612
rect 54846 14600 54852 14612
rect 54352 14572 54852 14600
rect 54352 14560 54358 14572
rect 54846 14560 54852 14572
rect 54904 14560 54910 14612
rect 31941 14535 31999 14541
rect 31941 14501 31953 14535
rect 31987 14532 31999 14535
rect 32416 14532 32444 14560
rect 31987 14504 32444 14532
rect 31987 14501 31999 14504
rect 31941 14495 31999 14501
rect 39577 14467 39635 14473
rect 39577 14433 39589 14467
rect 39623 14464 39635 14467
rect 39776 14464 39804 14560
rect 48501 14535 48559 14541
rect 48501 14501 48513 14535
rect 48547 14532 48559 14535
rect 49418 14532 49424 14544
rect 48547 14504 49424 14532
rect 48547 14501 48559 14504
rect 48501 14495 48559 14501
rect 49418 14492 49424 14504
rect 49476 14492 49482 14544
rect 50522 14492 50528 14544
rect 50580 14532 50586 14544
rect 51445 14535 51503 14541
rect 50580 14504 50844 14532
rect 50580 14492 50586 14504
rect 50816 14473 50844 14504
rect 51445 14501 51457 14535
rect 51491 14532 51503 14535
rect 57241 14535 57299 14541
rect 51491 14504 52868 14532
rect 51491 14501 51503 14504
rect 51445 14495 51503 14501
rect 39623 14436 39804 14464
rect 50801 14467 50859 14473
rect 39623 14433 39635 14436
rect 39577 14427 39635 14433
rect 50801 14433 50813 14467
rect 50847 14433 50859 14467
rect 50801 14427 50859 14433
rect 20211 14368 20484 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 2148 14300 2544 14328
rect 6104 14300 9536 14328
rect 16853 14331 16911 14337
rect 2516 14272 2544 14300
rect 2498 14220 2504 14272
rect 2556 14220 2562 14272
rect 6270 14220 6276 14272
rect 6328 14260 6334 14272
rect 6546 14260 6552 14272
rect 6328 14232 6552 14260
rect 6328 14220 6334 14232
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7208 14269 7236 14300
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 20456 14328 20484 14368
rect 20625 14399 20683 14405
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 20772 14368 21649 14396
rect 20772 14356 20778 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 25406 14356 25412 14408
rect 25464 14356 25470 14408
rect 26237 14399 26295 14405
rect 26237 14365 26249 14399
rect 26283 14396 26295 14399
rect 26786 14396 26792 14408
rect 26283 14368 26792 14396
rect 26283 14365 26295 14368
rect 26237 14359 26295 14365
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 30834 14356 30840 14408
rect 30892 14356 30898 14408
rect 34330 14356 34336 14408
rect 34388 14356 34394 14408
rect 34974 14356 34980 14408
rect 35032 14396 35038 14408
rect 35253 14399 35311 14405
rect 35253 14396 35265 14399
rect 35032 14368 35265 14396
rect 35032 14356 35038 14368
rect 35253 14365 35265 14368
rect 35299 14365 35311 14399
rect 35253 14359 35311 14365
rect 38105 14399 38163 14405
rect 38105 14365 38117 14399
rect 38151 14396 38163 14399
rect 38562 14396 38568 14408
rect 38151 14368 38568 14396
rect 38151 14365 38163 14368
rect 38105 14359 38163 14365
rect 38562 14356 38568 14368
rect 38620 14356 38626 14408
rect 40402 14356 40408 14408
rect 40460 14356 40466 14408
rect 43070 14356 43076 14408
rect 43128 14356 43134 14408
rect 44085 14399 44143 14405
rect 44085 14365 44097 14399
rect 44131 14396 44143 14399
rect 44910 14396 44916 14408
rect 44131 14368 44916 14396
rect 44131 14365 44143 14368
rect 44085 14359 44143 14365
rect 44910 14356 44916 14368
rect 44968 14356 44974 14408
rect 49142 14356 49148 14408
rect 49200 14356 49206 14408
rect 50816 14396 50844 14427
rect 52086 14424 52092 14476
rect 52144 14424 52150 14476
rect 52840 14473 52868 14504
rect 57241 14501 57253 14535
rect 57287 14532 57299 14535
rect 57287 14504 57928 14532
rect 57287 14501 57299 14504
rect 57241 14495 57299 14501
rect 57900 14473 57928 14504
rect 52825 14467 52883 14473
rect 52825 14433 52837 14467
rect 52871 14433 52883 14467
rect 56597 14467 56655 14473
rect 56597 14464 56609 14467
rect 52825 14427 52883 14433
rect 56336 14436 56609 14464
rect 50816 14368 53604 14396
rect 22480 14328 22508 14356
rect 16899 14300 17632 14328
rect 20456 14300 22508 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17604 14272 17632 14300
rect 24026 14288 24032 14340
rect 24084 14328 24090 14340
rect 24673 14331 24731 14337
rect 24673 14328 24685 14331
rect 24084 14300 24685 14328
rect 24084 14288 24090 14300
rect 24673 14297 24685 14300
rect 24719 14328 24731 14331
rect 24719 14300 26096 14328
rect 24719 14297 24731 14300
rect 24673 14291 24731 14297
rect 26068 14272 26096 14300
rect 30190 14288 30196 14340
rect 30248 14328 30254 14340
rect 31110 14328 31116 14340
rect 30248 14300 31116 14328
rect 30248 14288 30254 14300
rect 31110 14288 31116 14300
rect 31168 14328 31174 14340
rect 37093 14331 37151 14337
rect 37093 14328 37105 14331
rect 31168 14300 37105 14328
rect 31168 14288 31174 14300
rect 37093 14297 37105 14300
rect 37139 14328 37151 14331
rect 37826 14328 37832 14340
rect 37139 14300 37832 14328
rect 37139 14297 37151 14300
rect 37093 14291 37151 14297
rect 37826 14288 37832 14300
rect 37884 14288 37890 14340
rect 39332 14331 39390 14337
rect 39332 14297 39344 14331
rect 39378 14328 39390 14331
rect 39853 14331 39911 14337
rect 39853 14328 39865 14331
rect 39378 14300 39865 14328
rect 39378 14297 39390 14300
rect 39332 14291 39390 14297
rect 39853 14297 39865 14300
rect 39899 14297 39911 14331
rect 39853 14291 39911 14297
rect 47946 14288 47952 14340
rect 48004 14328 48010 14340
rect 48593 14331 48651 14337
rect 48593 14328 48605 14331
rect 48004 14300 48605 14328
rect 48004 14288 48010 14300
rect 48593 14297 48605 14300
rect 48639 14297 48651 14331
rect 48593 14291 48651 14297
rect 49605 14331 49663 14337
rect 49605 14297 49617 14331
rect 49651 14328 49663 14331
rect 50890 14328 50896 14340
rect 49651 14300 50896 14328
rect 49651 14297 49663 14300
rect 49605 14291 49663 14297
rect 50890 14288 50896 14300
rect 50948 14288 50954 14340
rect 51077 14331 51135 14337
rect 51077 14297 51089 14331
rect 51123 14328 51135 14331
rect 51537 14331 51595 14337
rect 51537 14328 51549 14331
rect 51123 14300 51549 14328
rect 51123 14297 51135 14300
rect 51077 14291 51135 14297
rect 51537 14297 51549 14300
rect 51583 14297 51595 14331
rect 53576 14328 53604 14368
rect 53650 14356 53656 14408
rect 53708 14356 53714 14408
rect 56336 14337 56364 14436
rect 56597 14433 56609 14436
rect 56643 14433 56655 14467
rect 56597 14427 56655 14433
rect 57885 14467 57943 14473
rect 57885 14433 57897 14467
rect 57931 14433 57943 14467
rect 57885 14427 57943 14433
rect 56321 14331 56379 14337
rect 56321 14328 56333 14331
rect 53576 14300 56333 14328
rect 51537 14291 51595 14297
rect 56321 14297 56333 14300
rect 56367 14297 56379 14331
rect 56321 14291 56379 14297
rect 56873 14331 56931 14337
rect 56873 14297 56885 14331
rect 56919 14328 56931 14331
rect 57882 14328 57888 14340
rect 56919 14300 57888 14328
rect 56919 14297 56931 14300
rect 56873 14291 56931 14297
rect 57882 14288 57888 14300
rect 57940 14288 57946 14340
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 8938 14220 8944 14272
rect 8996 14220 9002 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10045 14263 10103 14269
rect 10045 14260 10057 14263
rect 9916 14232 10057 14260
rect 9916 14220 9922 14232
rect 10045 14229 10057 14232
rect 10091 14229 10103 14263
rect 10045 14223 10103 14229
rect 14829 14263 14887 14269
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 15286 14260 15292 14272
rect 14875 14232 15292 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 16942 14220 16948 14272
rect 17000 14220 17006 14272
rect 17586 14220 17592 14272
rect 17644 14220 17650 14272
rect 17770 14220 17776 14272
rect 17828 14220 17834 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 20533 14263 20591 14269
rect 20533 14260 20545 14263
rect 18472 14232 20545 14260
rect 18472 14220 18478 14232
rect 20533 14229 20545 14232
rect 20579 14260 20591 14263
rect 20990 14260 20996 14272
rect 20579 14232 20996 14260
rect 20579 14229 20591 14232
rect 20533 14223 20591 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21082 14220 21088 14272
rect 21140 14220 21146 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 25590 14220 25596 14272
rect 25648 14220 25654 14272
rect 26050 14220 26056 14272
rect 26108 14260 26114 14272
rect 26881 14263 26939 14269
rect 26881 14260 26893 14263
rect 26108 14232 26893 14260
rect 26108 14220 26114 14232
rect 26881 14229 26893 14232
rect 26927 14260 26939 14263
rect 29730 14260 29736 14272
rect 26927 14232 29736 14260
rect 26927 14229 26939 14232
rect 26881 14223 26939 14229
rect 29730 14220 29736 14232
rect 29788 14220 29794 14272
rect 30282 14220 30288 14272
rect 30340 14220 30346 14272
rect 32214 14220 32220 14272
rect 32272 14220 32278 14272
rect 32858 14220 32864 14272
rect 32916 14260 32922 14272
rect 33137 14263 33195 14269
rect 33137 14260 33149 14263
rect 32916 14232 33149 14260
rect 32916 14220 32922 14232
rect 33137 14229 33149 14232
rect 33183 14229 33195 14263
rect 33137 14223 33195 14229
rect 33778 14220 33784 14272
rect 33836 14220 33842 14272
rect 34698 14220 34704 14272
rect 34756 14220 34762 14272
rect 37458 14220 37464 14272
rect 37516 14220 37522 14272
rect 42518 14220 42524 14272
rect 42576 14220 42582 14272
rect 43441 14263 43499 14269
rect 43441 14229 43453 14263
rect 43487 14260 43499 14263
rect 43806 14260 43812 14272
rect 43487 14232 43812 14260
rect 43487 14229 43499 14232
rect 43441 14223 43499 14229
rect 43806 14220 43812 14232
rect 43864 14220 43870 14272
rect 44545 14263 44603 14269
rect 44545 14229 44557 14263
rect 44591 14260 44603 14263
rect 44634 14260 44640 14272
rect 44591 14232 44640 14260
rect 44591 14229 44603 14232
rect 44545 14223 44603 14229
rect 44634 14220 44640 14232
rect 44692 14220 44698 14272
rect 47026 14220 47032 14272
rect 47084 14260 47090 14272
rect 47397 14263 47455 14269
rect 47397 14260 47409 14263
rect 47084 14232 47409 14260
rect 47084 14220 47090 14232
rect 47397 14229 47409 14232
rect 47443 14229 47455 14263
rect 47397 14223 47455 14229
rect 50522 14220 50528 14272
rect 50580 14260 50586 14272
rect 50985 14263 51043 14269
rect 50985 14260 50997 14263
rect 50580 14232 50997 14260
rect 50580 14220 50586 14232
rect 50985 14229 50997 14232
rect 51031 14229 51043 14263
rect 50985 14223 51043 14229
rect 53006 14220 53012 14272
rect 53064 14260 53070 14272
rect 53101 14263 53159 14269
rect 53101 14260 53113 14263
rect 53064 14232 53113 14260
rect 53064 14220 53070 14232
rect 53101 14229 53113 14232
rect 53147 14229 53159 14263
rect 53101 14223 53159 14229
rect 56778 14220 56784 14272
rect 56836 14220 56842 14272
rect 57330 14220 57336 14272
rect 57388 14220 57394 14272
rect 1104 14170 59040 14192
rect 1104 14118 15394 14170
rect 15446 14118 15458 14170
rect 15510 14118 15522 14170
rect 15574 14118 15586 14170
rect 15638 14118 15650 14170
rect 15702 14118 29838 14170
rect 29890 14118 29902 14170
rect 29954 14118 29966 14170
rect 30018 14118 30030 14170
rect 30082 14118 30094 14170
rect 30146 14118 44282 14170
rect 44334 14118 44346 14170
rect 44398 14118 44410 14170
rect 44462 14118 44474 14170
rect 44526 14118 44538 14170
rect 44590 14118 58726 14170
rect 58778 14118 58790 14170
rect 58842 14118 58854 14170
rect 58906 14118 58918 14170
rect 58970 14118 58982 14170
rect 59034 14118 59040 14170
rect 1104 14096 59040 14118
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 2924 14028 3617 14056
rect 2924 14016 2930 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 3786 14016 3792 14068
rect 3844 14056 3850 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 3844 14028 4077 14056
rect 3844 14016 3850 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 4065 14019 4123 14025
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14056 6239 14059
rect 6638 14056 6644 14068
rect 6227 14028 6644 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8938 14056 8944 14068
rect 8067 14028 8944 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9122 14016 9128 14068
rect 9180 14016 9186 14068
rect 10229 14059 10287 14065
rect 10229 14025 10241 14059
rect 10275 14056 10287 14059
rect 10594 14056 10600 14068
rect 10275 14028 10600 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12710 14056 12716 14068
rect 12584 14028 12716 14056
rect 12584 14016 12590 14028
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 12986 14016 12992 14068
rect 13044 14016 13050 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 16945 14059 17003 14065
rect 13780 14028 16528 14056
rect 13780 14016 13786 14028
rect 2498 13988 2504 14000
rect 2056 13960 2504 13988
rect 2056 13932 2084 13960
rect 2498 13948 2504 13960
rect 2556 13988 2562 14000
rect 5068 13991 5126 13997
rect 2556 13960 4844 13988
rect 2556 13948 2562 13960
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 2096 13892 2145 13920
rect 2096 13880 2102 13892
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 2133 13883 2191 13889
rect 2222 13880 2228 13932
rect 2280 13920 2286 13932
rect 2389 13923 2447 13929
rect 2389 13920 2401 13923
rect 2280 13892 2401 13920
rect 2280 13880 2286 13892
rect 2389 13889 2401 13892
rect 2435 13889 2447 13923
rect 2389 13883 2447 13889
rect 3970 13880 3976 13932
rect 4028 13880 4034 13932
rect 4816 13929 4844 13960
rect 5068 13957 5080 13991
rect 5114 13988 5126 13991
rect 5258 13988 5264 14000
rect 5114 13960 5264 13988
rect 5114 13957 5126 13960
rect 5068 13951 5126 13957
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13889 4859 13923
rect 5828 13920 5856 14016
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 8757 13991 8815 13997
rect 8757 13957 8769 13991
rect 8803 13988 8815 13991
rect 9140 13988 9168 14016
rect 9490 13988 9496 14000
rect 8803 13960 9496 13988
rect 8803 13957 8815 13960
rect 8757 13951 8815 13957
rect 6730 13920 6736 13932
rect 5828 13892 6736 13920
rect 4801 13883 4859 13889
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 7926 13920 7932 13932
rect 6788 13892 7932 13920
rect 6788 13880 6794 13892
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4706 13852 4712 13864
rect 4295 13824 4712 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 8588 13852 8616 13948
rect 7837 13815 7895 13821
rect 8404 13824 8616 13852
rect 3510 13744 3516 13796
rect 3568 13744 3574 13796
rect 7852 13784 7880 13815
rect 8404 13793 8432 13824
rect 8389 13787 8447 13793
rect 7852 13756 7972 13784
rect 7944 13716 7972 13756
rect 8389 13753 8401 13787
rect 8435 13753 8447 13787
rect 8389 13747 8447 13753
rect 8772 13716 8800 13951
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 11900 13988 11928 14016
rect 10612 13960 11928 13988
rect 14124 13991 14182 13997
rect 10612 13929 10640 13960
rect 14124 13957 14136 13991
rect 14170 13988 14182 13991
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 14170 13960 14565 13988
rect 14170 13957 14182 13960
rect 14124 13951 14182 13957
rect 14553 13957 14565 13960
rect 14599 13957 14611 13991
rect 14553 13951 14611 13957
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 10735 13892 11529 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 14918 13920 14924 13932
rect 11517 13883 11575 13889
rect 14384 13892 14924 13920
rect 14384 13864 14412 13892
rect 14918 13880 14924 13892
rect 14976 13920 14982 13932
rect 15470 13920 15476 13932
rect 14976 13892 15476 13920
rect 14976 13880 14982 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13852 10195 13855
rect 10778 13852 10784 13864
rect 10183 13824 10784 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 10778 13812 10784 13824
rect 10836 13852 10842 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10836 13824 10885 13852
rect 10836 13812 10842 13824
rect 10873 13821 10885 13824
rect 10919 13852 10931 13855
rect 11054 13852 11060 13864
rect 10919 13824 11060 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 12066 13852 12072 13864
rect 11204 13824 12072 13852
rect 11204 13812 11210 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 14366 13812 14372 13864
rect 14424 13812 14430 13864
rect 15194 13812 15200 13864
rect 15252 13812 15258 13864
rect 16500 13861 16528 14028
rect 16945 14025 16957 14059
rect 16991 14056 17003 14059
rect 17218 14056 17224 14068
rect 16991 14028 17224 14056
rect 16991 14025 17003 14028
rect 16945 14019 17003 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17313 14059 17371 14065
rect 17313 14025 17325 14059
rect 17359 14056 17371 14059
rect 17770 14056 17776 14068
rect 17359 14028 17776 14056
rect 17359 14025 17371 14028
rect 17313 14019 17371 14025
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 20070 14016 20076 14068
rect 20128 14016 20134 14068
rect 20257 14059 20315 14065
rect 20257 14025 20269 14059
rect 20303 14056 20315 14059
rect 20622 14056 20628 14068
rect 20303 14028 20628 14056
rect 20303 14025 20315 14028
rect 20257 14019 20315 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 22278 14016 22284 14068
rect 22336 14016 22342 14068
rect 24854 14016 24860 14068
rect 24912 14016 24918 14068
rect 25317 14059 25375 14065
rect 25317 14025 25329 14059
rect 25363 14025 25375 14059
rect 25317 14019 25375 14025
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 18432 13920 18460 14016
rect 20088 13988 20116 14016
rect 22296 13988 22324 14016
rect 24204 13991 24262 13997
rect 20088 13960 21956 13988
rect 22296 13960 24164 13988
rect 17451 13892 18460 13920
rect 21381 13923 21439 13929
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 21381 13889 21393 13923
rect 21427 13920 21439 13923
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21427 13892 21833 13920
rect 21427 13889 21439 13892
rect 21381 13883 21439 13889
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 16500 13784 16528 13815
rect 17586 13812 17592 13864
rect 17644 13812 17650 13864
rect 18598 13812 18604 13864
rect 18656 13852 18662 13864
rect 19242 13852 19248 13864
rect 18656 13824 19248 13852
rect 18656 13812 18662 13824
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19426 13852 19432 13864
rect 19383 13824 19432 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13852 21695 13855
rect 21928 13852 21956 13960
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13920 23995 13923
rect 24026 13920 24032 13932
rect 23983 13892 24032 13920
rect 23983 13889 23995 13892
rect 23937 13883 23995 13889
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 24136 13920 24164 13960
rect 24204 13957 24216 13991
rect 24250 13988 24262 13991
rect 24872 13988 24900 14016
rect 24250 13960 24900 13988
rect 25332 13988 25360 14019
rect 25406 14016 25412 14068
rect 25464 14016 25470 14068
rect 25590 14016 25596 14068
rect 25648 14056 25654 14068
rect 25869 14059 25927 14065
rect 25869 14056 25881 14059
rect 25648 14028 25881 14056
rect 25648 14016 25654 14028
rect 25869 14025 25881 14028
rect 25915 14025 25927 14059
rect 25869 14019 25927 14025
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 27709 14059 27767 14065
rect 27709 14056 27721 14059
rect 26660 14028 27721 14056
rect 26660 14016 26666 14028
rect 27709 14025 27721 14028
rect 27755 14025 27767 14059
rect 27709 14019 27767 14025
rect 28077 14059 28135 14065
rect 28077 14025 28089 14059
rect 28123 14056 28135 14059
rect 28350 14056 28356 14068
rect 28123 14028 28356 14056
rect 28123 14025 28135 14028
rect 28077 14019 28135 14025
rect 28350 14016 28356 14028
rect 28408 14016 28414 14068
rect 30009 14059 30067 14065
rect 30009 14025 30021 14059
rect 30055 14056 30067 14059
rect 30190 14056 30196 14068
rect 30055 14028 30196 14056
rect 30055 14025 30067 14028
rect 30009 14019 30067 14025
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 30469 14059 30527 14065
rect 30469 14025 30481 14059
rect 30515 14056 30527 14059
rect 30834 14056 30840 14068
rect 30515 14028 30840 14056
rect 30515 14025 30527 14028
rect 30469 14019 30527 14025
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 30926 14016 30932 14068
rect 30984 14016 30990 14068
rect 33962 14016 33968 14068
rect 34020 14056 34026 14068
rect 34425 14059 34483 14065
rect 34425 14056 34437 14059
rect 34020 14028 34437 14056
rect 34020 14016 34026 14028
rect 34425 14025 34437 14028
rect 34471 14025 34483 14059
rect 34425 14019 34483 14025
rect 34532 14028 34928 14056
rect 34532 13988 34560 14028
rect 34793 13991 34851 13997
rect 34793 13988 34805 13991
rect 25332 13960 26832 13988
rect 24250 13957 24262 13960
rect 24204 13951 24262 13957
rect 26804 13932 26832 13960
rect 28966 13960 34560 13988
rect 34624 13960 34805 13988
rect 24136 13892 24992 13920
rect 21683 13824 22094 13852
rect 21683 13821 21695 13824
rect 21637 13815 21695 13821
rect 18230 13784 18236 13796
rect 16500 13756 18236 13784
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 22066 13728 22094 13824
rect 22370 13812 22376 13864
rect 22428 13812 22434 13864
rect 24964 13852 24992 13892
rect 25774 13880 25780 13932
rect 25832 13880 25838 13932
rect 25884 13892 26096 13920
rect 25884 13852 25912 13892
rect 24964 13824 25912 13852
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13821 26019 13855
rect 26068 13852 26096 13892
rect 26786 13880 26792 13932
rect 26844 13880 26850 13932
rect 28966 13920 28994 13960
rect 27724 13892 28994 13920
rect 30837 13923 30895 13929
rect 27157 13855 27215 13861
rect 27157 13852 27169 13855
rect 26068 13824 27169 13852
rect 25961 13815 26019 13821
rect 27157 13821 27169 13824
rect 27203 13852 27215 13855
rect 27433 13855 27491 13861
rect 27433 13852 27445 13855
rect 27203 13824 27445 13852
rect 27203 13821 27215 13824
rect 27157 13815 27215 13821
rect 27433 13821 27445 13824
rect 27479 13821 27491 13855
rect 27433 13815 27491 13821
rect 25222 13744 25228 13796
rect 25280 13784 25286 13796
rect 25976 13784 26004 13815
rect 27522 13812 27528 13864
rect 27580 13852 27586 13864
rect 27617 13855 27675 13861
rect 27617 13852 27629 13855
rect 27580 13824 27629 13852
rect 27580 13812 27586 13824
rect 27617 13821 27629 13824
rect 27663 13821 27675 13855
rect 27617 13815 27675 13821
rect 26513 13787 26571 13793
rect 26513 13784 26525 13787
rect 25280 13756 26525 13784
rect 25280 13744 25286 13756
rect 26513 13753 26525 13756
rect 26559 13784 26571 13787
rect 27724 13784 27752 13892
rect 30837 13889 30849 13923
rect 30883 13920 30895 13923
rect 31297 13923 31355 13929
rect 31297 13920 31309 13923
rect 30883 13892 31309 13920
rect 30883 13889 30895 13892
rect 30837 13883 30895 13889
rect 31297 13889 31309 13892
rect 31343 13889 31355 13923
rect 32858 13920 32864 13932
rect 31297 13883 31355 13889
rect 32324 13892 32864 13920
rect 32324 13864 32352 13892
rect 32858 13880 32864 13892
rect 32916 13920 32922 13932
rect 33220 13923 33278 13929
rect 32916 13892 32996 13920
rect 32916 13880 32922 13892
rect 27798 13812 27804 13864
rect 27856 13852 27862 13864
rect 28721 13855 28779 13861
rect 28721 13852 28733 13855
rect 27856 13824 28733 13852
rect 27856 13812 27862 13824
rect 28721 13821 28733 13824
rect 28767 13821 28779 13855
rect 28721 13815 28779 13821
rect 31110 13812 31116 13864
rect 31168 13812 31174 13864
rect 31202 13812 31208 13864
rect 31260 13852 31266 13864
rect 31849 13855 31907 13861
rect 31849 13852 31861 13855
rect 31260 13824 31861 13852
rect 31260 13812 31266 13824
rect 31849 13821 31861 13824
rect 31895 13821 31907 13855
rect 31849 13815 31907 13821
rect 26559 13756 27752 13784
rect 31864 13784 31892 13815
rect 32306 13812 32312 13864
rect 32364 13812 32370 13864
rect 32674 13812 32680 13864
rect 32732 13812 32738 13864
rect 32968 13861 32996 13892
rect 33220 13889 33232 13923
rect 33266 13920 33278 13923
rect 33778 13920 33784 13932
rect 33266 13892 33784 13920
rect 33266 13889 33278 13892
rect 33220 13883 33278 13889
rect 33778 13880 33784 13892
rect 33836 13880 33842 13932
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 34624 13920 34652 13960
rect 34793 13957 34805 13960
rect 34839 13957 34851 13991
rect 34900 13988 34928 14028
rect 37458 14016 37464 14068
rect 37516 14056 37522 14068
rect 37645 14059 37703 14065
rect 37645 14056 37657 14059
rect 37516 14028 37657 14056
rect 37516 14016 37522 14028
rect 37645 14025 37657 14028
rect 37691 14025 37703 14059
rect 37645 14019 37703 14025
rect 39025 14059 39083 14065
rect 39025 14025 39037 14059
rect 39071 14056 39083 14059
rect 39298 14056 39304 14068
rect 39071 14028 39304 14056
rect 39071 14025 39083 14028
rect 39025 14019 39083 14025
rect 39298 14016 39304 14028
rect 39356 14016 39362 14068
rect 39485 14059 39543 14065
rect 39485 14025 39497 14059
rect 39531 14056 39543 14059
rect 40402 14056 40408 14068
rect 39531 14028 40408 14056
rect 39531 14025 39543 14028
rect 39485 14019 39543 14025
rect 40402 14016 40408 14028
rect 40460 14016 40466 14068
rect 47946 14016 47952 14068
rect 48004 14016 48010 14068
rect 48317 14059 48375 14065
rect 48317 14025 48329 14059
rect 48363 14025 48375 14059
rect 48317 14019 48375 14025
rect 49421 14059 49479 14065
rect 49421 14025 49433 14059
rect 49467 14056 49479 14059
rect 50614 14056 50620 14068
rect 49467 14028 50620 14056
rect 49467 14025 49479 14028
rect 49421 14019 49479 14025
rect 41598 13988 41604 14000
rect 34900 13960 41604 13988
rect 34793 13951 34851 13957
rect 41598 13948 41604 13960
rect 41656 13948 41662 14000
rect 35805 13923 35863 13929
rect 35805 13920 35817 13923
rect 34204 13892 34652 13920
rect 34716 13892 35817 13920
rect 34204 13880 34210 13892
rect 32953 13855 33011 13861
rect 32953 13821 32965 13855
rect 32999 13821 33011 13855
rect 32953 13815 33011 13821
rect 31864 13756 32996 13784
rect 26559 13753 26571 13756
rect 26513 13747 26571 13753
rect 32968 13728 32996 13756
rect 34238 13744 34244 13796
rect 34296 13784 34302 13796
rect 34333 13787 34391 13793
rect 34333 13784 34345 13787
rect 34296 13756 34345 13784
rect 34296 13744 34302 13756
rect 34333 13753 34345 13756
rect 34379 13784 34391 13787
rect 34716 13784 34744 13892
rect 35805 13889 35817 13892
rect 35851 13889 35863 13923
rect 35805 13883 35863 13889
rect 37734 13880 37740 13932
rect 37792 13920 37798 13932
rect 39117 13923 39175 13929
rect 39117 13920 39129 13923
rect 37792 13892 39129 13920
rect 37792 13880 37798 13892
rect 39117 13889 39129 13892
rect 39163 13889 39175 13923
rect 40494 13920 40500 13932
rect 39117 13883 39175 13889
rect 39500 13892 40500 13920
rect 34790 13812 34796 13864
rect 34848 13852 34854 13864
rect 34885 13855 34943 13861
rect 34885 13852 34897 13855
rect 34848 13824 34897 13852
rect 34848 13812 34854 13824
rect 34885 13821 34897 13824
rect 34931 13821 34943 13855
rect 34885 13815 34943 13821
rect 35023 13855 35081 13861
rect 35023 13821 35035 13855
rect 35069 13852 35081 13855
rect 35342 13852 35348 13864
rect 35069 13824 35348 13852
rect 35069 13821 35081 13824
rect 35023 13815 35081 13821
rect 35342 13812 35348 13824
rect 35400 13812 35406 13864
rect 37093 13855 37151 13861
rect 37093 13821 37105 13855
rect 37139 13852 37151 13855
rect 37139 13824 37320 13852
rect 37139 13821 37151 13824
rect 37093 13815 37151 13821
rect 34379 13756 34744 13784
rect 35360 13784 35388 13812
rect 37292 13793 37320 13824
rect 37826 13812 37832 13864
rect 37884 13812 37890 13864
rect 38838 13812 38844 13864
rect 38896 13852 38902 13864
rect 39500 13852 39528 13892
rect 40494 13880 40500 13892
rect 40552 13880 40558 13932
rect 43248 13923 43306 13929
rect 43248 13889 43260 13923
rect 43294 13920 43306 13923
rect 44453 13923 44511 13929
rect 44453 13920 44465 13923
rect 43294 13892 44465 13920
rect 43294 13889 43306 13892
rect 43248 13883 43306 13889
rect 44453 13889 44465 13892
rect 44499 13889 44511 13923
rect 48332 13920 48360 14019
rect 50614 14016 50620 14028
rect 50672 14056 50678 14068
rect 50672 14028 51074 14056
rect 50672 14016 50678 14028
rect 50890 13948 50896 14000
rect 50948 13948 50954 14000
rect 48961 13923 49019 13929
rect 48961 13920 48973 13923
rect 48332 13892 48973 13920
rect 44453 13883 44511 13889
rect 48961 13889 48973 13892
rect 49007 13889 49019 13923
rect 48961 13883 49019 13889
rect 50545 13923 50603 13929
rect 50545 13889 50557 13923
rect 50591 13920 50603 13923
rect 50801 13923 50859 13929
rect 50591 13892 50752 13920
rect 50591 13889 50603 13892
rect 50545 13883 50603 13889
rect 38896 13824 39528 13852
rect 38896 13812 38902 13824
rect 39574 13812 39580 13864
rect 39632 13812 39638 13864
rect 42610 13812 42616 13864
rect 42668 13852 42674 13864
rect 42981 13855 43039 13861
rect 42981 13852 42993 13855
rect 42668 13824 42993 13852
rect 42668 13812 42674 13824
rect 42981 13821 42993 13824
rect 43027 13821 43039 13855
rect 42981 13815 43039 13821
rect 44266 13812 44272 13864
rect 44324 13852 44330 13864
rect 45005 13855 45063 13861
rect 45005 13852 45017 13855
rect 44324 13824 45017 13852
rect 44324 13812 44330 13824
rect 45005 13821 45017 13824
rect 45051 13821 45063 13855
rect 45005 13815 45063 13821
rect 45278 13812 45284 13864
rect 45336 13852 45342 13864
rect 46566 13852 46572 13864
rect 45336 13824 46572 13852
rect 45336 13812 45342 13824
rect 46566 13812 46572 13824
rect 46624 13812 46630 13864
rect 47394 13812 47400 13864
rect 47452 13812 47458 13864
rect 47765 13855 47823 13861
rect 47765 13821 47777 13855
rect 47811 13821 47823 13855
rect 47765 13815 47823 13821
rect 47857 13855 47915 13861
rect 47857 13821 47869 13855
rect 47903 13852 47915 13855
rect 47946 13852 47952 13864
rect 47903 13824 47952 13852
rect 47903 13821 47915 13824
rect 47857 13815 47915 13821
rect 37277 13787 37335 13793
rect 35360 13756 36584 13784
rect 34379 13753 34391 13756
rect 34333 13747 34391 13753
rect 7944 13688 8800 13716
rect 11330 13676 11336 13728
rect 11388 13676 11394 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 14458 13716 14464 13728
rect 11940 13688 14464 13716
rect 11940 13676 11946 13688
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 17954 13676 17960 13728
rect 18012 13676 18018 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18693 13719 18751 13725
rect 18693 13716 18705 13719
rect 18196 13688 18705 13716
rect 18196 13676 18202 13688
rect 18693 13685 18705 13688
rect 18739 13685 18751 13719
rect 22066 13688 22100 13728
rect 18693 13679 18751 13685
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 28166 13676 28172 13728
rect 28224 13676 28230 13728
rect 29270 13676 29276 13728
rect 29328 13676 29334 13728
rect 30377 13719 30435 13725
rect 30377 13685 30389 13719
rect 30423 13716 30435 13719
rect 31386 13716 31392 13728
rect 30423 13688 31392 13716
rect 30423 13685 30435 13688
rect 30377 13679 30435 13685
rect 31386 13676 31392 13688
rect 31444 13676 31450 13728
rect 32122 13676 32128 13728
rect 32180 13676 32186 13728
rect 32950 13676 32956 13728
rect 33008 13676 33014 13728
rect 35250 13676 35256 13728
rect 35308 13676 35314 13728
rect 36446 13676 36452 13728
rect 36504 13676 36510 13728
rect 36556 13716 36584 13756
rect 37277 13753 37289 13787
rect 37323 13753 37335 13787
rect 37277 13747 37335 13753
rect 38102 13744 38108 13796
rect 38160 13784 38166 13796
rect 38381 13787 38439 13793
rect 38381 13784 38393 13787
rect 38160 13756 38393 13784
rect 38160 13744 38166 13756
rect 38381 13753 38393 13756
rect 38427 13753 38439 13787
rect 38381 13747 38439 13753
rect 38286 13716 38292 13728
rect 36556 13688 38292 13716
rect 38286 13676 38292 13688
rect 38344 13716 38350 13728
rect 39114 13716 39120 13728
rect 38344 13688 39120 13716
rect 38344 13676 38350 13688
rect 39114 13676 39120 13688
rect 39172 13676 39178 13728
rect 40218 13676 40224 13728
rect 40276 13676 40282 13728
rect 42242 13676 42248 13728
rect 42300 13716 42306 13728
rect 43162 13716 43168 13728
rect 42300 13688 43168 13716
rect 42300 13676 42306 13688
rect 43162 13676 43168 13688
rect 43220 13676 43226 13728
rect 44361 13719 44419 13725
rect 44361 13685 44373 13719
rect 44407 13716 44419 13719
rect 44910 13716 44916 13728
rect 44407 13688 44916 13716
rect 44407 13685 44419 13688
rect 44361 13679 44419 13685
rect 44910 13676 44916 13688
rect 44968 13676 44974 13728
rect 46750 13676 46756 13728
rect 46808 13676 46814 13728
rect 47026 13676 47032 13728
rect 47084 13716 47090 13728
rect 47780 13716 47808 13815
rect 47946 13812 47952 13824
rect 48004 13812 48010 13864
rect 50724 13852 50752 13892
rect 50801 13889 50813 13923
rect 50847 13920 50859 13923
rect 50908 13920 50936 13948
rect 50847 13892 50936 13920
rect 51046 13920 51074 14028
rect 52638 14016 52644 14068
rect 52696 14056 52702 14068
rect 53009 14059 53067 14065
rect 53009 14056 53021 14059
rect 52696 14028 53021 14056
rect 52696 14016 52702 14028
rect 53009 14025 53021 14028
rect 53055 14025 53067 14059
rect 53009 14019 53067 14025
rect 53193 14059 53251 14065
rect 53193 14025 53205 14059
rect 53239 14056 53251 14059
rect 53650 14056 53656 14068
rect 53239 14028 53656 14056
rect 53239 14025 53251 14028
rect 53193 14019 53251 14025
rect 52181 13923 52239 13929
rect 52181 13920 52193 13923
rect 51046 13892 52193 13920
rect 50847 13889 50859 13892
rect 50801 13883 50859 13889
rect 52181 13889 52193 13892
rect 52227 13889 52239 13923
rect 52181 13883 52239 13889
rect 50893 13855 50951 13861
rect 50893 13852 50905 13855
rect 50724 13824 50905 13852
rect 50893 13821 50905 13824
rect 50939 13821 50951 13855
rect 50893 13815 50951 13821
rect 51258 13812 51264 13864
rect 51316 13852 51322 13864
rect 51445 13855 51503 13861
rect 51445 13852 51457 13855
rect 51316 13824 51457 13852
rect 51316 13812 51322 13824
rect 51445 13821 51457 13824
rect 51491 13821 51503 13855
rect 51445 13815 51503 13821
rect 53024 13784 53052 14019
rect 53650 14016 53656 14028
rect 53708 14016 53714 14068
rect 57330 14016 57336 14068
rect 57388 14016 57394 14068
rect 57882 14016 57888 14068
rect 57940 14016 57946 14068
rect 56588 13991 56646 13997
rect 56588 13957 56600 13991
rect 56634 13988 56646 13991
rect 57348 13988 57376 14016
rect 56634 13960 57376 13988
rect 56634 13957 56646 13960
rect 56588 13951 56646 13957
rect 53561 13923 53619 13929
rect 53561 13889 53573 13923
rect 53607 13920 53619 13923
rect 54021 13923 54079 13929
rect 54021 13920 54033 13923
rect 53607 13892 54033 13920
rect 53607 13889 53619 13892
rect 53561 13883 53619 13889
rect 54021 13889 54033 13892
rect 54067 13889 54079 13923
rect 54021 13883 54079 13889
rect 53650 13812 53656 13864
rect 53708 13812 53714 13864
rect 53745 13855 53803 13861
rect 53745 13821 53757 13855
rect 53791 13821 53803 13855
rect 53745 13815 53803 13821
rect 54665 13855 54723 13861
rect 54665 13821 54677 13855
rect 54711 13852 54723 13855
rect 54938 13852 54944 13864
rect 54711 13824 54944 13852
rect 54711 13821 54723 13824
rect 54665 13815 54723 13821
rect 53760 13784 53788 13815
rect 54938 13812 54944 13824
rect 54996 13812 55002 13864
rect 55306 13812 55312 13864
rect 55364 13812 55370 13864
rect 56321 13855 56379 13861
rect 56321 13852 56333 13855
rect 56152 13824 56333 13852
rect 53024 13756 53788 13784
rect 56152 13728 56180 13824
rect 56321 13821 56333 13824
rect 56367 13821 56379 13855
rect 58437 13855 58495 13861
rect 58437 13852 58449 13855
rect 56321 13815 56379 13821
rect 57716 13824 58449 13852
rect 57716 13796 57744 13824
rect 58437 13821 58449 13824
rect 58483 13821 58495 13855
rect 58437 13815 58495 13821
rect 57698 13744 57704 13796
rect 57756 13744 57762 13796
rect 47084 13688 47808 13716
rect 47084 13676 47090 13688
rect 48406 13676 48412 13728
rect 48464 13676 48470 13728
rect 51166 13676 51172 13728
rect 51224 13716 51230 13728
rect 51629 13719 51687 13725
rect 51629 13716 51641 13719
rect 51224 13688 51641 13716
rect 51224 13676 51230 13688
rect 51629 13685 51641 13688
rect 51675 13685 51687 13719
rect 51629 13679 51687 13685
rect 54754 13676 54760 13728
rect 54812 13676 54818 13728
rect 56134 13676 56140 13728
rect 56192 13676 56198 13728
rect 56318 13676 56324 13728
rect 56376 13716 56382 13728
rect 57606 13716 57612 13728
rect 56376 13688 57612 13716
rect 56376 13676 56382 13688
rect 57606 13676 57612 13688
rect 57664 13676 57670 13728
rect 1104 13626 58880 13648
rect 1104 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 22616 13626
rect 22668 13574 22680 13626
rect 22732 13574 22744 13626
rect 22796 13574 22808 13626
rect 22860 13574 22872 13626
rect 22924 13574 37060 13626
rect 37112 13574 37124 13626
rect 37176 13574 37188 13626
rect 37240 13574 37252 13626
rect 37304 13574 37316 13626
rect 37368 13574 51504 13626
rect 51556 13574 51568 13626
rect 51620 13574 51632 13626
rect 51684 13574 51696 13626
rect 51748 13574 51760 13626
rect 51812 13574 58880 13626
rect 1104 13552 58880 13574
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 14921 13515 14979 13521
rect 12124 13484 13032 13512
rect 12124 13472 12130 13484
rect 10873 13447 10931 13453
rect 10873 13413 10885 13447
rect 10919 13444 10931 13447
rect 10919 13416 12204 13444
rect 10919 13413 10931 13416
rect 10873 13407 10931 13413
rect 12176 13388 12204 13416
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12667 13379 12725 13385
rect 12667 13376 12679 13379
rect 12216 13348 12679 13376
rect 12216 13336 12222 13348
rect 12667 13345 12679 13348
rect 12713 13345 12725 13379
rect 12667 13339 12725 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 13004 13376 13032 13484
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 15194 13512 15200 13524
rect 14967 13484 15200 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15528 13484 16129 13512
rect 15528 13472 15534 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 16117 13475 16175 13481
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 18598 13512 18604 13524
rect 17727 13484 18604 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 15102 13444 15108 13456
rect 14200 13416 15108 13444
rect 14200 13388 14228 13416
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 12851 13348 13032 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13136 13348 13492 13376
rect 13136 13336 13142 13348
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 11330 13308 11336 13320
rect 9539 13280 11336 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 11900 13308 11928 13336
rect 11471 13280 11928 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 13464 13308 13492 13348
rect 13538 13336 13544 13388
rect 13596 13336 13602 13388
rect 14182 13336 14188 13388
rect 14240 13336 14246 13388
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 14516 13348 15393 13376
rect 14516 13336 14522 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 15565 13379 15623 13385
rect 15565 13345 15577 13379
rect 15611 13376 15623 13379
rect 15746 13376 15752 13388
rect 15611 13348 15752 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16132 13376 16160 13475
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 18690 13472 18696 13524
rect 18748 13512 18754 13524
rect 19061 13515 19119 13521
rect 19061 13512 19073 13515
rect 18748 13484 19073 13512
rect 18748 13472 18754 13484
rect 19061 13481 19073 13484
rect 19107 13512 19119 13515
rect 19334 13512 19340 13524
rect 19107 13484 19340 13512
rect 19107 13481 19119 13484
rect 19061 13475 19119 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19426 13472 19432 13524
rect 19484 13472 19490 13524
rect 21453 13515 21511 13521
rect 21453 13481 21465 13515
rect 21499 13512 21511 13515
rect 22370 13512 22376 13524
rect 21499 13484 22376 13512
rect 21499 13481 21511 13484
rect 21453 13475 21511 13481
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 26050 13512 26056 13524
rect 25547 13484 26056 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 27522 13512 27528 13524
rect 26160 13484 27528 13512
rect 18509 13447 18567 13453
rect 17880 13416 18276 13444
rect 16298 13376 16304 13388
rect 16132 13348 16304 13376
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 17880 13385 17908 13416
rect 18248 13388 18276 13416
rect 18509 13413 18521 13447
rect 18555 13444 18567 13447
rect 19444 13444 19472 13472
rect 22278 13444 22284 13456
rect 18555 13416 19472 13444
rect 20272 13416 22284 13444
rect 18555 13413 18567 13416
rect 18509 13407 18567 13413
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 18012 13348 18061 13376
rect 18012 13336 18018 13348
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 18049 13339 18107 13345
rect 18230 13336 18236 13388
rect 18288 13336 18294 13388
rect 19518 13336 19524 13388
rect 19576 13376 19582 13388
rect 20272 13385 20300 13416
rect 22278 13404 22284 13416
rect 22336 13404 22342 13456
rect 24397 13447 24455 13453
rect 24397 13413 24409 13447
rect 24443 13413 24455 13447
rect 26160 13444 26188 13484
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 27798 13472 27804 13524
rect 27856 13472 27862 13524
rect 31205 13515 31263 13521
rect 31205 13481 31217 13515
rect 31251 13512 31263 13515
rect 32674 13512 32680 13524
rect 31251 13484 32680 13512
rect 31251 13481 31263 13484
rect 31205 13475 31263 13481
rect 32674 13472 32680 13484
rect 32732 13512 32738 13524
rect 34701 13515 34759 13521
rect 32732 13484 33364 13512
rect 32732 13472 32738 13484
rect 24397 13407 24455 13413
rect 25884 13416 26188 13444
rect 20257 13379 20315 13385
rect 20257 13376 20269 13379
rect 19576 13348 20269 13376
rect 19576 13336 19582 13348
rect 20257 13345 20269 13348
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13376 20959 13379
rect 21174 13376 21180 13388
rect 20947 13348 21180 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 24213 13379 24271 13385
rect 24213 13345 24225 13379
rect 24259 13376 24271 13379
rect 24412 13376 24440 13407
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 24259 13348 24440 13376
rect 24504 13348 24961 13376
rect 24259 13345 24271 13348
rect 24213 13339 24271 13345
rect 13725 13311 13783 13317
rect 13464 13280 13584 13308
rect 9760 13243 9818 13249
rect 9760 13209 9772 13243
rect 9806 13240 9818 13243
rect 10410 13240 10416 13252
rect 9806 13212 10416 13240
rect 9806 13209 9818 13212
rect 9760 13203 9818 13209
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 13556 13240 13584 13280
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 14090 13308 14096 13320
rect 13771 13280 14096 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14734 13308 14740 13320
rect 14415 13280 14740 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 16568 13311 16626 13317
rect 16568 13277 16580 13311
rect 16614 13308 16626 13311
rect 18138 13308 18144 13320
rect 16614 13280 18144 13308
rect 16614 13277 16626 13280
rect 16568 13271 16626 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19668 13280 19993 13308
rect 19668 13268 19674 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20162 13268 20168 13320
rect 20220 13308 20226 13320
rect 20990 13308 20996 13320
rect 20220 13280 20996 13308
rect 20220 13268 20226 13280
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 24118 13308 24124 13320
rect 23676 13280 24124 13308
rect 13556 13212 16160 13240
rect 16132 13184 16160 13212
rect 18414 13200 18420 13252
rect 18472 13240 18478 13252
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 18472 13212 20085 13240
rect 18472 13200 18478 13212
rect 20073 13209 20085 13212
rect 20119 13209 20131 13243
rect 20073 13203 20131 13209
rect 23477 13243 23535 13249
rect 23477 13209 23489 13243
rect 23523 13240 23535 13243
rect 23676 13240 23704 13280
rect 24118 13268 24124 13280
rect 24176 13308 24182 13320
rect 24504 13308 24532 13348
rect 24949 13345 24961 13348
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 25774 13336 25780 13388
rect 25832 13336 25838 13388
rect 25884 13385 25912 13416
rect 26970 13404 26976 13456
rect 27028 13444 27034 13456
rect 27065 13447 27123 13453
rect 27065 13444 27077 13447
rect 27028 13416 27077 13444
rect 27028 13404 27034 13416
rect 27065 13413 27077 13416
rect 27111 13413 27123 13447
rect 27065 13407 27123 13413
rect 25869 13379 25927 13385
rect 25869 13345 25881 13379
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 26326 13336 26332 13388
rect 26384 13376 26390 13388
rect 27709 13379 27767 13385
rect 26384 13348 26556 13376
rect 26384 13336 26390 13348
rect 24176 13280 24532 13308
rect 24857 13311 24915 13317
rect 24176 13268 24182 13280
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 25792 13308 25820 13336
rect 26528 13317 26556 13348
rect 27709 13345 27721 13379
rect 27755 13376 27767 13379
rect 27816 13376 27844 13472
rect 27755 13348 27844 13376
rect 27755 13345 27767 13348
rect 27709 13339 27767 13345
rect 31386 13336 31392 13388
rect 31444 13336 31450 13388
rect 31573 13379 31631 13385
rect 31573 13345 31585 13379
rect 31619 13376 31631 13379
rect 32122 13376 32128 13388
rect 31619 13348 32128 13376
rect 31619 13345 31631 13348
rect 31573 13339 31631 13345
rect 32122 13336 32128 13348
rect 32180 13336 32186 13388
rect 32861 13379 32919 13385
rect 32861 13376 32873 13379
rect 32324 13348 32873 13376
rect 24903 13280 25820 13308
rect 26513 13311 26571 13317
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 26513 13277 26525 13311
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 26602 13268 26608 13320
rect 26660 13317 26666 13320
rect 26660 13311 26709 13317
rect 26660 13277 26663 13311
rect 26697 13277 26709 13311
rect 26660 13271 26709 13277
rect 26660 13268 26666 13271
rect 26786 13268 26792 13320
rect 26844 13268 26850 13320
rect 27525 13311 27583 13317
rect 27525 13277 27537 13311
rect 27571 13308 27583 13311
rect 27798 13308 27804 13320
rect 27571 13280 27804 13308
rect 27571 13277 27583 13280
rect 27525 13271 27583 13277
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 29181 13311 29239 13317
rect 29181 13277 29193 13311
rect 29227 13308 29239 13311
rect 29270 13308 29276 13320
rect 29227 13280 29276 13308
rect 29227 13277 29239 13280
rect 29181 13271 29239 13277
rect 29270 13268 29276 13280
rect 29328 13308 29334 13320
rect 29730 13308 29736 13320
rect 29328 13280 29736 13308
rect 29328 13268 29334 13280
rect 29730 13268 29736 13280
rect 29788 13308 29794 13320
rect 29825 13311 29883 13317
rect 29825 13308 29837 13311
rect 29788 13280 29837 13308
rect 29788 13268 29794 13280
rect 29825 13277 29837 13280
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 30926 13268 30932 13320
rect 30984 13308 30990 13320
rect 31478 13308 31484 13320
rect 30984 13280 31484 13308
rect 30984 13268 30990 13280
rect 31478 13268 31484 13280
rect 31536 13308 31542 13320
rect 31665 13311 31723 13317
rect 31665 13308 31677 13311
rect 31536 13280 31677 13308
rect 31536 13268 31542 13280
rect 31665 13277 31677 13280
rect 31711 13277 31723 13311
rect 32324 13308 32352 13348
rect 32861 13345 32873 13348
rect 32907 13345 32919 13379
rect 32861 13339 32919 13345
rect 32950 13336 32956 13388
rect 33008 13385 33014 13388
rect 33008 13379 33057 13385
rect 33008 13345 33011 13379
rect 33045 13345 33057 13379
rect 33008 13339 33057 13345
rect 33137 13379 33195 13385
rect 33137 13345 33149 13379
rect 33183 13376 33195 13379
rect 33336 13376 33364 13484
rect 34701 13481 34713 13515
rect 34747 13512 34759 13515
rect 34974 13512 34980 13524
rect 34747 13484 34980 13512
rect 34747 13481 34759 13484
rect 34701 13475 34759 13481
rect 34974 13472 34980 13484
rect 35032 13472 35038 13524
rect 35342 13472 35348 13524
rect 35400 13472 35406 13524
rect 37461 13515 37519 13521
rect 37461 13481 37473 13515
rect 37507 13512 37519 13515
rect 38286 13512 38292 13524
rect 37507 13484 38292 13512
rect 37507 13481 37519 13484
rect 37461 13475 37519 13481
rect 38286 13472 38292 13484
rect 38344 13512 38350 13524
rect 38746 13512 38752 13524
rect 38344 13484 38752 13512
rect 38344 13472 38350 13484
rect 38746 13472 38752 13484
rect 38804 13472 38810 13524
rect 40494 13472 40500 13524
rect 40552 13512 40558 13524
rect 43349 13515 43407 13521
rect 43349 13512 43361 13515
rect 40552 13484 43361 13512
rect 40552 13472 40558 13484
rect 43349 13481 43361 13484
rect 43395 13481 43407 13515
rect 43349 13475 43407 13481
rect 33413 13447 33471 13453
rect 33413 13413 33425 13447
rect 33459 13444 33471 13447
rect 33502 13444 33508 13456
rect 33459 13416 33508 13444
rect 33459 13413 33471 13416
rect 33413 13407 33471 13413
rect 33502 13404 33508 13416
rect 33560 13404 33566 13456
rect 33594 13404 33600 13456
rect 33652 13444 33658 13456
rect 34333 13447 34391 13453
rect 34333 13444 34345 13447
rect 33652 13416 34345 13444
rect 33652 13404 33658 13416
rect 34333 13413 34345 13416
rect 34379 13444 34391 13447
rect 34422 13444 34428 13456
rect 34379 13416 34428 13444
rect 34379 13413 34391 13416
rect 34333 13407 34391 13413
rect 34422 13404 34428 13416
rect 34480 13444 34486 13456
rect 35360 13444 35388 13472
rect 34480 13416 35388 13444
rect 34480 13404 34486 13416
rect 35802 13404 35808 13456
rect 35860 13404 35866 13456
rect 38102 13444 38108 13456
rect 37108 13416 38108 13444
rect 33183 13348 33364 13376
rect 33873 13379 33931 13385
rect 33183 13345 33195 13348
rect 33137 13339 33195 13345
rect 33873 13345 33885 13379
rect 33919 13376 33931 13379
rect 34238 13376 34244 13388
rect 33919 13348 34244 13376
rect 33919 13345 33931 13348
rect 33873 13339 33931 13345
rect 33008 13336 33014 13339
rect 34238 13336 34244 13348
rect 34296 13336 34302 13388
rect 35345 13379 35403 13385
rect 35345 13345 35357 13379
rect 35391 13376 35403 13379
rect 35820 13376 35848 13404
rect 35391 13348 35848 13376
rect 35391 13345 35403 13348
rect 35345 13339 35403 13345
rect 31665 13271 31723 13277
rect 32140 13280 32352 13308
rect 34057 13311 34115 13317
rect 32140 13252 32168 13280
rect 34057 13277 34069 13311
rect 34103 13308 34115 13311
rect 34606 13308 34612 13320
rect 34103 13280 34612 13308
rect 34103 13277 34115 13280
rect 34057 13271 34115 13277
rect 34606 13268 34612 13280
rect 34664 13268 34670 13320
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 35158 13308 35164 13320
rect 34848 13280 35164 13308
rect 34848 13268 34854 13280
rect 35158 13268 35164 13280
rect 35216 13268 35222 13320
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 36081 13311 36139 13317
rect 36081 13308 36093 13311
rect 35860 13280 36093 13308
rect 35860 13268 35866 13280
rect 36081 13277 36093 13280
rect 36127 13308 36139 13311
rect 37108 13308 37136 13416
rect 38102 13404 38108 13416
rect 38160 13404 38166 13456
rect 38396 13416 38608 13444
rect 38013 13379 38071 13385
rect 38013 13345 38025 13379
rect 38059 13376 38071 13379
rect 38396 13376 38424 13416
rect 38059 13348 38424 13376
rect 38059 13345 38071 13348
rect 38013 13339 38071 13345
rect 38470 13336 38476 13388
rect 38528 13336 38534 13388
rect 38580 13376 38608 13416
rect 39574 13376 39580 13388
rect 38580 13348 39580 13376
rect 39574 13336 39580 13348
rect 39632 13336 39638 13388
rect 40034 13336 40040 13388
rect 40092 13336 40098 13388
rect 42518 13336 42524 13388
rect 42576 13376 42582 13388
rect 42797 13379 42855 13385
rect 42797 13376 42809 13379
rect 42576 13348 42809 13376
rect 42576 13336 42582 13348
rect 42797 13345 42809 13348
rect 42843 13345 42855 13379
rect 42797 13339 42855 13345
rect 42981 13379 43039 13385
rect 42981 13345 42993 13379
rect 43027 13376 43039 13379
rect 43162 13376 43168 13388
rect 43027 13348 43168 13376
rect 43027 13345 43039 13348
rect 42981 13339 43039 13345
rect 43162 13336 43168 13348
rect 43220 13336 43226 13388
rect 43364 13376 43392 13475
rect 44266 13472 44272 13524
rect 44324 13472 44330 13524
rect 49142 13472 49148 13524
rect 49200 13512 49206 13524
rect 49237 13515 49295 13521
rect 49237 13512 49249 13515
rect 49200 13484 49249 13512
rect 49200 13472 49206 13484
rect 49237 13481 49249 13484
rect 49283 13512 49295 13515
rect 49510 13512 49516 13524
rect 49283 13484 49516 13512
rect 49283 13481 49295 13484
rect 49237 13475 49295 13481
rect 49510 13472 49516 13484
rect 49568 13472 49574 13524
rect 50893 13515 50951 13521
rect 50893 13481 50905 13515
rect 50939 13512 50951 13515
rect 51258 13512 51264 13524
rect 50939 13484 51264 13512
rect 50939 13481 50951 13484
rect 50893 13475 50951 13481
rect 51258 13472 51264 13484
rect 51316 13472 51322 13524
rect 55324 13484 56456 13512
rect 55324 13456 55352 13484
rect 51721 13447 51779 13453
rect 50356 13416 51672 13444
rect 50356 13388 50384 13416
rect 43625 13379 43683 13385
rect 43625 13376 43637 13379
rect 43364 13348 43637 13376
rect 43625 13345 43637 13348
rect 43671 13345 43683 13379
rect 43625 13339 43683 13345
rect 43806 13336 43812 13388
rect 43864 13336 43870 13388
rect 46290 13336 46296 13388
rect 46348 13376 46354 13388
rect 46385 13379 46443 13385
rect 46385 13376 46397 13379
rect 46348 13348 46397 13376
rect 46348 13336 46354 13348
rect 46385 13345 46397 13348
rect 46431 13345 46443 13379
rect 46385 13339 46443 13345
rect 36127 13280 37136 13308
rect 37829 13311 37887 13317
rect 36127 13277 36139 13280
rect 36081 13271 36139 13277
rect 37829 13277 37841 13311
rect 37875 13277 37887 13311
rect 37829 13271 37887 13277
rect 23523 13212 23704 13240
rect 23523 13209 23535 13212
rect 23477 13203 23535 13209
rect 23676 13184 23704 13212
rect 28936 13243 28994 13249
rect 28936 13209 28948 13243
rect 28982 13240 28994 13243
rect 29086 13240 29092 13252
rect 28982 13212 29092 13240
rect 28982 13209 28994 13212
rect 28936 13203 28994 13209
rect 29086 13200 29092 13212
rect 29144 13200 29150 13252
rect 30092 13243 30150 13249
rect 30092 13209 30104 13243
rect 30138 13240 30150 13243
rect 31294 13240 31300 13252
rect 30138 13212 31300 13240
rect 30138 13209 30150 13212
rect 30092 13203 30150 13209
rect 31294 13200 31300 13212
rect 31352 13200 31358 13252
rect 32122 13200 32128 13252
rect 32180 13200 32186 13252
rect 34146 13200 34152 13252
rect 34204 13200 34210 13252
rect 36348 13243 36406 13249
rect 36348 13209 36360 13243
rect 36394 13240 36406 13243
rect 36814 13240 36820 13252
rect 36394 13212 36820 13240
rect 36394 13209 36406 13212
rect 36348 13203 36406 13209
rect 36814 13200 36820 13212
rect 36872 13200 36878 13252
rect 7098 13132 7104 13184
rect 7156 13132 7162 13184
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11054 13172 11060 13184
rect 11011 13144 11060 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 11296 13144 11345 13172
rect 11296 13132 11302 13144
rect 11333 13141 11345 13144
rect 11379 13141 11391 13175
rect 11333 13135 11391 13141
rect 11885 13175 11943 13181
rect 11885 13141 11897 13175
rect 11931 13172 11943 13175
rect 13262 13172 13268 13184
rect 11931 13144 13268 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14458 13132 14464 13184
rect 14516 13132 14522 13184
rect 14826 13132 14832 13184
rect 14884 13132 14890 13184
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 19334 13172 19340 13184
rect 18187 13144 19340 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19610 13132 19616 13184
rect 19668 13132 19674 13184
rect 23566 13132 23572 13184
rect 23624 13132 23630 13184
rect 23658 13132 23664 13184
rect 23716 13132 23722 13184
rect 24762 13132 24768 13184
rect 24820 13132 24826 13184
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 26234 13172 26240 13184
rect 25832 13144 26240 13172
rect 25832 13132 25838 13144
rect 26234 13132 26240 13144
rect 26292 13172 26298 13184
rect 31110 13172 31116 13184
rect 26292 13144 31116 13172
rect 26292 13132 26298 13144
rect 31110 13132 31116 13144
rect 31168 13132 31174 13184
rect 32030 13132 32036 13184
rect 32088 13132 32094 13184
rect 32217 13175 32275 13181
rect 32217 13141 32229 13175
rect 32263 13172 32275 13175
rect 34164 13172 34192 13200
rect 32263 13144 34192 13172
rect 32263 13141 32275 13144
rect 32217 13135 32275 13141
rect 35066 13132 35072 13184
rect 35124 13132 35130 13184
rect 35158 13132 35164 13184
rect 35216 13132 35222 13184
rect 37844 13172 37872 13271
rect 38746 13268 38752 13320
rect 38804 13268 38810 13320
rect 38838 13268 38844 13320
rect 38896 13317 38902 13320
rect 38896 13311 38924 13317
rect 38912 13277 38924 13311
rect 38896 13271 38924 13277
rect 38896 13268 38902 13271
rect 39022 13268 39028 13320
rect 39080 13268 39086 13320
rect 40218 13268 40224 13320
rect 40276 13268 40282 13320
rect 40310 13268 40316 13320
rect 40368 13308 40374 13320
rect 40865 13311 40923 13317
rect 40865 13308 40877 13311
rect 40368 13280 40877 13308
rect 40368 13268 40374 13280
rect 40865 13277 40877 13280
rect 40911 13277 40923 13311
rect 43180 13308 43208 13336
rect 45554 13308 45560 13320
rect 43180 13280 45560 13308
rect 40865 13271 40923 13277
rect 45554 13268 45560 13280
rect 45612 13268 45618 13320
rect 45738 13268 45744 13320
rect 45796 13268 45802 13320
rect 46400 13308 46428 13339
rect 50338 13336 50344 13388
rect 50396 13336 50402 13388
rect 51077 13379 51135 13385
rect 51077 13345 51089 13379
rect 51123 13376 51135 13379
rect 51534 13376 51540 13388
rect 51123 13348 51540 13376
rect 51123 13345 51135 13348
rect 51077 13339 51135 13345
rect 51534 13336 51540 13348
rect 51592 13336 51598 13388
rect 47857 13311 47915 13317
rect 47857 13308 47869 13311
rect 46400 13280 47869 13308
rect 47857 13277 47869 13280
rect 47903 13308 47915 13311
rect 48590 13308 48596 13320
rect 47903 13280 48596 13308
rect 47903 13277 47915 13280
rect 47857 13271 47915 13277
rect 48590 13268 48596 13280
rect 48648 13268 48654 13320
rect 49694 13308 49700 13320
rect 49160 13280 49700 13308
rect 41132 13243 41190 13249
rect 39500 13212 40172 13240
rect 38194 13172 38200 13184
rect 37844 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 38562 13132 38568 13184
rect 38620 13172 38626 13184
rect 38838 13172 38844 13184
rect 38620 13144 38844 13172
rect 38620 13132 38626 13144
rect 38838 13132 38844 13144
rect 38896 13132 38902 13184
rect 38930 13132 38936 13184
rect 38988 13172 38994 13184
rect 39500 13172 39528 13212
rect 38988 13144 39528 13172
rect 38988 13132 38994 13144
rect 39666 13132 39672 13184
rect 39724 13132 39730 13184
rect 40144 13181 40172 13212
rect 41132 13209 41144 13243
rect 41178 13240 41190 13243
rect 41598 13240 41604 13252
rect 41178 13212 41604 13240
rect 41178 13209 41190 13212
rect 41132 13203 41190 13209
rect 41598 13200 41604 13212
rect 41656 13200 41662 13252
rect 43070 13240 43076 13252
rect 42260 13212 43076 13240
rect 40129 13175 40187 13181
rect 40129 13141 40141 13175
rect 40175 13141 40187 13175
rect 40129 13135 40187 13141
rect 40586 13132 40592 13184
rect 40644 13132 40650 13184
rect 42260 13181 42288 13212
rect 43070 13200 43076 13212
rect 43128 13200 43134 13252
rect 46652 13243 46710 13249
rect 46652 13209 46664 13243
rect 46698 13240 46710 13243
rect 46750 13240 46756 13252
rect 46698 13212 46756 13240
rect 46698 13209 46710 13212
rect 46652 13203 46710 13209
rect 46750 13200 46756 13212
rect 46808 13200 46814 13252
rect 48124 13243 48182 13249
rect 48124 13209 48136 13243
rect 48170 13240 48182 13243
rect 48406 13240 48412 13252
rect 48170 13212 48412 13240
rect 48170 13209 48182 13212
rect 48124 13203 48182 13209
rect 48406 13200 48412 13212
rect 48464 13200 48470 13252
rect 42245 13175 42303 13181
rect 42245 13141 42257 13175
rect 42291 13141 42303 13175
rect 42245 13135 42303 13141
rect 42334 13132 42340 13184
rect 42392 13132 42398 13184
rect 42705 13175 42763 13181
rect 42705 13141 42717 13175
rect 42751 13172 42763 13175
rect 43806 13172 43812 13184
rect 42751 13144 43812 13172
rect 42751 13141 42763 13144
rect 42705 13135 42763 13141
rect 43806 13132 43812 13144
rect 43864 13172 43870 13184
rect 43901 13175 43959 13181
rect 43901 13172 43913 13175
rect 43864 13144 43913 13172
rect 43864 13132 43870 13144
rect 43901 13141 43913 13144
rect 43947 13141 43959 13175
rect 43901 13135 43959 13141
rect 44818 13132 44824 13184
rect 44876 13132 44882 13184
rect 45186 13132 45192 13184
rect 45244 13132 45250 13184
rect 47765 13175 47823 13181
rect 47765 13141 47777 13175
rect 47811 13172 47823 13175
rect 49160 13172 49188 13280
rect 49694 13268 49700 13280
rect 49752 13308 49758 13320
rect 49881 13311 49939 13317
rect 49881 13308 49893 13311
rect 49752 13280 49893 13308
rect 49752 13268 49758 13280
rect 49881 13277 49893 13280
rect 49927 13277 49939 13311
rect 49881 13271 49939 13277
rect 50433 13311 50491 13317
rect 50433 13277 50445 13311
rect 50479 13308 50491 13311
rect 51166 13308 51172 13320
rect 50479 13280 51172 13308
rect 50479 13277 50491 13280
rect 50433 13271 50491 13277
rect 51166 13268 51172 13280
rect 51224 13268 51230 13320
rect 51644 13308 51672 13416
rect 51721 13413 51733 13447
rect 51767 13444 51779 13447
rect 52362 13444 52368 13456
rect 51767 13416 52368 13444
rect 51767 13413 51779 13416
rect 51721 13407 51779 13413
rect 52362 13404 52368 13416
rect 52420 13404 52426 13456
rect 54113 13447 54171 13453
rect 54113 13413 54125 13447
rect 54159 13444 54171 13447
rect 54159 13416 54984 13444
rect 54159 13413 54171 13416
rect 54113 13407 54171 13413
rect 54956 13388 54984 13416
rect 55306 13404 55312 13456
rect 55364 13404 55370 13456
rect 54297 13379 54355 13385
rect 54297 13376 54309 13379
rect 54128 13348 54309 13376
rect 54128 13320 54156 13348
rect 54297 13345 54309 13348
rect 54343 13345 54355 13379
rect 54297 13339 54355 13345
rect 54481 13379 54539 13385
rect 54481 13345 54493 13379
rect 54527 13376 54539 13379
rect 54754 13376 54760 13388
rect 54527 13348 54760 13376
rect 54527 13345 54539 13348
rect 54481 13339 54539 13345
rect 54754 13336 54760 13348
rect 54812 13336 54818 13388
rect 54938 13336 54944 13388
rect 54996 13376 55002 13388
rect 56091 13379 56149 13385
rect 56091 13376 56103 13379
rect 54996 13348 56103 13376
rect 54996 13336 55002 13348
rect 56091 13345 56103 13348
rect 56137 13345 56149 13379
rect 56091 13339 56149 13345
rect 56229 13379 56287 13385
rect 56229 13345 56241 13379
rect 56275 13376 56287 13379
rect 56428 13376 56456 13484
rect 58253 13447 58311 13453
rect 58253 13444 58265 13447
rect 56612 13416 58265 13444
rect 56612 13388 56640 13416
rect 56275 13348 56456 13376
rect 56275 13345 56287 13348
rect 56229 13339 56287 13345
rect 56502 13336 56508 13388
rect 56560 13336 56566 13388
rect 56594 13336 56600 13388
rect 56652 13336 56658 13388
rect 56965 13379 57023 13385
rect 56965 13345 56977 13379
rect 57011 13376 57023 13379
rect 57698 13376 57704 13388
rect 57011 13348 57704 13376
rect 57011 13345 57023 13348
rect 56965 13339 57023 13345
rect 57698 13336 57704 13348
rect 57756 13336 57762 13388
rect 57808 13385 57836 13416
rect 58253 13413 58265 13416
rect 58299 13413 58311 13447
rect 58253 13407 58311 13413
rect 57793 13379 57851 13385
rect 57793 13345 57805 13379
rect 57839 13345 57851 13379
rect 57793 13339 57851 13345
rect 52089 13311 52147 13317
rect 52089 13308 52101 13311
rect 51644 13280 52101 13308
rect 52089 13277 52101 13280
rect 52135 13308 52147 13311
rect 52270 13308 52276 13320
rect 52135 13280 52276 13308
rect 52135 13277 52147 13280
rect 52089 13271 52147 13277
rect 52270 13268 52276 13280
rect 52328 13268 52334 13320
rect 53006 13317 53012 13320
rect 52733 13311 52791 13317
rect 52733 13308 52745 13311
rect 52472 13280 52745 13308
rect 49234 13200 49240 13252
rect 49292 13240 49298 13252
rect 51353 13243 51411 13249
rect 51353 13240 51365 13243
rect 49292 13212 51365 13240
rect 49292 13200 49298 13212
rect 51353 13209 51365 13212
rect 51399 13209 51411 13243
rect 51353 13203 51411 13209
rect 52472 13184 52500 13280
rect 52733 13277 52745 13280
rect 52779 13277 52791 13311
rect 53000 13308 53012 13317
rect 52967 13280 53012 13308
rect 52733 13271 52791 13277
rect 53000 13271 53012 13280
rect 53006 13268 53012 13271
rect 53064 13268 53070 13320
rect 54110 13268 54116 13320
rect 54168 13268 54174 13320
rect 55950 13268 55956 13320
rect 56008 13268 56014 13320
rect 57146 13268 57152 13320
rect 57204 13268 57210 13320
rect 57606 13268 57612 13320
rect 57664 13268 57670 13320
rect 54573 13243 54631 13249
rect 54573 13209 54585 13243
rect 54619 13240 54631 13243
rect 57701 13243 57759 13249
rect 57701 13240 57713 13243
rect 54619 13212 55168 13240
rect 54619 13209 54631 13212
rect 54573 13203 54631 13209
rect 55140 13184 55168 13212
rect 56980 13212 57713 13240
rect 47811 13144 49188 13172
rect 47811 13141 47823 13144
rect 47765 13135 47823 13141
rect 49326 13132 49332 13184
rect 49384 13132 49390 13184
rect 50522 13132 50528 13184
rect 50580 13132 50586 13184
rect 50798 13132 50804 13184
rect 50856 13172 50862 13184
rect 51261 13175 51319 13181
rect 51261 13172 51273 13175
rect 50856 13144 51273 13172
rect 50856 13132 50862 13144
rect 51261 13141 51273 13144
rect 51307 13141 51319 13175
rect 51261 13135 51319 13141
rect 52454 13132 52460 13184
rect 52512 13132 52518 13184
rect 54938 13132 54944 13184
rect 54996 13132 55002 13184
rect 55122 13132 55128 13184
rect 55180 13132 55186 13184
rect 55309 13175 55367 13181
rect 55309 13141 55321 13175
rect 55355 13172 55367 13175
rect 56980 13172 57008 13212
rect 57701 13209 57713 13212
rect 57747 13209 57759 13243
rect 57701 13203 57759 13209
rect 55355 13144 57008 13172
rect 57241 13175 57299 13181
rect 55355 13141 55367 13144
rect 55309 13135 55367 13141
rect 57241 13141 57253 13175
rect 57287 13172 57299 13175
rect 57514 13172 57520 13184
rect 57287 13144 57520 13172
rect 57287 13141 57299 13144
rect 57241 13135 57299 13141
rect 57514 13132 57520 13144
rect 57572 13132 57578 13184
rect 1104 13082 59040 13104
rect 1104 13030 15394 13082
rect 15446 13030 15458 13082
rect 15510 13030 15522 13082
rect 15574 13030 15586 13082
rect 15638 13030 15650 13082
rect 15702 13030 29838 13082
rect 29890 13030 29902 13082
rect 29954 13030 29966 13082
rect 30018 13030 30030 13082
rect 30082 13030 30094 13082
rect 30146 13030 44282 13082
rect 44334 13030 44346 13082
rect 44398 13030 44410 13082
rect 44462 13030 44474 13082
rect 44526 13030 44538 13082
rect 44590 13030 58726 13082
rect 58778 13030 58790 13082
rect 58842 13030 58854 13082
rect 58906 13030 58918 13082
rect 58970 13030 58982 13082
rect 59034 13030 59040 13082
rect 1104 13008 59040 13030
rect 2038 12928 2044 12980
rect 2096 12928 2102 12980
rect 6365 12971 6423 12977
rect 6365 12937 6377 12971
rect 6411 12968 6423 12971
rect 6454 12968 6460 12980
rect 6411 12940 6460 12968
rect 6411 12937 6423 12940
rect 6365 12931 6423 12937
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11146 12968 11152 12980
rect 11011 12940 11152 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 11388 12940 12817 12968
rect 11388 12928 11394 12940
rect 12805 12937 12817 12940
rect 12851 12937 12863 12971
rect 12805 12931 12863 12937
rect 2056 12900 2084 12928
rect 8018 12900 8024 12912
rect 1596 12872 2084 12900
rect 4172 12872 5304 12900
rect 1596 12841 1624 12872
rect 4172 12844 4200 12872
rect 1854 12841 1860 12844
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1848 12795 1860 12841
rect 1854 12792 1860 12795
rect 1912 12792 1918 12844
rect 4154 12792 4160 12844
rect 4212 12792 4218 12844
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 5276 12841 5304 12872
rect 7760 12872 8024 12900
rect 7760 12841 7788 12872
rect 8018 12860 8024 12872
rect 8076 12900 8082 12912
rect 8113 12903 8171 12909
rect 8113 12900 8125 12903
rect 8076 12872 8125 12900
rect 8076 12860 8082 12872
rect 8113 12869 8125 12872
rect 8159 12900 8171 12903
rect 11348 12900 11376 12928
rect 12158 12900 12164 12912
rect 8159 12872 11376 12900
rect 12084 12872 12164 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 9600 12841 9628 12872
rect 9858 12841 9864 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4488 12804 5089 12832
rect 4488 12792 4494 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12832 6239 12835
rect 7478 12835 7536 12841
rect 7478 12832 7490 12835
rect 6227 12804 7490 12832
rect 6227 12801 6239 12804
rect 6181 12795 6239 12801
rect 7478 12801 7490 12804
rect 7524 12801 7536 12835
rect 7478 12795 7536 12801
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12801 9643 12835
rect 9852 12832 9864 12841
rect 9819 12804 9864 12832
rect 9585 12795 9643 12801
rect 9852 12795 9864 12804
rect 9858 12792 9864 12795
rect 9916 12792 9922 12844
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 12084 12841 12112 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 12268 12872 12449 12900
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11296 12804 11529 12832
rect 11296 12792 11302 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2976 12736 3065 12764
rect 2976 12705 3004 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 5534 12724 5540 12776
rect 5592 12724 5598 12776
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 12268 12764 12296 12872
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12820 12900 12848 12931
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 13630 12968 13636 12980
rect 13504 12940 13636 12968
rect 13504 12928 13510 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14826 12928 14832 12980
rect 14884 12928 14890 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18322 12968 18328 12980
rect 18095 12940 18328 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18322 12928 18328 12940
rect 18380 12968 18386 12980
rect 19058 12968 19064 12980
rect 18380 12940 19064 12968
rect 18380 12928 18386 12940
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 20162 12968 20168 12980
rect 19392 12940 20168 12968
rect 19392 12928 19398 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20622 12928 20628 12980
rect 20680 12928 20686 12980
rect 23566 12928 23572 12980
rect 23624 12928 23630 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 24820 12940 24869 12968
rect 24820 12928 24826 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 24857 12931 24915 12937
rect 25866 12928 25872 12980
rect 25924 12968 25930 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 25924 12940 26341 12968
rect 25924 12928 25930 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 26329 12931 26387 12937
rect 26602 12928 26608 12980
rect 26660 12928 26666 12980
rect 26789 12971 26847 12977
rect 26789 12937 26801 12971
rect 26835 12968 26847 12971
rect 27614 12968 27620 12980
rect 26835 12940 27620 12968
rect 26835 12937 26847 12940
rect 26789 12931 26847 12937
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 27801 12971 27859 12977
rect 27801 12937 27813 12971
rect 27847 12968 27859 12971
rect 28166 12968 28172 12980
rect 27847 12940 28172 12968
rect 27847 12937 27859 12940
rect 27801 12931 27859 12937
rect 28166 12928 28172 12940
rect 28224 12928 28230 12980
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29273 12971 29331 12977
rect 29273 12968 29285 12971
rect 29144 12940 29285 12968
rect 29144 12928 29150 12940
rect 29273 12937 29285 12940
rect 29319 12937 29331 12971
rect 29273 12931 29331 12937
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 31662 12968 31668 12980
rect 29788 12940 31668 12968
rect 29788 12928 29794 12940
rect 14366 12900 14372 12912
rect 12820 12872 14372 12900
rect 12437 12863 12495 12869
rect 14366 12860 14372 12872
rect 14424 12900 14430 12912
rect 14424 12872 14504 12900
rect 14424 12860 14430 12872
rect 13078 12832 13084 12844
rect 11664 12736 12296 12764
rect 12406 12804 13084 12832
rect 11664 12724 11670 12736
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12665 3019 12699
rect 2961 12659 3019 12665
rect 3694 12588 3700 12640
rect 3752 12588 3758 12640
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12406 12628 12434 12804
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 14476 12841 14504 12872
rect 14205 12835 14263 12841
rect 14205 12801 14217 12835
rect 14251 12832 14263 12835
rect 14461 12835 14519 12841
rect 14251 12804 14412 12832
rect 14251 12801 14263 12804
rect 14205 12795 14263 12801
rect 14384 12764 14412 12804
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14844 12832 14872 12928
rect 16942 12909 16948 12912
rect 16936 12900 16948 12909
rect 16903 12872 16948 12900
rect 16936 12863 16948 12872
rect 16942 12860 16948 12863
rect 17000 12860 17006 12912
rect 18414 12860 18420 12912
rect 18472 12860 18478 12912
rect 20254 12860 20260 12912
rect 20312 12860 20318 12912
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14844 12804 15117 12832
rect 14461 12795 14519 12801
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 16298 12792 16304 12844
rect 16356 12832 16362 12844
rect 16666 12832 16672 12844
rect 16356 12804 16672 12832
rect 16356 12792 16362 12804
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12832 18383 12835
rect 18432 12832 18460 12860
rect 18371 12804 18460 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 19058 12792 19064 12844
rect 19116 12841 19122 12844
rect 19116 12835 19165 12841
rect 19116 12801 19119 12835
rect 19153 12801 19165 12835
rect 19116 12795 19165 12801
rect 19116 12792 19122 12795
rect 19242 12792 19248 12844
rect 19300 12792 19306 12844
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20640 12832 20668 12928
rect 20027 12804 20668 12832
rect 23584 12832 23612 12928
rect 26620 12900 26648 12928
rect 25516 12872 26648 12900
rect 25516 12841 25544 12872
rect 23641 12835 23699 12841
rect 23641 12832 23653 12835
rect 23584 12804 23653 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 23641 12801 23653 12804
rect 23687 12801 23699 12835
rect 23641 12795 23699 12801
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12801 25559 12835
rect 25501 12795 25559 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14384 12736 14565 12764
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 14553 12727 14611 12733
rect 18616 12736 18981 12764
rect 15565 12699 15623 12705
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 15746 12696 15752 12708
rect 15611 12668 15752 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 15746 12656 15752 12668
rect 15804 12696 15810 12708
rect 15804 12668 16344 12696
rect 15804 12656 15810 12668
rect 16316 12640 16344 12668
rect 11296 12600 12434 12628
rect 13081 12631 13139 12637
rect 11296 12588 11302 12600
rect 13081 12597 13093 12631
rect 13127 12628 13139 12631
rect 14090 12628 14096 12640
rect 13127 12600 14096 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 16114 12588 16120 12640
rect 16172 12588 16178 12640
rect 16298 12588 16304 12640
rect 16356 12588 16362 12640
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 18616 12628 18644 12736
rect 18969 12733 18981 12736
rect 19015 12764 19027 12767
rect 19521 12767 19579 12773
rect 19015 12736 19472 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 19444 12696 19472 12736
rect 19521 12733 19533 12767
rect 19567 12764 19579 12767
rect 19812 12764 19840 12792
rect 19567 12736 19840 12764
rect 20165 12767 20223 12773
rect 19567 12733 19579 12736
rect 19521 12727 19579 12733
rect 20165 12733 20177 12767
rect 20211 12764 20223 12767
rect 20622 12764 20628 12776
rect 20211 12736 20628 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 20806 12724 20812 12776
rect 20864 12724 20870 12776
rect 23385 12767 23443 12773
rect 23385 12764 23397 12767
rect 23216 12736 23397 12764
rect 19886 12696 19892 12708
rect 19444 12668 19892 12696
rect 19886 12656 19892 12668
rect 19944 12696 19950 12708
rect 22186 12696 22192 12708
rect 19944 12668 22192 12696
rect 19944 12656 19950 12668
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 23216 12640 23244 12736
rect 23385 12733 23397 12736
rect 23431 12733 23443 12767
rect 23385 12727 23443 12733
rect 24765 12699 24823 12705
rect 24765 12665 24777 12699
rect 24811 12696 24823 12699
rect 25516 12696 25544 12795
rect 25774 12724 25780 12776
rect 25832 12764 25838 12776
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 25832 12736 25881 12764
rect 25832 12724 25838 12736
rect 25869 12733 25881 12736
rect 25915 12733 25927 12767
rect 25869 12727 25927 12733
rect 26145 12767 26203 12773
rect 26145 12733 26157 12767
rect 26191 12733 26203 12767
rect 26436 12764 26464 12795
rect 27890 12792 27896 12844
rect 27948 12832 27954 12844
rect 29638 12832 29644 12844
rect 27948 12804 29644 12832
rect 27948 12792 27954 12804
rect 29638 12792 29644 12804
rect 29696 12792 29702 12844
rect 29840 12841 29868 12940
rect 31662 12928 31668 12940
rect 31720 12968 31726 12980
rect 32306 12968 32312 12980
rect 31720 12940 32312 12968
rect 31720 12928 31726 12940
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 34241 12971 34299 12977
rect 34241 12937 34253 12971
rect 34287 12968 34299 12971
rect 34330 12968 34336 12980
rect 34287 12940 34336 12968
rect 34287 12937 34299 12940
rect 34241 12931 34299 12937
rect 34330 12928 34336 12940
rect 34388 12928 34394 12980
rect 34609 12971 34667 12977
rect 34609 12937 34621 12971
rect 34655 12968 34667 12971
rect 35250 12968 35256 12980
rect 34655 12940 35256 12968
rect 34655 12937 34667 12940
rect 34609 12931 34667 12937
rect 35250 12928 35256 12940
rect 35308 12928 35314 12980
rect 37093 12971 37151 12977
rect 37093 12937 37105 12971
rect 37139 12968 37151 12971
rect 38562 12968 38568 12980
rect 37139 12940 38568 12968
rect 37139 12937 37151 12940
rect 37093 12931 37151 12937
rect 38562 12928 38568 12940
rect 38620 12928 38626 12980
rect 38749 12971 38807 12977
rect 38749 12937 38761 12971
rect 38795 12968 38807 12971
rect 39574 12968 39580 12980
rect 38795 12940 39580 12968
rect 38795 12937 38807 12940
rect 38749 12931 38807 12937
rect 39574 12928 39580 12940
rect 39632 12928 39638 12980
rect 41598 12928 41604 12980
rect 41656 12928 41662 12980
rect 42334 12928 42340 12980
rect 42392 12928 42398 12980
rect 43070 12928 43076 12980
rect 43128 12968 43134 12980
rect 43990 12968 43996 12980
rect 43128 12940 43996 12968
rect 43128 12928 43134 12940
rect 43990 12928 43996 12940
rect 44048 12928 44054 12980
rect 45005 12971 45063 12977
rect 45005 12937 45017 12971
rect 45051 12968 45063 12971
rect 45738 12968 45744 12980
rect 45051 12940 45744 12968
rect 45051 12937 45063 12940
rect 45005 12931 45063 12937
rect 30092 12903 30150 12909
rect 30092 12869 30104 12903
rect 30138 12900 30150 12903
rect 30282 12900 30288 12912
rect 30138 12872 30288 12900
rect 30138 12869 30150 12872
rect 30092 12863 30150 12869
rect 30282 12860 30288 12872
rect 30340 12860 30346 12912
rect 31294 12860 31300 12912
rect 31352 12860 31358 12912
rect 32030 12860 32036 12912
rect 32088 12860 32094 12912
rect 33904 12903 33962 12909
rect 33904 12869 33916 12903
rect 33950 12900 33962 12903
rect 34698 12900 34704 12912
rect 33950 12872 34704 12900
rect 33950 12869 33962 12872
rect 33904 12863 33962 12869
rect 34698 12860 34704 12872
rect 34756 12860 34762 12912
rect 35980 12903 36038 12909
rect 35980 12869 35992 12903
rect 36026 12900 36038 12903
rect 36446 12900 36452 12912
rect 36026 12872 36452 12900
rect 36026 12869 36038 12872
rect 35980 12863 36038 12869
rect 36446 12860 36452 12872
rect 36504 12860 36510 12912
rect 37550 12860 37556 12912
rect 37608 12900 37614 12912
rect 37645 12903 37703 12909
rect 37645 12900 37657 12903
rect 37608 12872 37657 12900
rect 37608 12860 37614 12872
rect 37645 12869 37657 12872
rect 37691 12900 37703 12903
rect 37734 12900 37740 12912
rect 37691 12872 37740 12900
rect 37691 12869 37703 12872
rect 37645 12863 37703 12869
rect 37734 12860 37740 12872
rect 37792 12860 37798 12912
rect 37826 12860 37832 12912
rect 37884 12860 37890 12912
rect 38010 12860 38016 12912
rect 38068 12900 38074 12912
rect 39022 12900 39028 12912
rect 38068 12872 39028 12900
rect 38068 12860 38074 12872
rect 39022 12860 39028 12872
rect 39080 12860 39086 12912
rect 39884 12903 39942 12909
rect 39884 12869 39896 12903
rect 39930 12900 39942 12903
rect 40221 12903 40279 12909
rect 40221 12900 40233 12903
rect 39930 12872 40233 12900
rect 39930 12869 39942 12872
rect 39884 12863 39942 12869
rect 40221 12869 40233 12872
rect 40267 12869 40279 12903
rect 40221 12863 40279 12869
rect 29825 12835 29883 12841
rect 29825 12801 29837 12835
rect 29871 12801 29883 12835
rect 29825 12795 29883 12801
rect 31941 12835 31999 12841
rect 31941 12801 31953 12835
rect 31987 12832 31999 12835
rect 32048 12832 32076 12860
rect 34330 12832 34336 12844
rect 31987 12804 32076 12832
rect 33152 12804 34336 12832
rect 31987 12801 31999 12804
rect 31941 12795 31999 12801
rect 27338 12764 27344 12776
rect 26436 12736 27344 12764
rect 26145 12727 26203 12733
rect 26160 12696 26188 12727
rect 27338 12724 27344 12736
rect 27396 12724 27402 12776
rect 27617 12767 27675 12773
rect 27617 12733 27629 12767
rect 27663 12733 27675 12767
rect 28629 12767 28687 12773
rect 28629 12764 28641 12767
rect 27617 12727 27675 12733
rect 28276 12736 28641 12764
rect 27062 12696 27068 12708
rect 24811 12668 25544 12696
rect 25884 12668 27068 12696
rect 24811 12665 24823 12668
rect 24765 12659 24823 12665
rect 25884 12640 25912 12668
rect 27062 12656 27068 12668
rect 27120 12656 27126 12708
rect 16448 12600 18644 12628
rect 16448 12588 16454 12600
rect 21174 12588 21180 12640
rect 21232 12588 21238 12640
rect 23198 12588 23204 12640
rect 23256 12588 23262 12640
rect 25866 12588 25872 12640
rect 25924 12588 25930 12640
rect 27430 12588 27436 12640
rect 27488 12628 27494 12640
rect 27632 12628 27660 12727
rect 28276 12705 28304 12736
rect 28629 12733 28641 12736
rect 28675 12733 28687 12767
rect 28629 12727 28687 12733
rect 31478 12724 31484 12776
rect 31536 12764 31542 12776
rect 33152 12764 33180 12804
rect 34330 12792 34336 12804
rect 34388 12832 34394 12844
rect 35066 12832 35072 12844
rect 34388 12804 35072 12832
rect 34388 12792 34394 12804
rect 31536 12736 33180 12764
rect 34149 12767 34207 12773
rect 31536 12724 31542 12736
rect 34149 12733 34161 12767
rect 34195 12764 34207 12767
rect 34514 12764 34520 12776
rect 34195 12736 34520 12764
rect 34195 12733 34207 12736
rect 34149 12727 34207 12733
rect 34514 12724 34520 12736
rect 34572 12724 34578 12776
rect 34716 12773 34744 12804
rect 35066 12792 35072 12804
rect 35124 12792 35130 12844
rect 35713 12835 35771 12841
rect 35713 12801 35725 12835
rect 35759 12832 35771 12835
rect 35802 12832 35808 12844
rect 35759 12804 35808 12832
rect 35759 12801 35771 12804
rect 35713 12795 35771 12801
rect 35802 12792 35808 12804
rect 35860 12792 35866 12844
rect 37844 12832 37872 12860
rect 39574 12832 39580 12844
rect 37844 12804 39580 12832
rect 39574 12792 39580 12804
rect 39632 12792 39638 12844
rect 42245 12835 42303 12841
rect 42245 12801 42257 12835
rect 42291 12832 42303 12835
rect 42352 12832 42380 12928
rect 43898 12841 43904 12844
rect 42291 12804 42380 12832
rect 43876 12835 43904 12841
rect 42291 12801 42303 12804
rect 42245 12795 42303 12801
rect 43876 12801 43888 12835
rect 43876 12795 43904 12801
rect 43898 12792 43904 12795
rect 43956 12792 43962 12844
rect 43990 12792 43996 12844
rect 44048 12792 44054 12844
rect 44729 12835 44787 12841
rect 44729 12801 44741 12835
rect 44775 12832 44787 12835
rect 45020 12832 45048 12931
rect 45738 12928 45744 12940
rect 45796 12928 45802 12980
rect 47394 12928 47400 12980
rect 47452 12968 47458 12980
rect 47581 12971 47639 12977
rect 47581 12968 47593 12971
rect 47452 12940 47593 12968
rect 47452 12928 47458 12940
rect 47581 12937 47593 12940
rect 47627 12937 47639 12971
rect 47581 12931 47639 12937
rect 47946 12928 47952 12980
rect 48004 12928 48010 12980
rect 48590 12928 48596 12980
rect 48648 12928 48654 12980
rect 49326 12968 49332 12980
rect 48700 12940 49332 12968
rect 46140 12903 46198 12909
rect 46140 12869 46152 12903
rect 46186 12900 46198 12903
rect 46477 12903 46535 12909
rect 46477 12900 46489 12903
rect 46186 12872 46489 12900
rect 46186 12869 46198 12872
rect 46140 12863 46198 12869
rect 46477 12869 46489 12872
rect 46523 12869 46535 12903
rect 46477 12863 46535 12869
rect 48041 12903 48099 12909
rect 48041 12869 48053 12903
rect 48087 12900 48099 12903
rect 48700 12900 48728 12940
rect 49326 12928 49332 12940
rect 49384 12928 49390 12980
rect 50522 12928 50528 12980
rect 50580 12968 50586 12980
rect 50985 12971 51043 12977
rect 50985 12968 50997 12971
rect 50580 12940 50997 12968
rect 50580 12928 50586 12940
rect 50985 12937 50997 12940
rect 51031 12968 51043 12971
rect 51074 12968 51080 12980
rect 51031 12940 51080 12968
rect 51031 12937 51043 12940
rect 50985 12931 51043 12937
rect 51074 12928 51080 12940
rect 51132 12928 51138 12980
rect 51534 12928 51540 12980
rect 51592 12968 51598 12980
rect 52270 12968 52276 12980
rect 51592 12940 52276 12968
rect 51592 12928 51598 12940
rect 52270 12928 52276 12940
rect 52328 12968 52334 12980
rect 52457 12971 52515 12977
rect 52457 12968 52469 12971
rect 52328 12940 52469 12968
rect 52328 12928 52334 12940
rect 52457 12937 52469 12940
rect 52503 12937 52515 12971
rect 52457 12931 52515 12937
rect 54938 12928 54944 12980
rect 54996 12928 55002 12980
rect 55214 12928 55220 12980
rect 55272 12968 55278 12980
rect 56502 12968 56508 12980
rect 55272 12940 56508 12968
rect 55272 12928 55278 12940
rect 56502 12928 56508 12940
rect 56560 12928 56566 12980
rect 56778 12928 56784 12980
rect 56836 12928 56842 12980
rect 57146 12928 57152 12980
rect 57204 12968 57210 12980
rect 57517 12971 57575 12977
rect 57517 12968 57529 12971
rect 57204 12940 57529 12968
rect 57204 12928 57210 12940
rect 57517 12937 57529 12940
rect 57563 12937 57575 12971
rect 57517 12931 57575 12937
rect 48087 12872 48728 12900
rect 48087 12869 48099 12872
rect 48041 12863 48099 12869
rect 44775 12804 45048 12832
rect 44775 12801 44787 12804
rect 44729 12795 44787 12801
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 46385 12835 46443 12841
rect 46385 12832 46397 12835
rect 46348 12804 46397 12832
rect 46348 12792 46354 12804
rect 46385 12801 46397 12804
rect 46431 12832 46443 12835
rect 46842 12832 46848 12844
rect 46431 12804 46848 12832
rect 46431 12801 46443 12804
rect 46385 12795 46443 12801
rect 46842 12792 46848 12804
rect 46900 12792 46906 12844
rect 49418 12792 49424 12844
rect 49476 12792 49482 12844
rect 49510 12792 49516 12844
rect 49568 12841 49574 12844
rect 49568 12835 49617 12841
rect 49568 12801 49571 12835
rect 49605 12801 49617 12835
rect 49568 12795 49617 12801
rect 49568 12792 49574 12795
rect 49694 12792 49700 12844
rect 49752 12792 49758 12844
rect 50614 12792 50620 12844
rect 50672 12792 50678 12844
rect 54956 12841 54984 12928
rect 55122 12860 55128 12912
rect 55180 12900 55186 12912
rect 56796 12900 56824 12928
rect 55180 12872 56824 12900
rect 55180 12860 55186 12872
rect 51077 12835 51135 12841
rect 51077 12801 51089 12835
rect 51123 12832 51135 12835
rect 51537 12835 51595 12841
rect 51537 12832 51549 12835
rect 51123 12804 51549 12832
rect 51123 12801 51135 12804
rect 51077 12795 51135 12801
rect 51537 12801 51549 12804
rect 51583 12801 51595 12835
rect 51537 12795 51595 12801
rect 53092 12835 53150 12841
rect 53092 12801 53104 12835
rect 53138 12832 53150 12835
rect 54297 12835 54355 12841
rect 54297 12832 54309 12835
rect 53138 12804 54309 12832
rect 53138 12801 53150 12804
rect 53092 12795 53150 12801
rect 54297 12801 54309 12804
rect 54343 12801 54355 12835
rect 54297 12795 54355 12801
rect 54941 12835 54999 12841
rect 54941 12801 54953 12835
rect 54987 12801 54999 12835
rect 54941 12795 54999 12801
rect 55677 12835 55735 12841
rect 55677 12801 55689 12835
rect 55723 12832 55735 12835
rect 55950 12832 55956 12844
rect 55723 12804 55956 12832
rect 55723 12801 55735 12804
rect 55677 12795 55735 12801
rect 55950 12792 55956 12804
rect 56008 12792 56014 12844
rect 56045 12835 56103 12841
rect 56045 12801 56057 12835
rect 56091 12832 56103 12835
rect 56134 12832 56140 12844
rect 56091 12804 56140 12832
rect 56091 12801 56103 12804
rect 56045 12795 56103 12801
rect 56134 12792 56140 12804
rect 56192 12792 56198 12844
rect 56404 12835 56462 12841
rect 56404 12801 56416 12835
rect 56450 12832 56462 12835
rect 57238 12832 57244 12844
rect 56450 12804 57244 12832
rect 56450 12801 56462 12804
rect 56404 12795 56462 12801
rect 57238 12792 57244 12804
rect 57296 12792 57302 12844
rect 57532 12832 57560 12931
rect 58437 12835 58495 12841
rect 58437 12832 58449 12835
rect 57532 12804 58449 12832
rect 58437 12801 58449 12804
rect 58483 12801 58495 12835
rect 58437 12795 58495 12801
rect 34701 12767 34759 12773
rect 34701 12733 34713 12767
rect 34747 12733 34759 12767
rect 34701 12727 34759 12733
rect 34885 12767 34943 12773
rect 34885 12733 34897 12767
rect 34931 12764 34943 12767
rect 35345 12767 35403 12773
rect 35345 12764 35357 12767
rect 34931 12736 35357 12764
rect 34931 12733 34943 12736
rect 34885 12727 34943 12733
rect 35345 12733 35357 12736
rect 35391 12764 35403 12767
rect 35526 12764 35532 12776
rect 35391 12736 35532 12764
rect 35391 12733 35403 12736
rect 35345 12727 35403 12733
rect 35526 12724 35532 12736
rect 35584 12724 35590 12776
rect 37734 12724 37740 12776
rect 37792 12724 37798 12776
rect 37921 12767 37979 12773
rect 37921 12733 37933 12767
rect 37967 12764 37979 12767
rect 40129 12767 40187 12773
rect 37967 12736 38654 12764
rect 37967 12733 37979 12736
rect 37921 12727 37979 12733
rect 28261 12699 28319 12705
rect 28261 12665 28273 12699
rect 28307 12665 28319 12699
rect 28261 12659 28319 12665
rect 31202 12656 31208 12708
rect 31260 12656 31266 12708
rect 36722 12656 36728 12708
rect 36780 12696 36786 12708
rect 37936 12696 37964 12727
rect 36780 12668 37964 12696
rect 36780 12656 36786 12668
rect 28718 12628 28724 12640
rect 27488 12600 28724 12628
rect 27488 12588 27494 12600
rect 28718 12588 28724 12600
rect 28776 12628 28782 12640
rect 32398 12628 32404 12640
rect 28776 12600 32404 12628
rect 28776 12588 28782 12600
rect 32398 12588 32404 12600
rect 32456 12588 32462 12640
rect 32769 12631 32827 12637
rect 32769 12597 32781 12631
rect 32815 12628 32827 12631
rect 34606 12628 34612 12640
rect 32815 12600 34612 12628
rect 32815 12597 32827 12600
rect 32769 12591 32827 12597
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 37277 12631 37335 12637
rect 37277 12597 37289 12631
rect 37323 12628 37335 12631
rect 37458 12628 37464 12640
rect 37323 12600 37464 12628
rect 37323 12597 37335 12600
rect 37277 12591 37335 12597
rect 37458 12588 37464 12600
rect 37516 12588 37522 12640
rect 37642 12588 37648 12640
rect 37700 12628 37706 12640
rect 38289 12631 38347 12637
rect 38289 12628 38301 12631
rect 37700 12600 38301 12628
rect 37700 12588 37706 12600
rect 38289 12597 38301 12600
rect 38335 12628 38347 12631
rect 38470 12628 38476 12640
rect 38335 12600 38476 12628
rect 38335 12597 38347 12600
rect 38289 12591 38347 12597
rect 38470 12588 38476 12600
rect 38528 12588 38534 12640
rect 38626 12628 38654 12736
rect 40129 12733 40141 12767
rect 40175 12764 40187 12767
rect 40310 12764 40316 12776
rect 40175 12736 40316 12764
rect 40175 12733 40187 12736
rect 40129 12727 40187 12733
rect 40310 12724 40316 12736
rect 40368 12724 40374 12776
rect 40586 12724 40592 12776
rect 40644 12764 40650 12776
rect 40773 12767 40831 12773
rect 40773 12764 40785 12767
rect 40644 12736 40785 12764
rect 40644 12724 40650 12736
rect 40773 12733 40785 12736
rect 40819 12733 40831 12767
rect 40773 12727 40831 12733
rect 41230 12724 41236 12776
rect 41288 12764 41294 12776
rect 42610 12764 42616 12776
rect 41288 12736 42616 12764
rect 41288 12724 41294 12736
rect 42610 12724 42616 12736
rect 42668 12724 42674 12776
rect 43717 12767 43775 12773
rect 43717 12733 43729 12767
rect 43763 12764 43775 12767
rect 44818 12764 44824 12776
rect 43763 12736 44824 12764
rect 43763 12733 43775 12736
rect 43717 12727 43775 12733
rect 44818 12724 44824 12736
rect 44876 12724 44882 12776
rect 44910 12724 44916 12776
rect 44968 12724 44974 12776
rect 47026 12724 47032 12776
rect 47084 12724 47090 12776
rect 47394 12724 47400 12776
rect 47452 12764 47458 12776
rect 48133 12767 48191 12773
rect 48133 12764 48145 12767
rect 47452 12736 48145 12764
rect 47452 12724 47458 12736
rect 48133 12733 48145 12736
rect 48179 12733 48191 12767
rect 48133 12727 48191 12733
rect 48777 12767 48835 12773
rect 48777 12733 48789 12767
rect 48823 12764 48835 12767
rect 49234 12764 49240 12776
rect 48823 12736 49240 12764
rect 48823 12733 48835 12736
rect 48777 12727 48835 12733
rect 49234 12724 49240 12736
rect 49292 12724 49298 12776
rect 49970 12764 49976 12776
rect 49896 12736 49976 12764
rect 42242 12656 42248 12708
rect 42300 12656 42306 12708
rect 44269 12699 44327 12705
rect 44269 12665 44281 12699
rect 44315 12696 44327 12699
rect 44315 12668 45508 12696
rect 44315 12665 44327 12668
rect 44269 12659 44327 12665
rect 42260 12628 42288 12656
rect 45480 12640 45508 12668
rect 38626 12600 42288 12628
rect 43073 12631 43131 12637
rect 43073 12597 43085 12631
rect 43119 12628 43131 12631
rect 44726 12628 44732 12640
rect 43119 12600 44732 12628
rect 43119 12597 43131 12600
rect 43073 12591 43131 12597
rect 44726 12588 44732 12600
rect 44784 12588 44790 12640
rect 45462 12588 45468 12640
rect 45520 12588 45526 12640
rect 47210 12588 47216 12640
rect 47268 12628 47274 12640
rect 48498 12628 48504 12640
rect 47268 12600 48504 12628
rect 47268 12588 47274 12600
rect 48498 12588 48504 12600
rect 48556 12628 48562 12640
rect 49896 12628 49924 12736
rect 49970 12724 49976 12736
rect 50028 12724 50034 12776
rect 50430 12724 50436 12776
rect 50488 12724 50494 12776
rect 50893 12767 50951 12773
rect 50893 12733 50905 12767
rect 50939 12764 50951 12767
rect 51350 12764 51356 12776
rect 50939 12736 51356 12764
rect 50939 12733 50951 12736
rect 50893 12727 50951 12733
rect 51350 12724 51356 12736
rect 51408 12724 51414 12776
rect 52089 12767 52147 12773
rect 52089 12733 52101 12767
rect 52135 12733 52147 12767
rect 52089 12727 52147 12733
rect 50448 12696 50476 12724
rect 52104 12696 52132 12727
rect 52454 12724 52460 12776
rect 52512 12764 52518 12776
rect 52825 12767 52883 12773
rect 52825 12764 52837 12767
rect 52512 12736 52837 12764
rect 52512 12724 52518 12736
rect 52825 12733 52837 12736
rect 52871 12733 52883 12767
rect 52825 12727 52883 12733
rect 50448 12668 52132 12696
rect 54205 12699 54263 12705
rect 54205 12665 54217 12699
rect 54251 12696 54263 12699
rect 55306 12696 55312 12708
rect 54251 12668 55312 12696
rect 54251 12665 54263 12668
rect 54205 12659 54263 12665
rect 55306 12656 55312 12668
rect 55364 12656 55370 12708
rect 48556 12600 49924 12628
rect 51445 12631 51503 12637
rect 48556 12588 48562 12600
rect 51445 12597 51457 12631
rect 51491 12628 51503 12631
rect 52178 12628 52184 12640
rect 51491 12600 52184 12628
rect 51491 12597 51503 12600
rect 51445 12591 51503 12597
rect 52178 12588 52184 12600
rect 52236 12588 52242 12640
rect 55214 12588 55220 12640
rect 55272 12588 55278 12640
rect 57606 12588 57612 12640
rect 57664 12628 57670 12640
rect 57885 12631 57943 12637
rect 57885 12628 57897 12631
rect 57664 12600 57897 12628
rect 57664 12588 57670 12600
rect 57885 12597 57897 12600
rect 57931 12597 57943 12631
rect 57885 12591 57943 12597
rect 1104 12538 58880 12560
rect 1104 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 22616 12538
rect 22668 12486 22680 12538
rect 22732 12486 22744 12538
rect 22796 12486 22808 12538
rect 22860 12486 22872 12538
rect 22924 12486 37060 12538
rect 37112 12486 37124 12538
rect 37176 12486 37188 12538
rect 37240 12486 37252 12538
rect 37304 12486 37316 12538
rect 37368 12486 51504 12538
rect 51556 12486 51568 12538
rect 51620 12486 51632 12538
rect 51684 12486 51696 12538
rect 51748 12486 51760 12538
rect 51812 12486 58880 12538
rect 1104 12464 58880 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 1912 12396 2237 12424
rect 1912 12384 1918 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 3694 12424 3700 12436
rect 2225 12387 2283 12393
rect 3436 12396 3700 12424
rect 3436 12288 3464 12396
rect 3694 12384 3700 12396
rect 3752 12424 3758 12436
rect 5445 12427 5503 12433
rect 3752 12396 5396 12424
rect 3752 12384 3758 12396
rect 5368 12356 5396 12396
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5534 12424 5540 12436
rect 5491 12396 5540 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6052 12396 10364 12424
rect 6052 12384 6058 12396
rect 10336 12356 10364 12396
rect 10410 12384 10416 12436
rect 10468 12384 10474 12436
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 14424 12396 15025 12424
rect 14424 12384 14430 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 19518 12424 19524 12436
rect 15013 12387 15071 12393
rect 19352 12396 19524 12424
rect 10778 12356 10784 12368
rect 3344 12260 3464 12288
rect 3620 12328 5304 12356
rect 5368 12328 6316 12356
rect 10336 12328 10784 12356
rect 3344 12229 3372 12260
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 2961 12223 3019 12229
rect 2961 12220 2973 12223
rect 2915 12192 2973 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2961 12189 2973 12192
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3620 12220 3648 12328
rect 5166 12288 5172 12300
rect 4172 12260 4568 12288
rect 4172 12232 4200 12260
rect 3467 12192 3648 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3160 12084 3188 12183
rect 3620 12096 3648 12192
rect 4154 12180 4160 12232
rect 4212 12180 4218 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 4264 12192 4353 12220
rect 4264 12096 4292 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4540 12220 4568 12260
rect 5092 12260 5172 12288
rect 5092 12229 5120 12260
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5276 12229 5304 12328
rect 6288 12300 6316 12328
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 12897 12359 12955 12365
rect 12897 12356 12909 12359
rect 12584 12328 12909 12356
rect 12584 12316 12590 12328
rect 12897 12325 12909 12328
rect 12943 12325 12955 12359
rect 12897 12319 12955 12325
rect 14734 12316 14740 12368
rect 14792 12316 14798 12368
rect 6270 12248 6276 12300
rect 6328 12248 6334 12300
rect 11054 12248 11060 12300
rect 11112 12248 11118 12300
rect 11624 12260 12848 12288
rect 4597 12223 4655 12229
rect 4597 12220 4609 12223
rect 4540 12192 4609 12220
rect 4341 12183 4399 12189
rect 4597 12189 4609 12192
rect 4643 12189 4655 12223
rect 4597 12183 4655 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4847 12192 4905 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12220 5319 12223
rect 5626 12220 5632 12232
rect 5307 12192 5632 12220
rect 5307 12189 5319 12192
rect 5261 12183 5319 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 6086 12220 6092 12232
rect 5767 12192 6092 12220
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 8018 12220 8024 12232
rect 6411 12192 8024 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 10183 12192 11161 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 5169 12155 5227 12161
rect 5169 12121 5181 12155
rect 5215 12121 5227 12155
rect 5169 12115 5227 12121
rect 6273 12155 6331 12161
rect 6273 12121 6285 12155
rect 6319 12152 6331 12155
rect 6610 12155 6668 12161
rect 6610 12152 6622 12155
rect 6319 12124 6622 12152
rect 6319 12121 6331 12124
rect 6273 12115 6331 12121
rect 6610 12121 6622 12124
rect 6656 12121 6668 12155
rect 9585 12155 9643 12161
rect 9585 12152 9597 12155
rect 6610 12115 6668 12121
rect 9508 12124 9597 12152
rect 3326 12084 3332 12096
rect 3160 12056 3332 12084
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 3602 12044 3608 12096
rect 3660 12044 3666 12096
rect 4246 12044 4252 12096
rect 4304 12044 4310 12096
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 4522 12084 4528 12096
rect 4479 12056 4528 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 5184 12084 5212 12115
rect 9508 12096 9536 12124
rect 9585 12121 9597 12124
rect 9631 12152 9643 12155
rect 11624 12152 11652 12260
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 9631 12124 11652 12152
rect 9631 12121 9643 12124
rect 9585 12115 9643 12121
rect 7098 12084 7104 12096
rect 5184 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12084 7162 12096
rect 7558 12084 7564 12096
rect 7156 12056 7564 12084
rect 7156 12044 7162 12056
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8812 12056 9229 12084
rect 8812 12044 8818 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 9490 12044 9496 12096
rect 9548 12044 9554 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11716 12084 11744 12183
rect 12820 12164 12848 12260
rect 13354 12248 13360 12300
rect 13412 12248 13418 12300
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13464 12152 13492 12251
rect 14090 12248 14096 12300
rect 14148 12248 14154 12300
rect 19352 12297 19380 12396
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 19981 12427 20039 12433
rect 19981 12393 19993 12427
rect 20027 12424 20039 12427
rect 20806 12424 20812 12436
rect 20027 12396 20812 12424
rect 20027 12393 20039 12396
rect 19981 12387 20039 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 27246 12424 27252 12436
rect 24872 12396 27252 12424
rect 24872 12368 24900 12396
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 27338 12384 27344 12436
rect 27396 12424 27402 12436
rect 27709 12427 27767 12433
rect 27709 12424 27721 12427
rect 27396 12396 27721 12424
rect 27396 12384 27402 12396
rect 27709 12393 27721 12396
rect 27755 12393 27767 12427
rect 27709 12387 27767 12393
rect 31662 12384 31668 12436
rect 31720 12384 31726 12436
rect 34333 12427 34391 12433
rect 34333 12393 34345 12427
rect 34379 12424 34391 12427
rect 34514 12424 34520 12436
rect 34379 12396 34520 12424
rect 34379 12393 34391 12396
rect 34333 12387 34391 12393
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 35158 12384 35164 12436
rect 35216 12424 35222 12436
rect 35345 12427 35403 12433
rect 35345 12424 35357 12427
rect 35216 12396 35357 12424
rect 35216 12384 35222 12396
rect 35345 12393 35357 12396
rect 35391 12393 35403 12427
rect 35345 12387 35403 12393
rect 36814 12384 36820 12436
rect 36872 12384 36878 12436
rect 37645 12427 37703 12433
rect 37645 12393 37657 12427
rect 37691 12424 37703 12427
rect 37734 12424 37740 12436
rect 37691 12396 37740 12424
rect 37691 12393 37703 12396
rect 37645 12387 37703 12393
rect 37734 12384 37740 12396
rect 37792 12384 37798 12436
rect 38102 12384 38108 12436
rect 38160 12424 38166 12436
rect 38565 12427 38623 12433
rect 38565 12424 38577 12427
rect 38160 12396 38577 12424
rect 38160 12384 38166 12396
rect 38565 12393 38577 12396
rect 38611 12393 38623 12427
rect 42150 12424 42156 12436
rect 38565 12387 38623 12393
rect 39040 12396 42156 12424
rect 24854 12356 24860 12368
rect 19444 12328 24860 12356
rect 19337 12291 19395 12297
rect 16132 12260 19288 12288
rect 16022 12152 16028 12164
rect 12860 12124 16028 12152
rect 12860 12112 12866 12124
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11204 12056 12081 12084
rect 11204 12044 11210 12056
rect 12069 12053 12081 12056
rect 12115 12084 12127 12087
rect 16132 12084 16160 12260
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 16850 12220 16856 12232
rect 16531 12192 16856 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 19260 12220 19288 12260
rect 19337 12257 19349 12291
rect 19383 12257 19395 12291
rect 19337 12251 19395 12257
rect 19444 12220 19472 12328
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 27617 12359 27675 12365
rect 27617 12325 27629 12359
rect 27663 12325 27675 12359
rect 27617 12319 27675 12325
rect 21637 12291 21695 12297
rect 21637 12257 21649 12291
rect 21683 12288 21695 12291
rect 22002 12288 22008 12300
rect 21683 12260 22008 12288
rect 21683 12257 21695 12260
rect 21637 12251 21695 12257
rect 22002 12248 22008 12260
rect 22060 12288 22066 12300
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 22060 12260 22385 12288
rect 22060 12248 22066 12260
rect 22373 12257 22385 12260
rect 22419 12257 22431 12291
rect 27632 12288 27660 12319
rect 37550 12316 37556 12368
rect 37608 12356 37614 12368
rect 38930 12356 38936 12368
rect 37608 12328 38936 12356
rect 37608 12316 37614 12328
rect 38930 12316 38936 12328
rect 38988 12316 38994 12368
rect 27798 12288 27804 12300
rect 27632 12260 27804 12288
rect 22373 12251 22431 12257
rect 27798 12248 27804 12260
rect 27856 12288 27862 12300
rect 28261 12291 28319 12297
rect 28261 12288 28273 12291
rect 27856 12260 28273 12288
rect 27856 12248 27862 12260
rect 28261 12257 28273 12260
rect 28307 12257 28319 12291
rect 28261 12251 28319 12257
rect 34698 12248 34704 12300
rect 34756 12248 34762 12300
rect 37458 12248 37464 12300
rect 37516 12248 37522 12300
rect 38286 12248 38292 12300
rect 38344 12248 38350 12300
rect 19260 12192 19472 12220
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19567 12192 20085 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 24026 12180 24032 12232
rect 24084 12180 24090 12232
rect 24946 12180 24952 12232
rect 25004 12180 25010 12232
rect 26237 12223 26295 12229
rect 26237 12189 26249 12223
rect 26283 12220 26295 12223
rect 26283 12192 26648 12220
rect 26283 12189 26295 12192
rect 26237 12183 26295 12189
rect 26620 12164 26648 12192
rect 26970 12180 26976 12232
rect 27028 12180 27034 12232
rect 27062 12180 27068 12232
rect 27120 12220 27126 12232
rect 27120 12192 29684 12220
rect 27120 12180 27126 12192
rect 17129 12155 17187 12161
rect 17129 12121 17141 12155
rect 17175 12152 17187 12155
rect 18690 12152 18696 12164
rect 17175 12124 18696 12152
rect 17175 12121 17187 12124
rect 17129 12115 17187 12121
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 19978 12152 19984 12164
rect 18923 12124 19984 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 19978 12112 19984 12124
rect 20036 12152 20042 12164
rect 21085 12155 21143 12161
rect 21085 12152 21097 12155
rect 20036 12124 21097 12152
rect 20036 12112 20042 12124
rect 21085 12121 21097 12124
rect 21131 12152 21143 12155
rect 22094 12152 22100 12164
rect 21131 12124 22100 12152
rect 21131 12121 21143 12124
rect 21085 12115 21143 12121
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 22189 12155 22247 12161
rect 22189 12121 22201 12155
rect 22235 12152 22247 12155
rect 22235 12124 24348 12152
rect 22235 12121 22247 12124
rect 22189 12115 22247 12121
rect 24320 12096 24348 12124
rect 24486 12112 24492 12164
rect 24544 12152 24550 12164
rect 26510 12161 26516 12164
rect 25593 12155 25651 12161
rect 25593 12152 25605 12155
rect 24544 12124 25605 12152
rect 24544 12112 24550 12124
rect 25593 12121 25605 12124
rect 25639 12152 25651 12155
rect 25639 12124 26004 12152
rect 25639 12121 25651 12124
rect 25593 12115 25651 12121
rect 12115 12056 16160 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19392 12056 19625 12084
rect 19392 12044 19398 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 21818 12044 21824 12096
rect 21876 12044 21882 12096
rect 22278 12044 22284 12096
rect 22336 12044 22342 12096
rect 23474 12044 23480 12096
rect 23532 12044 23538 12096
rect 24302 12044 24308 12096
rect 24360 12044 24366 12096
rect 24394 12044 24400 12096
rect 24452 12044 24458 12096
rect 25866 12044 25872 12096
rect 25924 12044 25930 12096
rect 25976 12084 26004 12124
rect 26504 12115 26516 12161
rect 26510 12112 26516 12115
rect 26568 12112 26574 12164
rect 26602 12112 26608 12164
rect 26660 12112 26666 12164
rect 26988 12084 27016 12180
rect 29546 12112 29552 12164
rect 29604 12112 29610 12164
rect 29656 12152 29684 12192
rect 31018 12180 31024 12232
rect 31076 12220 31082 12232
rect 36170 12220 36176 12232
rect 31076 12192 36176 12220
rect 31076 12180 31082 12192
rect 36170 12180 36176 12192
rect 36228 12180 36234 12232
rect 36262 12180 36268 12232
rect 36320 12180 36326 12232
rect 36722 12180 36728 12232
rect 36780 12220 36786 12232
rect 39040 12220 39068 12396
rect 42150 12384 42156 12396
rect 42208 12384 42214 12436
rect 46842 12384 46848 12436
rect 46900 12384 46906 12436
rect 47026 12384 47032 12436
rect 47084 12384 47090 12436
rect 48498 12384 48504 12436
rect 48556 12384 48562 12436
rect 48590 12384 48596 12436
rect 48648 12424 48654 12436
rect 49329 12427 49387 12433
rect 49329 12424 49341 12427
rect 48648 12396 49341 12424
rect 48648 12384 48654 12396
rect 49329 12393 49341 12396
rect 49375 12424 49387 12427
rect 52454 12424 52460 12436
rect 49375 12396 52460 12424
rect 49375 12393 49387 12396
rect 49329 12387 49387 12393
rect 42613 12359 42671 12365
rect 42613 12325 42625 12359
rect 42659 12356 42671 12359
rect 43898 12356 43904 12368
rect 42659 12328 43904 12356
rect 42659 12325 42671 12328
rect 42613 12319 42671 12325
rect 43898 12316 43904 12328
rect 43956 12356 43962 12368
rect 45741 12359 45799 12365
rect 43956 12328 44220 12356
rect 43956 12316 43962 12328
rect 42518 12248 42524 12300
rect 42576 12288 42582 12300
rect 42702 12288 42708 12300
rect 42576 12260 42708 12288
rect 42576 12248 42582 12260
rect 42702 12248 42708 12260
rect 42760 12288 42766 12300
rect 43257 12291 43315 12297
rect 43257 12288 43269 12291
rect 42760 12260 43269 12288
rect 42760 12248 42766 12260
rect 43257 12257 43269 12260
rect 43303 12288 43315 12291
rect 43990 12288 43996 12300
rect 43303 12260 43996 12288
rect 43303 12257 43315 12260
rect 43257 12251 43315 12257
rect 43990 12248 43996 12260
rect 44048 12248 44054 12300
rect 44192 12297 44220 12328
rect 45741 12325 45753 12359
rect 45787 12356 45799 12359
rect 47044 12356 47072 12384
rect 45787 12328 47072 12356
rect 50157 12359 50215 12365
rect 45787 12325 45799 12328
rect 45741 12319 45799 12325
rect 50157 12325 50169 12359
rect 50203 12356 50215 12359
rect 50430 12356 50436 12368
rect 50203 12328 50436 12356
rect 50203 12325 50215 12328
rect 50157 12319 50215 12325
rect 50430 12316 50436 12328
rect 50488 12316 50494 12368
rect 51552 12300 51580 12396
rect 52454 12384 52460 12396
rect 52512 12424 52518 12436
rect 52549 12427 52607 12433
rect 52549 12424 52561 12427
rect 52512 12396 52561 12424
rect 52512 12384 52518 12396
rect 52549 12393 52561 12396
rect 52595 12424 52607 12427
rect 52917 12427 52975 12433
rect 52917 12424 52929 12427
rect 52595 12396 52929 12424
rect 52595 12393 52607 12396
rect 52549 12387 52607 12393
rect 52917 12393 52929 12396
rect 52963 12393 52975 12427
rect 52917 12387 52975 12393
rect 54110 12384 54116 12436
rect 54168 12424 54174 12436
rect 54294 12424 54300 12436
rect 54168 12396 54300 12424
rect 54168 12384 54174 12396
rect 54294 12384 54300 12396
rect 54352 12384 54358 12436
rect 57238 12384 57244 12436
rect 57296 12384 57302 12436
rect 57149 12359 57207 12365
rect 57149 12325 57161 12359
rect 57195 12325 57207 12359
rect 57149 12319 57207 12325
rect 44177 12291 44235 12297
rect 44177 12257 44189 12291
rect 44223 12257 44235 12291
rect 44177 12251 44235 12257
rect 45097 12291 45155 12297
rect 45097 12257 45109 12291
rect 45143 12257 45155 12291
rect 45097 12251 45155 12257
rect 41230 12220 41236 12232
rect 36780 12192 39068 12220
rect 40420 12192 41236 12220
rect 36780 12180 36786 12192
rect 33137 12155 33195 12161
rect 33137 12152 33149 12155
rect 29656 12124 33149 12152
rect 33137 12121 33149 12124
rect 33183 12152 33195 12155
rect 33318 12152 33324 12164
rect 33183 12124 33324 12152
rect 33183 12121 33195 12124
rect 33137 12115 33195 12121
rect 33318 12112 33324 12124
rect 33376 12112 33382 12164
rect 38102 12112 38108 12164
rect 38160 12152 38166 12164
rect 40310 12152 40316 12164
rect 38160 12124 40316 12152
rect 38160 12112 38166 12124
rect 40310 12112 40316 12124
rect 40368 12152 40374 12164
rect 40420 12161 40448 12192
rect 41230 12180 41236 12192
rect 41288 12180 41294 12232
rect 45112 12220 45140 12251
rect 45462 12248 45468 12300
rect 45520 12288 45526 12300
rect 46109 12291 46167 12297
rect 46109 12288 46121 12291
rect 45520 12260 46121 12288
rect 45520 12248 45526 12260
rect 46109 12257 46121 12260
rect 46155 12288 46167 12291
rect 47210 12288 47216 12300
rect 46155 12260 47216 12288
rect 46155 12257 46167 12260
rect 46109 12251 46167 12257
rect 47210 12248 47216 12260
rect 47268 12248 47274 12300
rect 51534 12248 51540 12300
rect 51592 12248 51598 12300
rect 52178 12248 52184 12300
rect 52236 12248 52242 12300
rect 54478 12248 54484 12300
rect 54536 12288 54542 12300
rect 56505 12291 56563 12297
rect 56505 12288 56517 12291
rect 54536 12260 56517 12288
rect 54536 12248 54542 12260
rect 41386 12192 45140 12220
rect 40405 12155 40463 12161
rect 40405 12152 40417 12155
rect 40368 12124 40417 12152
rect 40368 12112 40374 12124
rect 40405 12121 40417 12124
rect 40451 12121 40463 12155
rect 40405 12115 40463 12121
rect 25976 12056 27016 12084
rect 30650 12044 30656 12096
rect 30708 12084 30714 12096
rect 30837 12087 30895 12093
rect 30837 12084 30849 12087
rect 30708 12056 30849 12084
rect 30708 12044 30714 12056
rect 30837 12053 30849 12056
rect 30883 12053 30895 12087
rect 30837 12047 30895 12053
rect 32030 12044 32036 12096
rect 32088 12044 32094 12096
rect 35710 12044 35716 12096
rect 35768 12044 35774 12096
rect 36446 12044 36452 12096
rect 36504 12084 36510 12096
rect 36630 12084 36636 12096
rect 36504 12056 36636 12084
rect 36504 12044 36510 12056
rect 36630 12044 36636 12056
rect 36688 12044 36694 12096
rect 40129 12087 40187 12093
rect 40129 12053 40141 12087
rect 40175 12084 40187 12087
rect 40218 12084 40224 12096
rect 40175 12056 40224 12084
rect 40175 12053 40187 12056
rect 40129 12047 40187 12053
rect 40218 12044 40224 12056
rect 40276 12084 40282 12096
rect 41386 12084 41414 12192
rect 41500 12155 41558 12161
rect 41500 12121 41512 12155
rect 41546 12152 41558 12155
rect 42426 12152 42432 12164
rect 41546 12124 42432 12152
rect 41546 12121 41558 12124
rect 41500 12115 41558 12121
rect 42426 12112 42432 12124
rect 42484 12112 42490 12164
rect 43073 12155 43131 12161
rect 43073 12121 43085 12155
rect 43119 12152 43131 12155
rect 43533 12155 43591 12161
rect 43533 12152 43545 12155
rect 43119 12124 43545 12152
rect 43119 12121 43131 12124
rect 43073 12115 43131 12121
rect 43533 12121 43545 12124
rect 43579 12121 43591 12155
rect 43533 12115 43591 12121
rect 44545 12155 44603 12161
rect 44545 12121 44557 12155
rect 44591 12152 44603 12155
rect 44634 12152 44640 12164
rect 44591 12124 44640 12152
rect 44591 12121 44603 12124
rect 44545 12115 44603 12121
rect 44634 12112 44640 12124
rect 44692 12112 44698 12164
rect 45112 12152 45140 12192
rect 45186 12180 45192 12232
rect 45244 12220 45250 12232
rect 45373 12223 45431 12229
rect 45373 12220 45385 12223
rect 45244 12192 45385 12220
rect 45244 12180 45250 12192
rect 45373 12189 45385 12192
rect 45419 12189 45431 12223
rect 45373 12183 45431 12189
rect 45554 12180 45560 12232
rect 45612 12220 45618 12232
rect 47394 12220 47400 12232
rect 45612 12192 47400 12220
rect 45612 12180 45618 12192
rect 47394 12180 47400 12192
rect 47452 12180 47458 12232
rect 46385 12155 46443 12161
rect 46385 12152 46397 12155
rect 45112 12124 46397 12152
rect 46385 12121 46397 12124
rect 46431 12121 46443 12155
rect 46385 12115 46443 12121
rect 51292 12155 51350 12161
rect 51292 12121 51304 12155
rect 51338 12152 51350 12155
rect 51338 12124 51488 12152
rect 51338 12121 51350 12124
rect 51292 12115 51350 12121
rect 40276 12056 41414 12084
rect 40276 12044 40282 12056
rect 42702 12044 42708 12096
rect 42760 12044 42766 12096
rect 42886 12044 42892 12096
rect 42944 12084 42950 12096
rect 43165 12087 43223 12093
rect 43165 12084 43177 12087
rect 42944 12056 43177 12084
rect 42944 12044 42950 12056
rect 43165 12053 43177 12056
rect 43211 12084 43223 12087
rect 43806 12084 43812 12096
rect 43211 12056 43812 12084
rect 43211 12053 43223 12056
rect 43165 12047 43223 12053
rect 43806 12044 43812 12056
rect 43864 12084 43870 12096
rect 45281 12087 45339 12093
rect 45281 12084 45293 12087
rect 43864 12056 45293 12084
rect 43864 12044 43870 12056
rect 45281 12053 45293 12056
rect 45327 12053 45339 12087
rect 45281 12047 45339 12053
rect 48774 12044 48780 12096
rect 48832 12084 48838 12096
rect 49418 12084 49424 12096
rect 48832 12056 49424 12084
rect 48832 12044 48838 12056
rect 49418 12044 49424 12056
rect 49476 12044 49482 12096
rect 51460 12084 51488 12124
rect 56244 12096 56272 12260
rect 56505 12257 56517 12260
rect 56551 12257 56563 12291
rect 57164 12288 57192 12319
rect 57793 12291 57851 12297
rect 57793 12288 57805 12291
rect 57164 12260 57805 12288
rect 56505 12251 56563 12257
rect 57793 12257 57805 12260
rect 57839 12257 57851 12291
rect 57793 12251 57851 12257
rect 56689 12223 56747 12229
rect 56689 12189 56701 12223
rect 56735 12220 56747 12223
rect 57606 12220 57612 12232
rect 56735 12192 57612 12220
rect 56735 12189 56747 12192
rect 56689 12183 56747 12189
rect 57606 12180 57612 12192
rect 57664 12180 57670 12232
rect 51629 12087 51687 12093
rect 51629 12084 51641 12087
rect 51460 12056 51641 12084
rect 51629 12053 51641 12056
rect 51675 12053 51687 12087
rect 51629 12047 51687 12053
rect 56226 12044 56232 12096
rect 56284 12044 56290 12096
rect 56778 12044 56784 12096
rect 56836 12084 56842 12096
rect 57606 12084 57612 12096
rect 56836 12056 57612 12084
rect 56836 12044 56842 12056
rect 57606 12044 57612 12056
rect 57664 12044 57670 12096
rect 1104 11994 59040 12016
rect 1104 11942 15394 11994
rect 15446 11942 15458 11994
rect 15510 11942 15522 11994
rect 15574 11942 15586 11994
rect 15638 11942 15650 11994
rect 15702 11942 29838 11994
rect 29890 11942 29902 11994
rect 29954 11942 29966 11994
rect 30018 11942 30030 11994
rect 30082 11942 30094 11994
rect 30146 11942 44282 11994
rect 44334 11942 44346 11994
rect 44398 11942 44410 11994
rect 44462 11942 44474 11994
rect 44526 11942 44538 11994
rect 44590 11942 58726 11994
rect 58778 11942 58790 11994
rect 58842 11942 58854 11994
rect 58906 11942 58918 11994
rect 58970 11942 58982 11994
rect 59034 11942 59040 11994
rect 1104 11920 59040 11942
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4246 11880 4252 11892
rect 4019 11852 4252 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 5169 11883 5227 11889
rect 4580 11852 5028 11880
rect 4580 11840 4586 11852
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 4203 11784 4568 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 3889 11747 3947 11753
rect 3889 11713 3901 11747
rect 3935 11744 3947 11747
rect 4065 11747 4123 11753
rect 3935 11716 4016 11744
rect 3935 11713 3947 11716
rect 3889 11707 3947 11713
rect 3988 11688 4016 11716
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4172 11744 4200 11775
rect 4540 11756 4568 11784
rect 4798 11772 4804 11824
rect 4856 11772 4862 11824
rect 4111 11716 4200 11744
rect 4341 11747 4399 11753
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4356 11676 4384 11707
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 4816 11744 4844 11772
rect 5000 11756 5028 11852
rect 5169 11849 5181 11883
rect 5215 11849 5227 11883
rect 5169 11843 5227 11849
rect 5184 11812 5212 11843
rect 6086 11840 6092 11892
rect 6144 11840 6150 11892
rect 7742 11840 7748 11892
rect 7800 11840 7806 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9732 11852 10548 11880
rect 9732 11840 9738 11852
rect 5721 11815 5779 11821
rect 5721 11812 5733 11815
rect 5184 11784 5733 11812
rect 5721 11781 5733 11784
rect 5767 11781 5779 11815
rect 5721 11775 5779 11781
rect 5813 11815 5871 11821
rect 5813 11781 5825 11815
rect 5859 11812 5871 11815
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 5859 11784 6837 11812
rect 5859 11781 5871 11784
rect 5813 11775 5871 11781
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 7760 11812 7788 11840
rect 6825 11775 6883 11781
rect 7484 11784 7788 11812
rect 10520 11812 10548 11852
rect 11146 11840 11152 11892
rect 11204 11840 11210 11892
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 19978 11880 19984 11892
rect 18187 11852 19984 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 13538 11812 13544 11824
rect 10520 11784 13544 11812
rect 4632 11716 4844 11744
rect 4632 11676 4660 11716
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 4028 11648 4660 11676
rect 4028 11636 4034 11648
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 4816 11608 4844 11639
rect 4356 11580 4844 11608
rect 4356 11552 4384 11580
rect 4908 11552 4936 11639
rect 5552 11552 5580 11707
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5684 11716 5917 11744
rect 5684 11704 5690 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6840 11676 6868 11775
rect 7484 11753 7512 11784
rect 13538 11772 13544 11784
rect 13596 11812 13602 11824
rect 16390 11812 16396 11824
rect 13596 11784 16396 11812
rect 13596 11772 13602 11784
rect 16390 11772 16396 11784
rect 16448 11772 16454 11824
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7558 11704 7564 11756
rect 7616 11704 7622 11756
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9398 11744 9404 11756
rect 9355 11716 9404 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9490 11704 9496 11756
rect 9548 11704 9554 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 9631 11716 9996 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 6840 11648 7665 11676
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 9508 11676 9536 11704
rect 9968 11688 9996 11716
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 18248 11753 18276 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 21818 11840 21824 11892
rect 21876 11840 21882 11892
rect 22278 11880 22284 11892
rect 22066 11852 22284 11880
rect 18500 11815 18558 11821
rect 18500 11781 18512 11815
rect 18546 11812 18558 11815
rect 20254 11812 20260 11824
rect 18546 11784 20260 11812
rect 18546 11781 18558 11784
rect 18500 11775 18558 11781
rect 20254 11772 20260 11784
rect 20312 11772 20318 11824
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16816 11716 17233 11744
rect 16816 11704 16822 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 19426 11744 19432 11756
rect 18380 11716 19432 11744
rect 18380 11704 18386 11716
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 21637 11747 21695 11753
rect 21637 11713 21649 11747
rect 21683 11744 21695 11747
rect 21836 11744 21864 11840
rect 21683 11716 21864 11744
rect 21683 11713 21695 11716
rect 21637 11707 21695 11713
rect 7653 11639 7711 11645
rect 8864 11648 9536 11676
rect 4338 11500 4344 11552
rect 4396 11500 4402 11552
rect 4890 11500 4896 11552
rect 4948 11500 4954 11552
rect 5534 11500 5540 11552
rect 5592 11500 5598 11552
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 6328 11512 7573 11540
rect 6328 11500 6334 11512
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7561 11503 7619 11509
rect 7926 11500 7932 11552
rect 7984 11500 7990 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8864 11549 8892 11648
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14608 11648 15025 11676
rect 14608 11636 14614 11648
rect 15013 11645 15025 11648
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 17310 11636 17316 11688
rect 17368 11636 17374 11688
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 19536 11648 20760 11676
rect 17420 11608 17448 11639
rect 16408 11580 17448 11608
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8076 11512 8861 11540
rect 8076 11500 8082 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8996 11512 9045 11540
rect 8996 11500 9002 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 9306 11500 9312 11552
rect 9364 11500 9370 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 14424 11512 14473 11540
rect 14424 11500 14430 11512
rect 14461 11509 14473 11512
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 16408 11549 16436 11580
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 15160 11512 16405 11540
rect 15160 11500 15166 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 19536 11540 19564 11648
rect 19613 11611 19671 11617
rect 19613 11577 19625 11611
rect 19659 11608 19671 11611
rect 20622 11608 20628 11620
rect 19659 11580 20628 11608
rect 19659 11577 19671 11580
rect 19613 11571 19671 11577
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 20732 11608 20760 11648
rect 20806 11636 20812 11688
rect 20864 11636 20870 11688
rect 21821 11679 21879 11685
rect 21821 11645 21833 11679
rect 21867 11676 21879 11679
rect 22066 11676 22094 11852
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 23474 11840 23480 11892
rect 23532 11840 23538 11892
rect 24026 11840 24032 11892
rect 24084 11840 24090 11892
rect 24394 11840 24400 11892
rect 24452 11880 24458 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 24452 11852 24501 11880
rect 24452 11840 24458 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 24489 11843 24547 11849
rect 25774 11840 25780 11892
rect 25832 11840 25838 11892
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 26973 11883 27031 11889
rect 26973 11880 26985 11883
rect 26568 11852 26985 11880
rect 26568 11840 26574 11852
rect 26973 11849 26985 11852
rect 27019 11849 27031 11883
rect 26973 11843 27031 11849
rect 31110 11840 31116 11892
rect 31168 11840 31174 11892
rect 32766 11840 32772 11892
rect 32824 11880 32830 11892
rect 33502 11880 33508 11892
rect 32824 11852 33508 11880
rect 32824 11840 32830 11852
rect 33502 11840 33508 11852
rect 33560 11840 33566 11892
rect 35897 11883 35955 11889
rect 35897 11849 35909 11883
rect 35943 11880 35955 11883
rect 36262 11880 36268 11892
rect 35943 11852 36268 11880
rect 35943 11849 35955 11852
rect 35897 11843 35955 11849
rect 36262 11840 36268 11852
rect 36320 11840 36326 11892
rect 36357 11883 36415 11889
rect 36357 11849 36369 11883
rect 36403 11880 36415 11883
rect 37093 11883 37151 11889
rect 36403 11852 37044 11880
rect 36403 11849 36415 11852
rect 36357 11843 36415 11849
rect 22824 11815 22882 11821
rect 22824 11781 22836 11815
rect 22870 11812 22882 11815
rect 23492 11812 23520 11840
rect 25792 11812 25820 11840
rect 36722 11812 36728 11824
rect 22870 11784 23520 11812
rect 23584 11784 25820 11812
rect 28920 11784 36728 11812
rect 22870 11781 22882 11784
rect 22824 11775 22882 11781
rect 23584 11744 23612 11784
rect 21867 11648 22094 11676
rect 22204 11716 23612 11744
rect 21867 11645 21879 11648
rect 21821 11639 21879 11645
rect 22204 11608 22232 11716
rect 24302 11704 24308 11756
rect 24360 11744 24366 11756
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 24360 11716 24409 11744
rect 24360 11704 24366 11716
rect 24397 11713 24409 11716
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 27614 11704 27620 11756
rect 27672 11704 27678 11756
rect 28920 11753 28948 11784
rect 36722 11772 36728 11784
rect 36780 11772 36786 11824
rect 28905 11747 28963 11753
rect 28905 11744 28917 11747
rect 28368 11716 28917 11744
rect 22462 11636 22468 11688
rect 22520 11636 22526 11688
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 20732 11580 22232 11608
rect 22278 11568 22284 11620
rect 22336 11608 22342 11620
rect 22572 11608 22600 11639
rect 23566 11636 23572 11688
rect 23624 11676 23630 11688
rect 24578 11676 24584 11688
rect 23624 11648 24584 11676
rect 23624 11636 23630 11648
rect 24578 11636 24584 11648
rect 24636 11636 24642 11688
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25498 11636 25504 11688
rect 25556 11636 25562 11688
rect 22336 11580 22600 11608
rect 22336 11568 22342 11580
rect 16632 11512 19564 11540
rect 16632 11500 16638 11512
rect 20254 11500 20260 11552
rect 20312 11500 20318 11552
rect 20993 11543 21051 11549
rect 20993 11509 21005 11543
rect 21039 11540 21051 11543
rect 21266 11540 21272 11552
rect 21039 11512 21272 11540
rect 21039 11509 21051 11512
rect 20993 11503 21051 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 22572 11540 22600 11580
rect 23937 11611 23995 11617
rect 23937 11577 23949 11611
rect 23983 11608 23995 11611
rect 24964 11608 24992 11636
rect 28368 11617 28396 11716
rect 28905 11713 28917 11716
rect 28951 11713 28963 11747
rect 35342 11744 35348 11756
rect 28905 11707 28963 11713
rect 30576 11716 35348 11744
rect 30576 11688 30604 11716
rect 35342 11704 35348 11716
rect 35400 11744 35406 11756
rect 35713 11747 35771 11753
rect 35713 11744 35725 11747
rect 35400 11716 35725 11744
rect 35400 11704 35406 11716
rect 35713 11713 35725 11716
rect 35759 11713 35771 11747
rect 35713 11707 35771 11713
rect 36265 11747 36323 11753
rect 36265 11713 36277 11747
rect 36311 11744 36323 11747
rect 36311 11716 36768 11744
rect 36311 11713 36323 11716
rect 36265 11707 36323 11713
rect 29086 11636 29092 11688
rect 29144 11676 29150 11688
rect 29273 11679 29331 11685
rect 29273 11676 29285 11679
rect 29144 11648 29285 11676
rect 29144 11636 29150 11648
rect 29273 11645 29285 11648
rect 29319 11676 29331 11679
rect 30558 11676 30564 11688
rect 29319 11648 30564 11676
rect 29319 11645 29331 11648
rect 29273 11639 29331 11645
rect 30558 11636 30564 11648
rect 30616 11636 30622 11688
rect 30653 11679 30711 11685
rect 30653 11645 30665 11679
rect 30699 11676 30711 11679
rect 30926 11676 30932 11688
rect 30699 11648 30932 11676
rect 30699 11645 30711 11648
rect 30653 11639 30711 11645
rect 30926 11636 30932 11648
rect 30984 11636 30990 11688
rect 33134 11636 33140 11688
rect 33192 11636 33198 11688
rect 34422 11636 34428 11688
rect 34480 11636 34486 11688
rect 35728 11676 35756 11707
rect 36449 11679 36507 11685
rect 36449 11676 36461 11679
rect 35728 11648 36461 11676
rect 36449 11645 36461 11648
rect 36495 11676 36507 11679
rect 36538 11676 36544 11688
rect 36495 11648 36544 11676
rect 36495 11645 36507 11648
rect 36449 11639 36507 11645
rect 36538 11636 36544 11648
rect 36596 11636 36602 11688
rect 28353 11611 28411 11617
rect 28353 11608 28365 11611
rect 23983 11580 24992 11608
rect 26068 11580 28365 11608
rect 23983 11577 23995 11580
rect 23937 11571 23995 11577
rect 23198 11540 23204 11552
rect 22572 11512 23204 11540
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 23658 11500 23664 11552
rect 23716 11540 23722 11552
rect 26068 11540 26096 11580
rect 28353 11577 28365 11580
rect 28399 11577 28411 11611
rect 31018 11608 31024 11620
rect 28353 11571 28411 11577
rect 29012 11580 31024 11608
rect 29012 11552 29040 11580
rect 31018 11568 31024 11580
rect 31076 11568 31082 11620
rect 32398 11568 32404 11620
rect 32456 11608 32462 11620
rect 36740 11608 36768 11716
rect 37016 11676 37044 11852
rect 37093 11849 37105 11883
rect 37139 11880 37151 11883
rect 37642 11880 37648 11892
rect 37139 11852 37648 11880
rect 37139 11849 37151 11852
rect 37093 11843 37151 11849
rect 37642 11840 37648 11852
rect 37700 11840 37706 11892
rect 38010 11840 38016 11892
rect 38068 11880 38074 11892
rect 38197 11883 38255 11889
rect 38197 11880 38209 11883
rect 38068 11852 38209 11880
rect 38068 11840 38074 11852
rect 38197 11849 38209 11852
rect 38243 11849 38255 11883
rect 38197 11843 38255 11849
rect 39114 11840 39120 11892
rect 39172 11840 39178 11892
rect 39574 11840 39580 11892
rect 39632 11840 39638 11892
rect 39666 11840 39672 11892
rect 39724 11840 39730 11892
rect 42426 11840 42432 11892
rect 42484 11840 42490 11892
rect 42702 11840 42708 11892
rect 42760 11840 42766 11892
rect 43990 11840 43996 11892
rect 44048 11880 44054 11892
rect 46934 11880 46940 11892
rect 44048 11852 46940 11880
rect 44048 11840 44054 11852
rect 46934 11840 46940 11852
rect 46992 11840 46998 11892
rect 51534 11840 51540 11892
rect 51592 11880 51598 11892
rect 51629 11883 51687 11889
rect 51629 11880 51641 11883
rect 51592 11852 51641 11880
rect 51592 11840 51598 11852
rect 51629 11849 51641 11852
rect 51675 11849 51687 11883
rect 51629 11843 51687 11849
rect 54570 11840 54576 11892
rect 54628 11880 54634 11892
rect 55122 11880 55128 11892
rect 54628 11852 55128 11880
rect 54628 11840 54634 11852
rect 55122 11840 55128 11852
rect 55180 11840 55186 11892
rect 37458 11676 37464 11688
rect 37016 11648 37464 11676
rect 37458 11636 37464 11648
rect 37516 11636 37522 11688
rect 37642 11636 37648 11688
rect 37700 11676 37706 11688
rect 37829 11679 37887 11685
rect 37829 11676 37841 11679
rect 37700 11648 37841 11676
rect 37700 11636 37706 11648
rect 37829 11645 37841 11648
rect 37875 11676 37887 11679
rect 38286 11676 38292 11688
rect 37875 11648 38292 11676
rect 37875 11645 37887 11648
rect 37829 11639 37887 11645
rect 38286 11636 38292 11648
rect 38344 11636 38350 11688
rect 39132 11676 39160 11840
rect 39592 11812 39620 11840
rect 42153 11815 42211 11821
rect 42153 11812 42165 11815
rect 39592 11784 42165 11812
rect 42153 11781 42165 11784
rect 42199 11812 42211 11815
rect 42518 11812 42524 11824
rect 42199 11784 42524 11812
rect 42199 11781 42211 11784
rect 42153 11775 42211 11781
rect 42518 11772 42524 11784
rect 42576 11772 42582 11824
rect 42720 11744 42748 11840
rect 43257 11815 43315 11821
rect 43257 11781 43269 11815
rect 43303 11812 43315 11815
rect 44174 11812 44180 11824
rect 43303 11784 44180 11812
rect 43303 11781 43315 11784
rect 43257 11775 43315 11781
rect 44174 11772 44180 11784
rect 44232 11772 44238 11824
rect 42981 11747 43039 11753
rect 42981 11744 42993 11747
rect 42720 11716 42993 11744
rect 42981 11713 42993 11716
rect 43027 11713 43039 11747
rect 42981 11707 43039 11713
rect 49970 11704 49976 11756
rect 50028 11744 50034 11756
rect 54113 11747 54171 11753
rect 54113 11744 54125 11747
rect 50028 11716 54125 11744
rect 50028 11704 50034 11716
rect 54113 11713 54125 11716
rect 54159 11744 54171 11747
rect 55214 11744 55220 11756
rect 54159 11716 55220 11744
rect 54159 11713 54171 11716
rect 54113 11707 54171 11713
rect 55214 11704 55220 11716
rect 55272 11704 55278 11756
rect 39393 11679 39451 11685
rect 39393 11676 39405 11679
rect 39132 11648 39405 11676
rect 39393 11645 39405 11648
rect 39439 11645 39451 11679
rect 39393 11639 39451 11645
rect 39577 11679 39635 11685
rect 39577 11645 39589 11679
rect 39623 11645 39635 11679
rect 39577 11639 39635 11645
rect 37277 11611 37335 11617
rect 37277 11608 37289 11611
rect 32456 11580 35848 11608
rect 36740 11580 37289 11608
rect 32456 11568 32462 11580
rect 23716 11512 26096 11540
rect 23716 11500 23722 11512
rect 26142 11500 26148 11552
rect 26200 11500 26206 11552
rect 26513 11543 26571 11549
rect 26513 11509 26525 11543
rect 26559 11540 26571 11543
rect 26602 11540 26608 11552
rect 26559 11512 26608 11540
rect 26559 11509 26571 11512
rect 26513 11503 26571 11509
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 28813 11543 28871 11549
rect 28813 11509 28825 11543
rect 28859 11540 28871 11543
rect 28994 11540 29000 11552
rect 28859 11512 29000 11540
rect 28859 11509 28871 11512
rect 28813 11503 28871 11509
rect 28994 11500 29000 11512
rect 29052 11500 29058 11552
rect 29454 11500 29460 11552
rect 29512 11540 29518 11552
rect 30009 11543 30067 11549
rect 30009 11540 30021 11543
rect 29512 11512 30021 11540
rect 29512 11500 29518 11512
rect 30009 11509 30021 11512
rect 30055 11509 30067 11543
rect 30009 11503 30067 11509
rect 33778 11500 33784 11552
rect 33836 11500 33842 11552
rect 33870 11500 33876 11552
rect 33928 11500 33934 11552
rect 35820 11540 35848 11580
rect 37277 11577 37289 11580
rect 37323 11577 37335 11611
rect 37277 11571 37335 11577
rect 37550 11568 37556 11620
rect 37608 11608 37614 11620
rect 39592 11608 39620 11639
rect 45094 11636 45100 11688
rect 45152 11636 45158 11688
rect 45646 11636 45652 11688
rect 45704 11636 45710 11688
rect 48406 11636 48412 11688
rect 48464 11676 48470 11688
rect 49602 11676 49608 11688
rect 48464 11648 49608 11676
rect 48464 11636 48470 11648
rect 49602 11636 49608 11648
rect 49660 11636 49666 11688
rect 50798 11636 50804 11688
rect 50856 11676 50862 11688
rect 51261 11679 51319 11685
rect 51261 11676 51273 11679
rect 50856 11648 51273 11676
rect 50856 11636 50862 11648
rect 51261 11645 51273 11648
rect 51307 11645 51319 11679
rect 51261 11639 51319 11645
rect 57146 11636 57152 11688
rect 57204 11636 57210 11688
rect 43622 11608 43628 11620
rect 37608 11580 39620 11608
rect 39684 11580 43628 11608
rect 37608 11568 37614 11580
rect 39684 11540 39712 11580
rect 43622 11568 43628 11580
rect 43680 11568 43686 11620
rect 43714 11568 43720 11620
rect 43772 11608 43778 11620
rect 44545 11611 44603 11617
rect 44545 11608 44557 11611
rect 43772 11580 44557 11608
rect 43772 11568 43778 11580
rect 44545 11577 44557 11580
rect 44591 11608 44603 11611
rect 44634 11608 44640 11620
rect 44591 11580 44640 11608
rect 44591 11577 44603 11580
rect 44545 11571 44603 11577
rect 44634 11568 44640 11580
rect 44692 11568 44698 11620
rect 50540 11580 51074 11608
rect 35820 11512 39712 11540
rect 40037 11543 40095 11549
rect 40037 11509 40049 11543
rect 40083 11540 40095 11543
rect 41506 11540 41512 11552
rect 40083 11512 41512 11540
rect 40083 11509 40095 11512
rect 40037 11503 40095 11509
rect 41506 11500 41512 11512
rect 41564 11500 41570 11552
rect 43254 11500 43260 11552
rect 43312 11540 43318 11552
rect 47118 11540 47124 11552
rect 43312 11512 47124 11540
rect 43312 11500 43318 11512
rect 47118 11500 47124 11512
rect 47176 11500 47182 11552
rect 47762 11500 47768 11552
rect 47820 11500 47826 11552
rect 50540 11549 50568 11580
rect 50249 11543 50307 11549
rect 50249 11509 50261 11543
rect 50295 11540 50307 11543
rect 50525 11543 50583 11549
rect 50525 11540 50537 11543
rect 50295 11512 50537 11540
rect 50295 11509 50307 11512
rect 50249 11503 50307 11509
rect 50525 11509 50537 11512
rect 50571 11509 50583 11543
rect 50525 11503 50583 11509
rect 50706 11500 50712 11552
rect 50764 11500 50770 11552
rect 51046 11540 51074 11580
rect 51258 11540 51264 11552
rect 51046 11512 51264 11540
rect 51258 11500 51264 11512
rect 51316 11500 51322 11552
rect 56594 11500 56600 11552
rect 56652 11500 56658 11552
rect 1104 11450 58880 11472
rect 1104 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 22616 11450
rect 22668 11398 22680 11450
rect 22732 11398 22744 11450
rect 22796 11398 22808 11450
rect 22860 11398 22872 11450
rect 22924 11398 37060 11450
rect 37112 11398 37124 11450
rect 37176 11398 37188 11450
rect 37240 11398 37252 11450
rect 37304 11398 37316 11450
rect 37368 11398 51504 11450
rect 51556 11398 51568 11450
rect 51620 11398 51632 11450
rect 51684 11398 51696 11450
rect 51748 11398 51760 11450
rect 51812 11398 58880 11450
rect 1104 11376 58880 11398
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 3436 11268 3464 11299
rect 3602 11296 3608 11348
rect 3660 11296 3666 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 3988 11268 4016 11299
rect 4154 11296 4160 11348
rect 4212 11296 4218 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4396 11308 4660 11336
rect 4396 11296 4402 11308
rect 3436 11240 4292 11268
rect 4264 11200 4292 11240
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4264 11172 4537 11200
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4632 11200 4660 11308
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 9306 11296 9312 11348
rect 9364 11296 9370 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 9916 11308 11529 11336
rect 9916 11296 9922 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 11940 11308 12173 11336
rect 11940 11296 11946 11308
rect 12161 11305 12173 11308
rect 12207 11336 12219 11339
rect 12802 11336 12808 11348
rect 12207 11308 12808 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13504 11308 13737 11336
rect 13504 11296 13510 11308
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 17368 11308 18429 11336
rect 17368 11296 17374 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18417 11299 18475 11305
rect 19429 11339 19487 11345
rect 19429 11305 19441 11339
rect 19475 11336 19487 11339
rect 19518 11336 19524 11348
rect 19475 11308 19524 11336
rect 19475 11305 19487 11308
rect 19429 11299 19487 11305
rect 19518 11296 19524 11308
rect 19576 11336 19582 11348
rect 20346 11336 20352 11348
rect 19576 11308 20352 11336
rect 19576 11296 19582 11308
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 22094 11336 22100 11348
rect 21192 11308 22100 11336
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 4632 11172 5641 11200
rect 4525 11163 4583 11169
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 9324 11200 9352 11296
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10597 11271 10655 11277
rect 10597 11268 10609 11271
rect 10100 11240 10609 11268
rect 10100 11228 10106 11240
rect 10597 11237 10609 11240
rect 10643 11237 10655 11271
rect 10597 11231 10655 11237
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 13541 11271 13599 11277
rect 13541 11268 13553 11271
rect 10836 11240 13553 11268
rect 10836 11228 10842 11240
rect 13541 11237 13553 11240
rect 13587 11268 13599 11271
rect 14090 11268 14096 11280
rect 13587 11240 14096 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11237 15531 11271
rect 15473 11231 15531 11237
rect 15488 11200 15516 11231
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 8812 11172 8984 11200
rect 9324 11172 11560 11200
rect 8812 11160 8818 11172
rect 3326 11092 3332 11144
rect 3384 11092 3390 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4057 11137 4115 11143
rect 4057 11134 4069 11137
rect 3988 11132 4069 11134
rect 3936 11106 4069 11132
rect 3936 11104 4016 11106
rect 3936 11092 3942 11104
rect 4057 11103 4069 11106
rect 4103 11103 4115 11137
rect 4057 11097 4115 11103
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4488 11104 4629 11132
rect 4488 11092 4494 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4755 11104 4844 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 3234 11024 3240 11076
rect 3292 11024 3298 11076
rect 3344 10996 3372 11092
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 3970 11064 3976 11076
rect 3651 11036 3976 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4356 11064 4384 11092
rect 4816 11076 4844 11104
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 8956 11141 8984 11172
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 5040 11104 5273 11132
rect 5040 11092 5046 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9674 11132 9680 11144
rect 9447 11104 9680 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10183 11104 10517 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 10505 11101 10517 11104
rect 10551 11132 10563 11135
rect 10551 11104 11192 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 4172 11036 4384 11064
rect 4172 10996 4200 11036
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 4908 11064 4936 11092
rect 8021 11067 8079 11073
rect 4908 11036 5488 11064
rect 3344 10968 4200 10996
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4706 10996 4712 11008
rect 4304 10968 4712 10996
rect 4304 10956 4310 10968
rect 4706 10956 4712 10968
rect 4764 10996 4770 11008
rect 5460 11005 5488 11036
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8757 11067 8815 11073
rect 8067 11036 8708 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 5353 10999 5411 11005
rect 5353 10996 5365 10999
rect 4764 10968 5365 10996
rect 4764 10956 4770 10968
rect 5353 10965 5365 10968
rect 5399 10965 5411 10999
rect 5353 10959 5411 10965
rect 5445 10999 5503 11005
rect 5445 10965 5457 10999
rect 5491 10996 5503 10999
rect 5626 10996 5632 11008
rect 5491 10968 5632 10996
rect 5491 10965 5503 10968
rect 5445 10959 5503 10965
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 8680 10996 8708 11036
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 9214 11064 9220 11076
rect 8803 11036 9220 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 11164 11073 11192 11104
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11532 11141 11560 11172
rect 11716 11172 14228 11200
rect 15488 11172 16129 11200
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 9916 11036 10793 11064
rect 9916 11024 9922 11036
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 11149 11067 11207 11073
rect 11149 11033 11161 11067
rect 11195 11064 11207 11067
rect 11716 11064 11744 11172
rect 11790 11092 11796 11144
rect 11848 11092 11854 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13964 11104 14105 11132
rect 13964 11092 13970 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14200 11132 14228 11172
rect 16117 11169 16129 11172
rect 16163 11200 16175 11203
rect 16482 11200 16488 11212
rect 16163 11172 16488 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 19610 11200 19616 11212
rect 18371 11172 19616 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 16592 11132 16620 11160
rect 14200 11104 16620 11132
rect 14093 11095 14151 11101
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16724 11104 16865 11132
rect 16724 11092 16730 11104
rect 16853 11101 16865 11104
rect 16899 11132 16911 11135
rect 18340 11132 18368 11163
rect 19610 11160 19616 11172
rect 19668 11200 19674 11212
rect 21192 11209 21220 11308
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 23293 11339 23351 11345
rect 23293 11305 23305 11339
rect 23339 11336 23351 11339
rect 24486 11336 24492 11348
rect 23339 11308 24492 11336
rect 23339 11305 23351 11308
rect 23293 11299 23351 11305
rect 24486 11296 24492 11308
rect 24544 11296 24550 11348
rect 24762 11296 24768 11348
rect 24820 11336 24826 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 24820 11308 25237 11336
rect 24820 11296 24826 11308
rect 25225 11305 25237 11308
rect 25271 11336 25283 11339
rect 25271 11308 27292 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 22462 11228 22468 11280
rect 22520 11268 22526 11280
rect 22557 11271 22615 11277
rect 22557 11268 22569 11271
rect 22520 11240 22569 11268
rect 22520 11228 22526 11240
rect 22557 11237 22569 11240
rect 22603 11268 22615 11271
rect 22603 11240 23980 11268
rect 22603 11237 22615 11240
rect 22557 11231 22615 11237
rect 23952 11212 23980 11240
rect 21177 11203 21235 11209
rect 19668 11172 19748 11200
rect 19668 11160 19674 11172
rect 16899 11104 18368 11132
rect 16899 11101 16911 11104
rect 16853 11095 16911 11101
rect 18966 11092 18972 11144
rect 19024 11092 19030 11144
rect 19720 11141 19748 11172
rect 21177 11169 21189 11203
rect 21223 11169 21235 11203
rect 21177 11163 21235 11169
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 21192 11132 21220 11163
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 23845 11203 23903 11209
rect 23845 11200 23857 11203
rect 23624 11172 23857 11200
rect 23624 11160 23630 11172
rect 23845 11169 23857 11172
rect 23891 11169 23903 11203
rect 23845 11163 23903 11169
rect 23934 11160 23940 11212
rect 23992 11160 23998 11212
rect 26602 11160 26608 11212
rect 26660 11160 26666 11212
rect 27264 11209 27292 11308
rect 29454 11296 29460 11348
rect 29512 11296 29518 11348
rect 30926 11296 30932 11348
rect 30984 11296 30990 11348
rect 33318 11296 33324 11348
rect 33376 11296 33382 11348
rect 37366 11296 37372 11348
rect 37424 11336 37430 11348
rect 37461 11339 37519 11345
rect 37461 11336 37473 11339
rect 37424 11308 37473 11336
rect 37424 11296 37430 11308
rect 37461 11305 37473 11308
rect 37507 11336 37519 11339
rect 38102 11336 38108 11348
rect 37507 11308 38108 11336
rect 37507 11305 37519 11308
rect 37461 11299 37519 11305
rect 38102 11296 38108 11308
rect 38160 11296 38166 11348
rect 38470 11296 38476 11348
rect 38528 11336 38534 11348
rect 38528 11308 38792 11336
rect 38528 11296 38534 11308
rect 28994 11268 29000 11280
rect 28828 11240 29000 11268
rect 28828 11209 28856 11240
rect 28994 11228 29000 11240
rect 29052 11228 29058 11280
rect 27249 11203 27307 11209
rect 27249 11169 27261 11203
rect 27295 11169 27307 11203
rect 27249 11163 27307 11169
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11169 28871 11203
rect 28813 11163 28871 11169
rect 28905 11203 28963 11209
rect 28905 11169 28917 11203
rect 28951 11200 28963 11203
rect 29472 11200 29500 11296
rect 28951 11172 29500 11200
rect 28951 11169 28963 11172
rect 28905 11163 28963 11169
rect 19751 11104 21220 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 21433 11135 21491 11141
rect 21433 11132 21445 11135
rect 21324 11104 21445 11132
rect 21324 11092 21330 11104
rect 21433 11101 21445 11104
rect 21479 11101 21491 11135
rect 21433 11095 21491 11101
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11132 22983 11135
rect 23198 11132 23204 11144
rect 22971 11104 23204 11132
rect 22971 11101 22983 11104
rect 22925 11095 22983 11101
rect 23198 11092 23204 11104
rect 23256 11132 23262 11144
rect 25133 11135 25191 11141
rect 25133 11132 25145 11135
rect 23256 11104 25145 11132
rect 23256 11092 23262 11104
rect 25133 11101 25145 11104
rect 25179 11132 25191 11135
rect 26620 11132 26648 11160
rect 25179 11104 26648 11132
rect 25179 11101 25191 11104
rect 25133 11095 25191 11101
rect 28534 11092 28540 11144
rect 28592 11092 28598 11144
rect 29549 11135 29607 11141
rect 29549 11101 29561 11135
rect 29595 11101 29607 11135
rect 29549 11095 29607 11101
rect 11195 11036 11744 11064
rect 13817 11067 13875 11073
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 13817 11033 13829 11067
rect 13863 11064 13875 11067
rect 14182 11064 14188 11076
rect 13863 11036 14188 11064
rect 13863 11033 13875 11036
rect 13817 11027 13875 11033
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 14366 11073 14372 11076
rect 14349 11067 14372 11073
rect 14349 11033 14361 11067
rect 14349 11027 14372 11033
rect 14366 11024 14372 11027
rect 14424 11024 14430 11076
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15565 11067 15623 11073
rect 15565 11064 15577 11067
rect 15344 11036 15577 11064
rect 15344 11024 15350 11036
rect 15565 11033 15577 11036
rect 15611 11033 15623 11067
rect 15565 11027 15623 11033
rect 18046 11024 18052 11076
rect 18104 11073 18110 11076
rect 18104 11027 18116 11073
rect 19972 11067 20030 11073
rect 19972 11033 19984 11067
rect 20018 11064 20030 11067
rect 20254 11064 20260 11076
rect 20018 11036 20260 11064
rect 20018 11033 20030 11036
rect 19972 11027 20030 11033
rect 18104 11024 18110 11027
rect 20254 11024 20260 11036
rect 20312 11024 20318 11076
rect 22462 11064 22468 11076
rect 21100 11036 22468 11064
rect 8846 10996 8852 11008
rect 8680 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9030 10956 9036 11008
rect 9088 10956 9094 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 11514 10996 11520 11008
rect 9456 10968 11520 10996
rect 9456 10956 9462 10968
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 11882 10996 11888 11008
rect 11747 10968 11888 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 16945 10999 17003 11005
rect 16945 10965 16957 10999
rect 16991 10996 17003 10999
rect 17218 10996 17224 11008
rect 16991 10968 17224 10996
rect 16991 10965 17003 10968
rect 16945 10959 17003 10965
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 20714 10996 20720 11008
rect 17644 10968 20720 10996
rect 17644 10956 17650 10968
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 21100 11005 21128 11036
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 23658 11064 23664 11076
rect 23124 11036 23664 11064
rect 21085 10999 21143 11005
rect 21085 10965 21097 10999
rect 21131 10965 21143 10999
rect 21085 10959 21143 10965
rect 21542 10956 21548 11008
rect 21600 10996 21606 11008
rect 23124 10996 23152 11036
rect 23658 11024 23664 11036
rect 23716 11024 23722 11076
rect 26142 11024 26148 11076
rect 26200 11064 26206 11076
rect 26338 11067 26396 11073
rect 26338 11064 26350 11067
rect 26200 11036 26350 11064
rect 26200 11024 26206 11036
rect 26338 11033 26350 11036
rect 26384 11033 26396 11067
rect 29564 11064 29592 11095
rect 31110 11092 31116 11144
rect 31168 11132 31174 11144
rect 31205 11135 31263 11141
rect 31205 11132 31217 11135
rect 31168 11104 31217 11132
rect 31168 11092 31174 11104
rect 31205 11101 31217 11104
rect 31251 11101 31263 11135
rect 31205 11095 31263 11101
rect 32398 11092 32404 11144
rect 32456 11092 32462 11144
rect 33336 11141 33364 11296
rect 36265 11271 36323 11277
rect 36265 11237 36277 11271
rect 36311 11268 36323 11271
rect 36722 11268 36728 11280
rect 36311 11240 36728 11268
rect 36311 11237 36323 11240
rect 36265 11231 36323 11237
rect 36722 11228 36728 11240
rect 36780 11268 36786 11280
rect 36780 11240 37504 11268
rect 36780 11228 36786 11240
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34572 11172 34897 11200
rect 34572 11160 34578 11172
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 34885 11163 34943 11169
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11101 33379 11135
rect 34900 11132 34928 11163
rect 36170 11160 36176 11212
rect 36228 11200 36234 11212
rect 36906 11200 36912 11212
rect 36228 11172 36912 11200
rect 36228 11160 36234 11172
rect 36906 11160 36912 11172
rect 36964 11160 36970 11212
rect 37476 11200 37504 11240
rect 37550 11228 37556 11280
rect 37608 11228 37614 11280
rect 38764 11277 38792 11308
rect 40770 11296 40776 11348
rect 40828 11336 40834 11348
rect 43717 11339 43775 11345
rect 43717 11336 43729 11339
rect 40828 11308 43729 11336
rect 40828 11296 40834 11308
rect 43717 11305 43729 11308
rect 43763 11336 43775 11339
rect 44174 11336 44180 11348
rect 43763 11308 44180 11336
rect 43763 11305 43775 11308
rect 43717 11299 43775 11305
rect 44174 11296 44180 11308
rect 44232 11296 44238 11348
rect 45094 11336 45100 11348
rect 44284 11308 45100 11336
rect 38749 11271 38807 11277
rect 38749 11237 38761 11271
rect 38795 11237 38807 11271
rect 42613 11271 42671 11277
rect 42613 11268 42625 11271
rect 38749 11231 38807 11237
rect 41984 11240 42625 11268
rect 37476 11172 37688 11200
rect 37366 11132 37372 11144
rect 34900 11104 37372 11132
rect 33321 11095 33379 11101
rect 37366 11092 37372 11104
rect 37424 11092 37430 11144
rect 37458 11092 37464 11144
rect 37516 11092 37522 11144
rect 26338 11027 26396 11033
rect 27724 11036 29592 11064
rect 29816 11067 29874 11073
rect 21600 10968 23152 10996
rect 21600 10956 21606 10968
rect 26694 10956 26700 11008
rect 26752 10956 26758 11008
rect 27614 10956 27620 11008
rect 27672 10996 27678 11008
rect 27724 11005 27752 11036
rect 29816 11033 29828 11067
rect 29862 11033 29874 11067
rect 29816 11027 29874 11033
rect 27709 10999 27767 11005
rect 27709 10996 27721 10999
rect 27672 10968 27721 10996
rect 27672 10956 27678 10968
rect 27709 10965 27721 10968
rect 27755 10965 27767 10999
rect 27709 10959 27767 10965
rect 27890 10956 27896 11008
rect 27948 10956 27954 11008
rect 28810 10956 28816 11008
rect 28868 10996 28874 11008
rect 28997 10999 29055 11005
rect 28997 10996 29009 10999
rect 28868 10968 29009 10996
rect 28868 10956 28874 10968
rect 28997 10965 29009 10968
rect 29043 10965 29055 10999
rect 28997 10959 29055 10965
rect 29362 10956 29368 11008
rect 29420 10956 29426 11008
rect 29730 10956 29736 11008
rect 29788 10996 29794 11008
rect 29840 10996 29868 11027
rect 30558 11024 30564 11076
rect 30616 11064 30622 11076
rect 31941 11067 31999 11073
rect 31941 11064 31953 11067
rect 30616 11036 31953 11064
rect 30616 11024 30622 11036
rect 31941 11033 31953 11036
rect 31987 11064 31999 11067
rect 32030 11064 32036 11076
rect 31987 11036 32036 11064
rect 31987 11033 31999 11036
rect 31941 11027 31999 11033
rect 32030 11024 32036 11036
rect 32088 11024 32094 11076
rect 33045 11067 33103 11073
rect 33045 11033 33057 11067
rect 33091 11033 33103 11067
rect 33045 11027 33103 11033
rect 29788 10968 29868 10996
rect 33060 10996 33088 11027
rect 34146 11024 34152 11076
rect 34204 11064 34210 11076
rect 34882 11064 34888 11076
rect 34204 11036 34888 11064
rect 34204 11024 34210 11036
rect 34882 11024 34888 11036
rect 34940 11024 34946 11076
rect 35152 11067 35210 11073
rect 35152 11033 35164 11067
rect 35198 11064 35210 11067
rect 35802 11064 35808 11076
rect 35198 11036 35808 11064
rect 35198 11033 35210 11036
rect 35152 11027 35210 11033
rect 35802 11024 35808 11036
rect 35860 11024 35866 11076
rect 36725 11067 36783 11073
rect 36725 11033 36737 11067
rect 36771 11064 36783 11067
rect 37476 11064 37504 11092
rect 36771 11036 37504 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 34606 10996 34612 11008
rect 33060 10968 34612 10996
rect 29788 10956 29794 10968
rect 34606 10956 34612 10968
rect 34664 10956 34670 11008
rect 36354 10956 36360 11008
rect 36412 10956 36418 11008
rect 36814 10956 36820 11008
rect 36872 10956 36878 11008
rect 37660 10996 37688 11172
rect 38010 11160 38016 11212
rect 38068 11200 38074 11212
rect 38378 11209 38384 11212
rect 38197 11203 38255 11209
rect 38197 11200 38209 11203
rect 38068 11172 38209 11200
rect 38068 11160 38074 11172
rect 38197 11169 38209 11172
rect 38243 11169 38255 11203
rect 38197 11163 38255 11169
rect 38356 11203 38384 11209
rect 38356 11169 38368 11203
rect 38356 11163 38384 11169
rect 38378 11160 38384 11163
rect 38436 11160 38442 11212
rect 39206 11160 39212 11212
rect 39264 11200 39270 11212
rect 41984 11209 42012 11240
rect 42613 11237 42625 11240
rect 42659 11237 42671 11271
rect 43254 11268 43260 11280
rect 42613 11231 42671 11237
rect 43180 11240 43260 11268
rect 43180 11209 43208 11240
rect 43254 11228 43260 11240
rect 43312 11228 43318 11280
rect 43622 11228 43628 11280
rect 43680 11228 43686 11280
rect 40405 11203 40463 11209
rect 40405 11200 40417 11203
rect 39264 11172 40417 11200
rect 39264 11160 39270 11172
rect 40405 11169 40417 11172
rect 40451 11169 40463 11203
rect 40405 11163 40463 11169
rect 41969 11203 42027 11209
rect 41969 11169 41981 11203
rect 42015 11169 42027 11203
rect 43165 11203 43223 11209
rect 43165 11200 43177 11203
rect 41969 11163 42027 11169
rect 42904 11172 43177 11200
rect 38470 11092 38476 11144
rect 38528 11092 38534 11144
rect 39393 11135 39451 11141
rect 39393 11101 39405 11135
rect 39439 11132 39451 11135
rect 39850 11132 39856 11144
rect 39439 11104 39856 11132
rect 39439 11101 39451 11104
rect 39393 11095 39451 11101
rect 39850 11092 39856 11104
rect 39908 11092 39914 11144
rect 41785 11135 41843 11141
rect 41785 11101 41797 11135
rect 41831 11132 41843 11135
rect 42904 11132 42932 11172
rect 43165 11169 43177 11172
rect 43211 11169 43223 11203
rect 43640 11200 43668 11228
rect 44284 11209 44312 11308
rect 45094 11296 45100 11308
rect 45152 11296 45158 11348
rect 50706 11296 50712 11348
rect 50764 11296 50770 11348
rect 50893 11339 50951 11345
rect 50893 11305 50905 11339
rect 50939 11336 50951 11339
rect 52917 11339 52975 11345
rect 50939 11308 51856 11336
rect 50939 11305 50951 11308
rect 50893 11299 50951 11305
rect 44729 11271 44787 11277
rect 44729 11237 44741 11271
rect 44775 11268 44787 11271
rect 47857 11271 47915 11277
rect 44775 11240 46336 11268
rect 44775 11237 44787 11240
rect 44729 11231 44787 11237
rect 44177 11203 44235 11209
rect 44177 11200 44189 11203
rect 43640 11172 44189 11200
rect 43165 11163 43223 11169
rect 44177 11169 44189 11172
rect 44223 11169 44235 11203
rect 44177 11163 44235 11169
rect 44269 11203 44327 11209
rect 44269 11169 44281 11203
rect 44315 11169 44327 11203
rect 45830 11200 45836 11212
rect 44269 11163 44327 11169
rect 44560 11172 45836 11200
rect 41831 11104 42932 11132
rect 43073 11135 43131 11141
rect 41831 11101 41843 11104
rect 41785 11095 41843 11101
rect 43073 11101 43085 11135
rect 43119 11132 43131 11135
rect 44192 11132 44220 11163
rect 44560 11132 44588 11172
rect 45830 11160 45836 11172
rect 45888 11160 45894 11212
rect 46308 11209 46336 11240
rect 47857 11237 47869 11271
rect 47903 11268 47915 11271
rect 48314 11268 48320 11280
rect 47903 11240 48320 11268
rect 47903 11237 47915 11240
rect 47857 11231 47915 11237
rect 48314 11228 48320 11240
rect 48372 11228 48378 11280
rect 46293 11203 46351 11209
rect 46293 11169 46305 11203
rect 46339 11169 46351 11203
rect 46293 11163 46351 11169
rect 46934 11160 46940 11212
rect 46992 11200 46998 11212
rect 47213 11203 47271 11209
rect 47213 11200 47225 11203
rect 46992 11172 47225 11200
rect 46992 11160 46998 11172
rect 47213 11169 47225 11172
rect 47259 11169 47271 11203
rect 47213 11163 47271 11169
rect 49973 11203 50031 11209
rect 49973 11169 49985 11203
rect 50019 11200 50031 11203
rect 50338 11200 50344 11212
rect 50019 11172 50344 11200
rect 50019 11169 50031 11172
rect 49973 11163 50031 11169
rect 50338 11160 50344 11172
rect 50396 11160 50402 11212
rect 50433 11203 50491 11209
rect 50433 11169 50445 11203
rect 50479 11200 50491 11203
rect 50724 11200 50752 11296
rect 50985 11271 51043 11277
rect 50985 11237 50997 11271
rect 51031 11268 51043 11271
rect 51166 11268 51172 11280
rect 51031 11240 51172 11268
rect 51031 11237 51043 11240
rect 50985 11231 51043 11237
rect 51166 11228 51172 11240
rect 51224 11228 51230 11280
rect 50479 11172 50752 11200
rect 50479 11169 50491 11172
rect 50433 11163 50491 11169
rect 51258 11160 51264 11212
rect 51316 11200 51322 11212
rect 51828 11209 51856 11308
rect 52917 11305 52929 11339
rect 52963 11336 52975 11339
rect 52963 11308 56272 11336
rect 52963 11305 52975 11308
rect 52917 11299 52975 11305
rect 51537 11203 51595 11209
rect 51537 11200 51549 11203
rect 51316 11172 51549 11200
rect 51316 11160 51322 11172
rect 51537 11169 51549 11172
rect 51583 11169 51595 11203
rect 51537 11163 51595 11169
rect 51813 11203 51871 11209
rect 51813 11169 51825 11203
rect 51859 11169 51871 11203
rect 51813 11163 51871 11169
rect 53024 11144 53052 11308
rect 54389 11271 54447 11277
rect 54389 11237 54401 11271
rect 54435 11268 54447 11271
rect 55398 11268 55404 11280
rect 54435 11240 55404 11268
rect 54435 11237 54447 11240
rect 54389 11231 54447 11237
rect 55398 11228 55404 11240
rect 55456 11228 55462 11280
rect 43119 11104 44128 11132
rect 44192 11104 44588 11132
rect 43119 11101 43131 11104
rect 43073 11095 43131 11101
rect 44100 11064 44128 11104
rect 44910 11092 44916 11144
rect 44968 11132 44974 11144
rect 45557 11135 45615 11141
rect 45557 11132 45569 11135
rect 44968 11104 45569 11132
rect 44968 11092 44974 11104
rect 45557 11101 45569 11104
rect 45603 11101 45615 11135
rect 45557 11095 45615 11101
rect 47397 11135 47455 11141
rect 47397 11101 47409 11135
rect 47443 11132 47455 11135
rect 47443 11104 48268 11132
rect 47443 11101 47455 11104
rect 47397 11095 47455 11101
rect 45005 11067 45063 11073
rect 45005 11064 45017 11067
rect 44100 11036 45017 11064
rect 45005 11033 45017 11036
rect 45051 11033 45063 11067
rect 45005 11027 45063 11033
rect 47486 11024 47492 11076
rect 47544 11024 47550 11076
rect 48240 11008 48268 11104
rect 48498 11092 48504 11144
rect 48556 11092 48562 11144
rect 51350 11092 51356 11144
rect 51408 11092 51414 11144
rect 53006 11092 53012 11144
rect 53064 11092 53070 11144
rect 54481 11135 54539 11141
rect 54481 11132 54493 11135
rect 53484 11104 54493 11132
rect 49510 11064 49516 11076
rect 48884 11036 49516 11064
rect 38470 10996 38476 11008
rect 37660 10968 38476 10996
rect 38470 10956 38476 10968
rect 38528 10956 38534 11008
rect 38746 10956 38752 11008
rect 38804 10996 38810 11008
rect 39853 10999 39911 11005
rect 39853 10996 39865 10999
rect 38804 10968 39865 10996
rect 38804 10956 38810 10968
rect 39853 10965 39865 10968
rect 39899 10965 39911 10999
rect 39853 10959 39911 10965
rect 42518 10956 42524 11008
rect 42576 10956 42582 11008
rect 42886 10956 42892 11008
rect 42944 10996 42950 11008
rect 42981 10999 43039 11005
rect 42981 10996 42993 10999
rect 42944 10968 42993 10996
rect 42944 10956 42950 10968
rect 42981 10965 42993 10968
rect 43027 10996 43039 10999
rect 44361 10999 44419 11005
rect 44361 10996 44373 10999
rect 43027 10968 44373 10996
rect 43027 10965 43039 10968
rect 42981 10959 43039 10965
rect 44361 10965 44373 10968
rect 44407 10965 44419 10999
rect 44361 10959 44419 10965
rect 45738 10956 45744 11008
rect 45796 10956 45802 11008
rect 46014 10956 46020 11008
rect 46072 10996 46078 11008
rect 46661 10999 46719 11005
rect 46661 10996 46673 10999
rect 46072 10968 46673 10996
rect 46072 10956 46078 10968
rect 46661 10965 46673 10968
rect 46707 10965 46719 10999
rect 46661 10959 46719 10965
rect 47946 10956 47952 11008
rect 48004 10956 48010 11008
rect 48222 10956 48228 11008
rect 48280 10956 48286 11008
rect 48774 10956 48780 11008
rect 48832 10996 48838 11008
rect 48884 11005 48912 11036
rect 49510 11024 49516 11036
rect 49568 11024 49574 11076
rect 50430 11024 50436 11076
rect 50488 11064 50494 11076
rect 50525 11067 50583 11073
rect 50525 11064 50537 11067
rect 50488 11036 50537 11064
rect 50488 11024 50494 11036
rect 50525 11033 50537 11036
rect 50571 11064 50583 11067
rect 51445 11067 51503 11073
rect 51445 11064 51457 11067
rect 50571 11036 51457 11064
rect 50571 11033 50583 11036
rect 50525 11027 50583 11033
rect 51445 11033 51457 11036
rect 51491 11033 51503 11067
rect 51445 11027 51503 11033
rect 53276 11067 53334 11073
rect 53276 11033 53288 11067
rect 53322 11033 53334 11067
rect 53276 11027 53334 11033
rect 48869 10999 48927 11005
rect 48869 10996 48881 10999
rect 48832 10968 48881 10996
rect 48832 10956 48838 10968
rect 48869 10965 48881 10968
rect 48915 10965 48927 10999
rect 48869 10959 48927 10965
rect 49142 10956 49148 11008
rect 49200 10996 49206 11008
rect 52270 10996 52276 11008
rect 49200 10968 52276 10996
rect 49200 10956 49206 10968
rect 52270 10956 52276 10968
rect 52328 10956 52334 11008
rect 52457 10999 52515 11005
rect 52457 10965 52469 10999
rect 52503 10996 52515 10999
rect 52638 10996 52644 11008
rect 52503 10968 52644 10996
rect 52503 10965 52515 10968
rect 52457 10959 52515 10965
rect 52638 10956 52644 10968
rect 52696 10956 52702 11008
rect 53300 10996 53328 11027
rect 53484 10996 53512 11104
rect 54481 11101 54493 11104
rect 54527 11101 54539 11135
rect 54481 11095 54539 11101
rect 55030 11092 55036 11144
rect 55088 11092 55094 11144
rect 56244 11141 56272 11308
rect 56594 11141 56600 11144
rect 56229 11135 56287 11141
rect 56229 11101 56241 11135
rect 56275 11132 56287 11135
rect 56321 11135 56379 11141
rect 56321 11132 56333 11135
rect 56275 11104 56333 11132
rect 56275 11101 56287 11104
rect 56229 11095 56287 11101
rect 56321 11101 56333 11104
rect 56367 11101 56379 11135
rect 56588 11132 56600 11141
rect 56555 11104 56600 11132
rect 56321 11095 56379 11101
rect 56588 11095 56600 11104
rect 56594 11092 56600 11095
rect 56652 11092 56658 11144
rect 58345 11135 58403 11141
rect 58345 11132 58357 11135
rect 57716 11104 58357 11132
rect 53300 10968 53512 10996
rect 56594 10956 56600 11008
rect 56652 10996 56658 11008
rect 57716 11005 57744 11104
rect 58345 11101 58357 11104
rect 58391 11101 58403 11135
rect 58345 11095 58403 11101
rect 57790 11024 57796 11076
rect 57848 11024 57854 11076
rect 57701 10999 57759 11005
rect 57701 10996 57713 10999
rect 56652 10968 57713 10996
rect 56652 10956 56658 10968
rect 57701 10965 57713 10968
rect 57747 10965 57759 10999
rect 57701 10959 57759 10965
rect 1104 10906 59040 10928
rect 1104 10854 15394 10906
rect 15446 10854 15458 10906
rect 15510 10854 15522 10906
rect 15574 10854 15586 10906
rect 15638 10854 15650 10906
rect 15702 10854 29838 10906
rect 29890 10854 29902 10906
rect 29954 10854 29966 10906
rect 30018 10854 30030 10906
rect 30082 10854 30094 10906
rect 30146 10854 44282 10906
rect 44334 10854 44346 10906
rect 44398 10854 44410 10906
rect 44462 10854 44474 10906
rect 44526 10854 44538 10906
rect 44590 10854 58726 10906
rect 58778 10854 58790 10906
rect 58842 10854 58854 10906
rect 58906 10854 58918 10906
rect 58970 10854 58982 10906
rect 59034 10854 59040 10906
rect 1104 10832 59040 10854
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 4856 10764 5641 10792
rect 4856 10752 4862 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 11333 10795 11391 10801
rect 5629 10755 5687 10761
rect 8680 10764 11284 10792
rect 4157 10727 4215 10733
rect 4157 10724 4169 10727
rect 3436 10696 4169 10724
rect 2866 10616 2872 10668
rect 2924 10616 2930 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3142 10656 3148 10668
rect 3099 10628 3148 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3436 10665 3464 10696
rect 4157 10693 4169 10696
rect 4203 10693 4215 10727
rect 4157 10687 4215 10693
rect 3421 10659 3479 10665
rect 3421 10656 3433 10659
rect 3200 10628 3433 10656
rect 3200 10616 3206 10628
rect 3421 10625 3433 10628
rect 3467 10625 3479 10659
rect 3878 10656 3884 10668
rect 3421 10619 3479 10625
rect 3528 10628 3884 10656
rect 3528 10597 3556 10628
rect 3878 10616 3884 10628
rect 3936 10656 3942 10668
rect 4062 10656 4068 10668
rect 3936 10628 4068 10656
rect 3936 10616 3942 10628
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4338 10616 4344 10668
rect 4396 10616 4402 10668
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10557 3571 10591
rect 5644 10588 5672 10616
rect 6086 10588 6092 10600
rect 5644 10560 6092 10588
rect 3513 10551 3571 10557
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8570 10588 8576 10600
rect 8527 10560 8576 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8570 10548 8576 10560
rect 8628 10588 8634 10600
rect 8680 10588 8708 10764
rect 11256 10736 11284 10764
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11422 10792 11428 10804
rect 11379 10764 11428 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 11790 10792 11796 10804
rect 11572 10764 11796 10792
rect 11572 10752 11578 10764
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 14550 10752 14556 10804
rect 14608 10752 14614 10804
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15286 10792 15292 10804
rect 15059 10764 15292 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 17126 10792 17132 10804
rect 16546 10764 17132 10792
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 9861 10727 9919 10733
rect 9861 10724 9873 10727
rect 9732 10696 9873 10724
rect 9732 10684 9738 10696
rect 9861 10693 9873 10696
rect 9907 10693 9919 10727
rect 9861 10687 9919 10693
rect 11238 10684 11244 10736
rect 11296 10684 11302 10736
rect 13906 10724 13912 10736
rect 13096 10696 13912 10724
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9490 10656 9496 10668
rect 8904 10628 9496 10656
rect 8904 10616 8910 10628
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10209 10659 10267 10665
rect 10209 10656 10221 10659
rect 10100 10628 10221 10656
rect 10100 10616 10106 10628
rect 10209 10625 10221 10628
rect 10255 10625 10267 10659
rect 10209 10619 10267 10625
rect 8628 10560 8708 10588
rect 8628 10548 8634 10560
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8812 10560 9045 10588
rect 8812 10548 8818 10560
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3326 10520 3332 10532
rect 2915 10492 3332 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 3789 10523 3847 10529
rect 3789 10489 3801 10523
rect 3835 10520 3847 10523
rect 4246 10520 4252 10532
rect 3835 10492 4252 10520
rect 3835 10489 3847 10492
rect 3789 10483 3847 10489
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 4341 10523 4399 10529
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 4430 10520 4436 10532
rect 4387 10492 4436 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 8956 10464 8984 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9950 10548 9956 10600
rect 10008 10548 10014 10600
rect 13096 10597 13124 10696
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 16546 10724 16574 10764
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 17644 10764 18061 10792
rect 17644 10752 17650 10764
rect 18049 10761 18061 10764
rect 18095 10792 18107 10795
rect 18966 10792 18972 10804
rect 18095 10764 18972 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10792 20499 10795
rect 20806 10792 20812 10804
rect 20487 10764 20812 10792
rect 20487 10761 20499 10764
rect 20441 10755 20499 10761
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 20901 10795 20959 10801
rect 20901 10761 20913 10795
rect 20947 10792 20959 10795
rect 22094 10792 22100 10804
rect 20947 10764 22100 10792
rect 20947 10761 20959 10764
rect 20901 10755 20959 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 22428 10764 22845 10792
rect 22428 10752 22434 10764
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 25409 10795 25467 10801
rect 22833 10755 22891 10761
rect 23216 10764 25268 10792
rect 14792 10696 16574 10724
rect 16936 10727 16994 10733
rect 14792 10684 14798 10696
rect 16936 10693 16948 10727
rect 16982 10724 16994 10727
rect 17034 10724 17040 10736
rect 16982 10696 17040 10724
rect 16982 10693 16994 10696
rect 16936 10687 16994 10693
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 17144 10724 17172 10752
rect 21545 10727 21603 10733
rect 21545 10724 21557 10727
rect 17144 10696 20392 10724
rect 13354 10665 13360 10668
rect 13348 10619 13360 10665
rect 13354 10616 13360 10619
rect 13412 10616 13418 10668
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 16758 10656 16764 10668
rect 14976 10628 16764 10656
rect 14976 10616 14982 10628
rect 16758 10616 16764 10628
rect 16816 10656 16822 10668
rect 17770 10656 17776 10668
rect 16816 10628 17776 10656
rect 16816 10616 16822 10628
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 19978 10616 19984 10668
rect 20036 10616 20042 10668
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12406 10560 13093 10588
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 6822 10452 6828 10464
rect 6687 10424 6828 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6822 10412 6828 10424
rect 6880 10452 6886 10464
rect 8018 10452 8024 10464
rect 6880 10424 8024 10452
rect 6880 10412 6886 10424
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8938 10412 8944 10464
rect 8996 10412 9002 10464
rect 9968 10452 9996 10548
rect 10870 10452 10876 10464
rect 9968 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10452 10934 10464
rect 12406 10452 12434 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14148 10560 15117 10588
rect 14148 10548 14154 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 12986 10480 12992 10532
rect 13044 10480 13050 10532
rect 14461 10523 14519 10529
rect 14461 10489 14473 10523
rect 14507 10520 14519 10523
rect 15838 10520 15844 10532
rect 14507 10492 15844 10520
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 15838 10480 15844 10492
rect 15896 10520 15902 10532
rect 15948 10520 15976 10551
rect 16666 10548 16672 10600
rect 16724 10548 16730 10600
rect 20364 10597 20392 10696
rect 20456 10696 21557 10724
rect 20456 10668 20484 10696
rect 21545 10693 21557 10696
rect 21591 10724 21603 10727
rect 23216 10724 23244 10764
rect 25240 10736 25268 10764
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 25498 10792 25504 10804
rect 25455 10764 25504 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 25777 10795 25835 10801
rect 25777 10761 25789 10795
rect 25823 10792 25835 10795
rect 26694 10792 26700 10804
rect 25823 10764 26700 10792
rect 25823 10761 25835 10764
rect 25777 10755 25835 10761
rect 26694 10752 26700 10764
rect 26752 10752 26758 10804
rect 29730 10752 29736 10804
rect 29788 10792 29794 10804
rect 30009 10795 30067 10801
rect 30009 10792 30021 10795
rect 29788 10764 30021 10792
rect 29788 10752 29794 10764
rect 30009 10761 30021 10764
rect 30055 10761 30067 10795
rect 30009 10755 30067 10761
rect 30650 10752 30656 10804
rect 30708 10792 30714 10804
rect 40497 10795 40555 10801
rect 30708 10764 39068 10792
rect 30708 10752 30714 10764
rect 21591 10696 23244 10724
rect 21591 10693 21603 10696
rect 21545 10687 21603 10693
rect 25222 10684 25228 10736
rect 25280 10724 25286 10736
rect 27430 10724 27436 10736
rect 25280 10696 27436 10724
rect 25280 10684 25286 10696
rect 27430 10684 27436 10696
rect 27488 10684 27494 10736
rect 27890 10684 27896 10736
rect 27948 10724 27954 10736
rect 28138 10727 28196 10733
rect 28138 10724 28150 10727
rect 27948 10696 28150 10724
rect 27948 10684 27954 10696
rect 28138 10693 28150 10696
rect 28184 10693 28196 10727
rect 28138 10687 28196 10693
rect 33260 10727 33318 10733
rect 33260 10693 33272 10727
rect 33306 10724 33318 10727
rect 33306 10696 33640 10724
rect 33306 10693 33318 10696
rect 33260 10687 33318 10693
rect 20438 10616 20444 10668
rect 20496 10616 20502 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 20855 10628 21833 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 23658 10616 23664 10668
rect 23716 10616 23722 10668
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 24673 10659 24731 10665
rect 24673 10625 24685 10659
rect 24719 10656 24731 10659
rect 24762 10656 24768 10668
rect 24719 10628 24768 10656
rect 24719 10625 24731 10628
rect 24673 10619 24731 10625
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 24857 10659 24915 10665
rect 24857 10625 24869 10659
rect 24903 10656 24915 10659
rect 24946 10656 24952 10668
rect 24903 10628 24952 10656
rect 24903 10625 24915 10628
rect 24857 10619 24915 10625
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 26510 10656 26516 10668
rect 25424 10628 26516 10656
rect 25424 10600 25452 10628
rect 20349 10591 20407 10597
rect 20349 10557 20361 10591
rect 20395 10588 20407 10591
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 20395 10560 21097 10588
rect 20395 10557 20407 10560
rect 20349 10551 20407 10557
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 15896 10492 15976 10520
rect 21100 10520 21128 10551
rect 22462 10548 22468 10600
rect 22520 10588 22526 10600
rect 23799 10591 23857 10597
rect 23799 10588 23811 10591
rect 22520 10560 23811 10588
rect 22520 10548 22526 10560
rect 23799 10557 23811 10560
rect 23845 10557 23857 10591
rect 23799 10551 23857 10557
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24213 10591 24271 10597
rect 24213 10588 24225 10591
rect 24176 10560 24225 10588
rect 24176 10548 24182 10560
rect 24213 10557 24225 10560
rect 24259 10588 24271 10591
rect 24486 10588 24492 10600
rect 24259 10560 24492 10588
rect 24259 10557 24271 10560
rect 24213 10551 24271 10557
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 25406 10548 25412 10600
rect 25464 10548 25470 10600
rect 25682 10548 25688 10600
rect 25740 10588 25746 10600
rect 25976 10597 26004 10628
rect 26510 10616 26516 10628
rect 26568 10616 26574 10668
rect 29362 10616 29368 10668
rect 29420 10616 29426 10668
rect 30926 10665 30932 10668
rect 30904 10659 30932 10665
rect 30904 10625 30916 10659
rect 30904 10619 30932 10625
rect 30926 10616 30932 10619
rect 30984 10616 30990 10668
rect 31018 10616 31024 10668
rect 31076 10616 31082 10668
rect 32766 10656 32772 10668
rect 31588 10628 32772 10656
rect 25869 10591 25927 10597
rect 25869 10588 25881 10591
rect 25740 10560 25881 10588
rect 25740 10548 25746 10560
rect 25869 10557 25881 10560
rect 25915 10557 25927 10591
rect 25869 10551 25927 10557
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 27614 10548 27620 10600
rect 27672 10588 27678 10600
rect 27893 10591 27951 10597
rect 27893 10588 27905 10591
rect 27672 10560 27905 10588
rect 27672 10548 27678 10560
rect 27893 10557 27905 10560
rect 27939 10557 27951 10591
rect 27893 10551 27951 10557
rect 30558 10548 30564 10600
rect 30616 10588 30622 10600
rect 30745 10591 30803 10597
rect 30745 10588 30757 10591
rect 30616 10560 30757 10588
rect 30616 10548 30622 10560
rect 30745 10557 30757 10560
rect 30791 10557 30803 10591
rect 30745 10551 30803 10557
rect 31294 10548 31300 10600
rect 31352 10588 31358 10600
rect 31588 10588 31616 10628
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 33410 10616 33416 10668
rect 33468 10656 33474 10668
rect 33505 10659 33563 10665
rect 33505 10656 33517 10659
rect 33468 10628 33517 10656
rect 33468 10616 33474 10628
rect 33505 10625 33517 10628
rect 33551 10625 33563 10659
rect 33612 10656 33640 10696
rect 33778 10684 33784 10736
rect 33836 10724 33842 10736
rect 34057 10727 34115 10733
rect 34057 10724 34069 10727
rect 33836 10696 34069 10724
rect 33836 10684 33842 10696
rect 34057 10693 34069 10696
rect 34103 10693 34115 10727
rect 34057 10687 34115 10693
rect 35428 10727 35486 10733
rect 35428 10693 35440 10727
rect 35474 10724 35486 10727
rect 35710 10724 35716 10736
rect 35474 10696 35716 10724
rect 35474 10693 35486 10696
rect 35428 10687 35486 10693
rect 35710 10684 35716 10696
rect 35768 10684 35774 10736
rect 36906 10684 36912 10736
rect 36964 10684 36970 10736
rect 39040 10733 39068 10764
rect 40497 10761 40509 10795
rect 40543 10792 40555 10795
rect 40770 10792 40776 10804
rect 40543 10764 40776 10792
rect 40543 10761 40555 10764
rect 40497 10755 40555 10761
rect 40770 10752 40776 10764
rect 40828 10752 40834 10804
rect 41230 10752 41236 10804
rect 41288 10792 41294 10804
rect 41325 10795 41383 10801
rect 41325 10792 41337 10795
rect 41288 10764 41337 10792
rect 41288 10752 41294 10764
rect 41325 10761 41337 10764
rect 41371 10792 41383 10795
rect 42153 10795 42211 10801
rect 42153 10792 42165 10795
rect 41371 10764 42165 10792
rect 41371 10761 41383 10764
rect 41325 10755 41383 10761
rect 42153 10761 42165 10764
rect 42199 10761 42211 10795
rect 42153 10755 42211 10761
rect 45281 10795 45339 10801
rect 45281 10761 45293 10795
rect 45327 10792 45339 10795
rect 45646 10792 45652 10804
rect 45327 10764 45652 10792
rect 45327 10761 45339 10764
rect 45281 10755 45339 10761
rect 39025 10727 39083 10733
rect 39025 10693 39037 10727
rect 39071 10693 39083 10727
rect 39025 10687 39083 10693
rect 33870 10656 33876 10668
rect 33612 10628 33876 10656
rect 33505 10619 33563 10625
rect 33870 10616 33876 10628
rect 33928 10616 33934 10668
rect 33965 10659 34023 10665
rect 33965 10625 33977 10659
rect 34011 10625 34023 10659
rect 33965 10619 34023 10625
rect 31352 10560 31616 10588
rect 31757 10591 31815 10597
rect 31352 10548 31358 10560
rect 31757 10557 31769 10591
rect 31803 10557 31815 10591
rect 31757 10551 31815 10557
rect 31941 10591 31999 10597
rect 31941 10557 31953 10591
rect 31987 10588 31999 10591
rect 31987 10560 32168 10588
rect 31987 10557 31999 10560
rect 31941 10551 31999 10557
rect 31772 10520 31800 10551
rect 21100 10492 23244 10520
rect 15896 10480 15902 10492
rect 10928 10424 12434 10452
rect 10928 10412 10934 10424
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 18322 10452 18328 10464
rect 16080 10424 18328 10452
rect 16080 10412 16086 10424
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19242 10452 19248 10464
rect 18748 10424 19248 10452
rect 18748 10412 18754 10424
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 23014 10412 23020 10464
rect 23072 10412 23078 10464
rect 23216 10452 23244 10492
rect 25240 10492 27936 10520
rect 31772 10492 31984 10520
rect 23750 10452 23756 10464
rect 23216 10424 23756 10452
rect 23750 10412 23756 10424
rect 23808 10452 23814 10464
rect 25240 10452 25268 10492
rect 23808 10424 25268 10452
rect 25317 10455 25375 10461
rect 23808 10412 23814 10424
rect 25317 10421 25329 10455
rect 25363 10452 25375 10455
rect 25406 10452 25412 10464
rect 25363 10424 25412 10452
rect 25363 10421 25375 10424
rect 25317 10415 25375 10421
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 27908 10452 27936 10492
rect 31956 10464 31984 10492
rect 28994 10452 29000 10464
rect 27908 10424 29000 10452
rect 28994 10412 29000 10424
rect 29052 10412 29058 10464
rect 29270 10412 29276 10464
rect 29328 10412 29334 10464
rect 30101 10455 30159 10461
rect 30101 10421 30113 10455
rect 30147 10452 30159 10455
rect 31202 10452 31208 10464
rect 30147 10424 31208 10452
rect 30147 10421 30159 10424
rect 30101 10415 30159 10421
rect 31202 10412 31208 10424
rect 31260 10412 31266 10464
rect 31938 10412 31944 10464
rect 31996 10412 32002 10464
rect 32140 10461 32168 10560
rect 33686 10548 33692 10600
rect 33744 10588 33750 10600
rect 33980 10588 34008 10619
rect 34514 10616 34520 10668
rect 34572 10656 34578 10668
rect 35161 10659 35219 10665
rect 35161 10656 35173 10659
rect 34572 10628 35173 10656
rect 34572 10616 34578 10628
rect 35161 10625 35173 10628
rect 35207 10625 35219 10659
rect 35161 10619 35219 10625
rect 37366 10616 37372 10668
rect 37424 10656 37430 10668
rect 37553 10659 37611 10665
rect 37553 10656 37565 10659
rect 37424 10628 37565 10656
rect 37424 10616 37430 10628
rect 37553 10625 37565 10628
rect 37599 10625 37611 10659
rect 37553 10619 37611 10625
rect 37642 10616 37648 10668
rect 37700 10656 37706 10668
rect 37809 10659 37867 10665
rect 37809 10656 37821 10659
rect 37700 10628 37821 10656
rect 37700 10616 37706 10628
rect 37809 10625 37821 10628
rect 37855 10625 37867 10659
rect 42168 10656 42196 10755
rect 45646 10752 45652 10764
rect 45704 10752 45710 10804
rect 47762 10752 47768 10804
rect 47820 10792 47826 10804
rect 47857 10795 47915 10801
rect 47857 10792 47869 10795
rect 47820 10764 47869 10792
rect 47820 10752 47826 10764
rect 47857 10761 47869 10764
rect 47903 10761 47915 10795
rect 47857 10755 47915 10761
rect 47946 10752 47952 10804
rect 48004 10752 48010 10804
rect 48317 10795 48375 10801
rect 48317 10761 48329 10795
rect 48363 10792 48375 10795
rect 48498 10792 48504 10804
rect 48363 10764 48504 10792
rect 48363 10761 48375 10764
rect 48317 10755 48375 10761
rect 48498 10752 48504 10764
rect 48556 10752 48562 10804
rect 50798 10792 50804 10804
rect 48608 10764 50660 10792
rect 43714 10724 43720 10736
rect 42444 10696 43720 10724
rect 42444 10668 42472 10696
rect 43714 10684 43720 10696
rect 43772 10724 43778 10736
rect 44168 10727 44226 10733
rect 43772 10696 43944 10724
rect 43772 10684 43778 10696
rect 42426 10656 42432 10668
rect 42168 10628 42432 10656
rect 37809 10619 37867 10625
rect 42426 10616 42432 10628
rect 42484 10616 42490 10668
rect 42518 10616 42524 10668
rect 42576 10656 42582 10668
rect 43916 10665 43944 10696
rect 44168 10693 44180 10727
rect 44214 10724 44226 10727
rect 45738 10724 45744 10736
rect 44214 10696 45744 10724
rect 44214 10693 44226 10696
rect 44168 10687 44226 10693
rect 45738 10684 45744 10696
rect 45796 10684 45802 10736
rect 46284 10727 46342 10733
rect 46284 10693 46296 10727
rect 46330 10724 46342 10727
rect 47964 10724 47992 10752
rect 46330 10696 47992 10724
rect 46330 10693 46342 10696
rect 46284 10687 46342 10693
rect 42685 10659 42743 10665
rect 42685 10656 42697 10659
rect 42576 10628 42697 10656
rect 42576 10616 42582 10628
rect 42685 10625 42697 10628
rect 42731 10625 42743 10659
rect 42685 10619 42743 10625
rect 43901 10659 43959 10665
rect 43901 10625 43913 10659
rect 43947 10625 43959 10659
rect 43901 10619 43959 10625
rect 44450 10616 44456 10668
rect 44508 10656 44514 10668
rect 47949 10659 48007 10665
rect 44508 10628 47808 10656
rect 44508 10616 44514 10628
rect 33744 10560 34008 10588
rect 34241 10591 34299 10597
rect 33744 10548 33750 10560
rect 34241 10557 34253 10591
rect 34287 10588 34299 10591
rect 34606 10588 34612 10600
rect 34287 10560 34612 10588
rect 34287 10557 34299 10560
rect 34241 10551 34299 10557
rect 34606 10548 34612 10560
rect 34664 10588 34670 10600
rect 34664 10560 34744 10588
rect 34664 10548 34670 10560
rect 33597 10523 33655 10529
rect 33597 10489 33609 10523
rect 33643 10520 33655 10523
rect 34422 10520 34428 10532
rect 33643 10492 34428 10520
rect 33643 10489 33655 10492
rect 33597 10483 33655 10489
rect 34422 10480 34428 10492
rect 34480 10480 34486 10532
rect 32125 10455 32183 10461
rect 32125 10421 32137 10455
rect 32171 10452 32183 10455
rect 33134 10452 33140 10464
rect 32171 10424 33140 10452
rect 32171 10421 32183 10424
rect 32125 10415 32183 10421
rect 33134 10412 33140 10424
rect 33192 10412 33198 10464
rect 34716 10461 34744 10560
rect 39206 10548 39212 10600
rect 39264 10548 39270 10600
rect 44910 10548 44916 10600
rect 44968 10548 44974 10600
rect 45649 10591 45707 10597
rect 45649 10557 45661 10591
rect 45695 10588 45707 10591
rect 45830 10588 45836 10600
rect 45695 10560 45836 10588
rect 45695 10557 45707 10560
rect 45649 10551 45707 10557
rect 45830 10548 45836 10560
rect 45888 10548 45894 10600
rect 46014 10548 46020 10600
rect 46072 10548 46078 10600
rect 47302 10548 47308 10600
rect 47360 10588 47366 10600
rect 47673 10591 47731 10597
rect 47673 10588 47685 10591
rect 47360 10560 47685 10588
rect 47360 10548 47366 10560
rect 47673 10557 47685 10560
rect 47719 10557 47731 10591
rect 47780 10588 47808 10628
rect 47949 10625 47961 10659
rect 47995 10656 48007 10659
rect 48222 10656 48228 10668
rect 47995 10628 48228 10656
rect 47995 10625 48007 10628
rect 47949 10619 48007 10625
rect 48222 10616 48228 10628
rect 48280 10616 48286 10668
rect 48608 10588 48636 10764
rect 49510 10616 49516 10668
rect 49568 10616 49574 10668
rect 49786 10616 49792 10668
rect 49844 10616 49850 10668
rect 47780 10560 48636 10588
rect 47673 10551 47731 10557
rect 49142 10548 49148 10600
rect 49200 10548 49206 10600
rect 49602 10548 49608 10600
rect 49660 10597 49666 10600
rect 49660 10591 49709 10597
rect 49660 10557 49663 10591
rect 49697 10557 49709 10591
rect 49660 10551 49709 10557
rect 49660 10548 49666 10551
rect 49970 10548 49976 10600
rect 50028 10588 50034 10600
rect 50065 10591 50123 10597
rect 50065 10588 50077 10591
rect 50028 10560 50077 10588
rect 50028 10548 50034 10560
rect 50065 10557 50077 10560
rect 50111 10557 50123 10591
rect 50065 10551 50123 10557
rect 50525 10591 50583 10597
rect 50525 10557 50537 10591
rect 50571 10557 50583 10591
rect 50632 10588 50660 10764
rect 50724 10764 50804 10792
rect 50724 10665 50752 10764
rect 50798 10752 50804 10764
rect 50856 10752 50862 10804
rect 56410 10792 56416 10804
rect 51046 10764 56416 10792
rect 50709 10659 50767 10665
rect 50709 10625 50721 10659
rect 50755 10625 50767 10659
rect 50709 10619 50767 10625
rect 51046 10588 51074 10764
rect 56410 10752 56416 10764
rect 56468 10752 56474 10804
rect 51936 10727 51994 10733
rect 51936 10693 51948 10727
rect 51982 10724 51994 10727
rect 52638 10724 52644 10736
rect 51982 10696 52644 10724
rect 51982 10693 51994 10696
rect 51936 10687 51994 10693
rect 52638 10684 52644 10696
rect 52696 10684 52702 10736
rect 52181 10659 52239 10665
rect 52181 10625 52193 10659
rect 52227 10656 52239 10659
rect 52454 10656 52460 10668
rect 52227 10628 52460 10656
rect 52227 10625 52239 10628
rect 52181 10619 52239 10625
rect 52454 10616 52460 10628
rect 52512 10656 52518 10668
rect 52549 10659 52607 10665
rect 52549 10656 52561 10659
rect 52512 10628 52561 10656
rect 52512 10616 52518 10628
rect 52549 10625 52561 10628
rect 52595 10656 52607 10659
rect 52917 10659 52975 10665
rect 52917 10656 52929 10659
rect 52595 10628 52929 10656
rect 52595 10625 52607 10628
rect 52549 10619 52607 10625
rect 52917 10625 52929 10628
rect 52963 10656 52975 10659
rect 53006 10656 53012 10668
rect 52963 10628 53012 10656
rect 52963 10625 52975 10628
rect 52917 10619 52975 10625
rect 53006 10616 53012 10628
rect 53064 10616 53070 10668
rect 53190 10665 53196 10668
rect 53184 10619 53196 10665
rect 53190 10616 53196 10619
rect 53248 10616 53254 10668
rect 55122 10616 55128 10668
rect 55180 10616 55186 10668
rect 55398 10616 55404 10668
rect 55456 10616 55462 10668
rect 56137 10659 56195 10665
rect 56137 10625 56149 10659
rect 56183 10656 56195 10659
rect 56594 10656 56600 10668
rect 56183 10628 56600 10656
rect 56183 10625 56195 10628
rect 56137 10619 56195 10625
rect 56594 10616 56600 10628
rect 56652 10616 56658 10668
rect 56781 10659 56839 10665
rect 56781 10625 56793 10659
rect 56827 10656 56839 10659
rect 56962 10656 56968 10668
rect 56827 10628 56968 10656
rect 56827 10625 56839 10628
rect 56781 10619 56839 10625
rect 56962 10616 56968 10628
rect 57020 10616 57026 10668
rect 54570 10588 54576 10600
rect 50632 10560 51074 10588
rect 54312 10560 54576 10588
rect 50525 10551 50583 10557
rect 36541 10523 36599 10529
rect 36541 10489 36553 10523
rect 36587 10520 36599 10523
rect 37550 10520 37556 10532
rect 36587 10492 37556 10520
rect 36587 10489 36599 10492
rect 36541 10483 36599 10489
rect 37550 10480 37556 10492
rect 37608 10480 37614 10532
rect 38933 10523 38991 10529
rect 38933 10489 38945 10523
rect 38979 10520 38991 10523
rect 39224 10520 39252 10548
rect 38979 10492 39252 10520
rect 38979 10489 38991 10492
rect 38933 10483 38991 10489
rect 34701 10455 34759 10461
rect 34701 10421 34713 10455
rect 34747 10452 34759 10455
rect 37734 10452 37740 10464
rect 34747 10424 37740 10452
rect 34747 10421 34759 10424
rect 34701 10415 34759 10421
rect 37734 10412 37740 10424
rect 37792 10412 37798 10464
rect 43809 10455 43867 10461
rect 43809 10421 43821 10455
rect 43855 10452 43867 10455
rect 43898 10452 43904 10464
rect 43855 10424 43904 10452
rect 43855 10421 43867 10424
rect 43809 10415 43867 10421
rect 43898 10412 43904 10424
rect 43956 10452 43962 10464
rect 44928 10452 44956 10548
rect 46032 10520 46060 10548
rect 45848 10492 46060 10520
rect 45848 10464 45876 10492
rect 43956 10424 44956 10452
rect 43956 10412 43962 10424
rect 45830 10412 45836 10464
rect 45888 10412 45894 10464
rect 47320 10452 47348 10548
rect 47397 10523 47455 10529
rect 47397 10489 47409 10523
rect 47443 10520 47455 10523
rect 48406 10520 48412 10532
rect 47443 10492 48412 10520
rect 47443 10489 47455 10492
rect 47397 10483 47455 10489
rect 48406 10480 48412 10492
rect 48464 10480 48470 10532
rect 49160 10520 49188 10548
rect 48608 10492 49188 10520
rect 48130 10452 48136 10464
rect 47320 10424 48136 10452
rect 48130 10412 48136 10424
rect 48188 10452 48194 10464
rect 48608 10461 48636 10492
rect 50540 10464 50568 10551
rect 54312 10529 54340 10560
rect 54570 10548 54576 10560
rect 54628 10588 54634 10600
rect 55263 10591 55321 10597
rect 55263 10588 55275 10591
rect 54628 10560 55275 10588
rect 54628 10548 54634 10560
rect 55263 10557 55275 10560
rect 55309 10557 55321 10591
rect 55263 10551 55321 10557
rect 56321 10591 56379 10597
rect 56321 10557 56333 10591
rect 56367 10557 56379 10591
rect 56321 10551 56379 10557
rect 56505 10591 56563 10597
rect 56505 10557 56517 10591
rect 56551 10588 56563 10591
rect 56551 10560 56640 10588
rect 56551 10557 56563 10560
rect 56505 10551 56563 10557
rect 54297 10523 54355 10529
rect 54297 10489 54309 10523
rect 54343 10489 54355 10523
rect 54297 10483 54355 10489
rect 55677 10523 55735 10529
rect 55677 10489 55689 10523
rect 55723 10489 55735 10523
rect 55677 10483 55735 10489
rect 48593 10455 48651 10461
rect 48593 10452 48605 10455
rect 48188 10424 48605 10452
rect 48188 10412 48194 10424
rect 48593 10421 48605 10424
rect 48639 10421 48651 10455
rect 48593 10415 48651 10421
rect 48869 10455 48927 10461
rect 48869 10421 48881 10455
rect 48915 10452 48927 10455
rect 50154 10452 50160 10464
rect 48915 10424 50160 10452
rect 48915 10421 48927 10424
rect 48869 10415 48927 10421
rect 50154 10412 50160 10424
rect 50212 10412 50218 10464
rect 50522 10412 50528 10464
rect 50580 10412 50586 10464
rect 54478 10412 54484 10464
rect 54536 10412 54542 10464
rect 55214 10412 55220 10464
rect 55272 10452 55278 10464
rect 55692 10452 55720 10483
rect 56336 10464 56364 10551
rect 56612 10464 56640 10560
rect 56686 10548 56692 10600
rect 56744 10548 56750 10600
rect 58437 10591 58495 10597
rect 58437 10557 58449 10591
rect 58483 10557 58495 10591
rect 58437 10551 58495 10557
rect 57149 10523 57207 10529
rect 57149 10489 57161 10523
rect 57195 10520 57207 10523
rect 58452 10520 58480 10551
rect 57195 10492 58480 10520
rect 57195 10489 57207 10492
rect 57149 10483 57207 10489
rect 55272 10424 55720 10452
rect 55272 10412 55278 10424
rect 56318 10412 56324 10464
rect 56376 10412 56382 10464
rect 56594 10412 56600 10464
rect 56652 10452 56658 10464
rect 56778 10452 56784 10464
rect 56652 10424 56784 10452
rect 56652 10412 56658 10424
rect 56778 10412 56784 10424
rect 56836 10452 56842 10464
rect 57425 10455 57483 10461
rect 57425 10452 57437 10455
rect 56836 10424 57437 10452
rect 56836 10412 56842 10424
rect 57425 10421 57437 10424
rect 57471 10421 57483 10455
rect 57425 10415 57483 10421
rect 57882 10412 57888 10464
rect 57940 10412 57946 10464
rect 1104 10362 58880 10384
rect 1104 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 22616 10362
rect 22668 10310 22680 10362
rect 22732 10310 22744 10362
rect 22796 10310 22808 10362
rect 22860 10310 22872 10362
rect 22924 10310 37060 10362
rect 37112 10310 37124 10362
rect 37176 10310 37188 10362
rect 37240 10310 37252 10362
rect 37304 10310 37316 10362
rect 37368 10310 51504 10362
rect 51556 10310 51568 10362
rect 51620 10310 51632 10362
rect 51684 10310 51696 10362
rect 51748 10310 51760 10362
rect 51812 10310 58880 10362
rect 1104 10288 58880 10310
rect 2866 10208 2872 10260
rect 2924 10208 2930 10260
rect 3142 10208 3148 10260
rect 3200 10208 3206 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 5868 10220 6745 10248
rect 5868 10208 5874 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 7742 10208 7748 10260
rect 7800 10208 7806 10260
rect 9122 10248 9128 10260
rect 7944 10220 9128 10248
rect 2884 10121 2912 10208
rect 6086 10140 6092 10192
rect 6144 10140 6150 10192
rect 7944 10189 7972 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9309 10251 9367 10257
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9398 10248 9404 10260
rect 9355 10220 9404 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10042 10248 10048 10260
rect 9723 10220 10048 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13354 10248 13360 10260
rect 13311 10220 13360 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 14918 10208 14924 10260
rect 14976 10208 14982 10260
rect 15378 10208 15384 10260
rect 15436 10208 15442 10260
rect 15838 10208 15844 10260
rect 15896 10208 15902 10260
rect 16298 10208 16304 10260
rect 16356 10248 16362 10260
rect 16356 10220 17724 10248
rect 16356 10208 16362 10220
rect 7929 10183 7987 10189
rect 7929 10149 7941 10183
rect 7975 10149 7987 10183
rect 7929 10143 7987 10149
rect 9030 10140 9036 10192
rect 9088 10180 9094 10192
rect 9585 10183 9643 10189
rect 9585 10180 9597 10183
rect 9088 10152 9597 10180
rect 9088 10140 9094 10152
rect 9585 10149 9597 10152
rect 9631 10149 9643 10183
rect 9585 10143 9643 10149
rect 14093 10183 14151 10189
rect 14093 10149 14105 10183
rect 14139 10149 14151 10183
rect 14936 10180 14964 10208
rect 14093 10143 14151 10149
rect 14568 10152 14964 10180
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10081 2927 10115
rect 4065 10115 4123 10121
rect 2869 10075 2927 10081
rect 3068 10084 3372 10112
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2655 10047 2713 10053
rect 2655 10013 2667 10047
rect 2701 10044 2713 10047
rect 2774 10044 2780 10056
rect 2701 10016 2780 10044
rect 2701 10013 2713 10016
rect 2655 10007 2713 10013
rect 2516 9976 2544 10007
rect 2774 10004 2780 10016
rect 2832 10044 2838 10056
rect 3068 10044 3096 10084
rect 3344 10053 3372 10084
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 6546 10112 6552 10124
rect 4111 10084 6552 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 3236 10047 3294 10053
rect 3236 10044 3248 10047
rect 2832 10016 3096 10044
rect 3215 10016 3248 10044
rect 2832 10004 2838 10016
rect 3236 10013 3248 10016
rect 3282 10013 3294 10047
rect 3236 10007 3294 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3050 9976 3056 9988
rect 2516 9948 3056 9976
rect 3050 9936 3056 9948
rect 3108 9976 3114 9988
rect 3252 9976 3280 10007
rect 4080 9976 4108 10075
rect 6546 10072 6552 10084
rect 6604 10112 6610 10124
rect 6604 10084 7604 10112
rect 6604 10072 6610 10084
rect 6333 10047 6391 10053
rect 6333 10013 6345 10047
rect 6379 10044 6391 10047
rect 6457 10047 6515 10053
rect 6379 10013 6408 10044
rect 6333 10007 6408 10013
rect 6457 10013 6469 10047
rect 6503 10044 6515 10047
rect 6822 10044 6828 10056
rect 6503 10016 6828 10044
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 6380 9976 6408 10007
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 6932 9976 6960 10007
rect 7576 9985 7604 10084
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 13909 10115 13967 10121
rect 9456 10084 9720 10112
rect 9456 10072 9462 10084
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8570 10044 8576 10056
rect 8159 10016 8576 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 3108 9948 4108 9976
rect 6288 9948 6960 9976
rect 7561 9979 7619 9985
rect 3108 9936 3114 9948
rect 6288 9920 6316 9948
rect 7561 9945 7573 9979
rect 7607 9976 7619 9979
rect 7650 9976 7656 9988
rect 7607 9948 7656 9976
rect 7607 9945 7619 9948
rect 7561 9939 7619 9945
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 7777 9979 7835 9985
rect 7777 9945 7789 9979
rect 7823 9976 7835 9979
rect 7944 9976 7972 10004
rect 7823 9948 7972 9976
rect 7823 9945 7835 9948
rect 7777 9939 7835 9945
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 8128 9908 8156 10007
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8938 10044 8944 10056
rect 8772 10016 8944 10044
rect 8662 9936 8668 9988
rect 8720 9936 8726 9988
rect 7515 9880 8156 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8772 9908 8800 10016
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9122 10053 9128 10056
rect 9111 10047 9128 10053
rect 9111 10013 9123 10047
rect 9111 10007 9128 10013
rect 9122 10004 9128 10007
rect 9180 10004 9186 10056
rect 9692 10053 9720 10084
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 14108 10112 14136 10143
rect 14568 10121 14596 10152
rect 13955 10084 14136 10112
rect 14553 10115 14611 10121
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14553 10081 14565 10115
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 14734 10072 14740 10124
rect 14792 10072 14798 10124
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 15396 10044 15424 10208
rect 15856 10112 15884 10208
rect 16347 10115 16405 10121
rect 16347 10112 16359 10115
rect 15856 10084 16359 10112
rect 16347 10081 16359 10084
rect 16393 10081 16405 10115
rect 16347 10075 16405 10081
rect 16482 10072 16488 10124
rect 16540 10072 16546 10124
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16724 10084 16773 10112
rect 16724 10072 16730 10084
rect 16761 10081 16773 10084
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 17218 10072 17224 10124
rect 17276 10072 17282 10124
rect 17586 10072 17592 10124
rect 17644 10072 17650 10124
rect 17696 10112 17724 10220
rect 19610 10208 19616 10260
rect 19668 10208 19674 10260
rect 20533 10251 20591 10257
rect 20533 10217 20545 10251
rect 20579 10248 20591 10251
rect 20898 10248 20904 10260
rect 20579 10220 20904 10248
rect 20579 10217 20591 10220
rect 20533 10211 20591 10217
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 23014 10208 23020 10260
rect 23072 10208 23078 10260
rect 25130 10208 25136 10260
rect 25188 10248 25194 10260
rect 26513 10251 26571 10257
rect 26513 10248 26525 10251
rect 25188 10220 26525 10248
rect 25188 10208 25194 10220
rect 26513 10217 26525 10220
rect 26559 10217 26571 10251
rect 26513 10211 26571 10217
rect 28534 10208 28540 10260
rect 28592 10208 28598 10260
rect 29270 10208 29276 10260
rect 29328 10208 29334 10260
rect 31726 10220 34192 10248
rect 20349 10183 20407 10189
rect 20349 10149 20361 10183
rect 20395 10180 20407 10183
rect 20714 10180 20720 10192
rect 20395 10152 20720 10180
rect 20395 10149 20407 10152
rect 20349 10143 20407 10149
rect 20714 10140 20720 10152
rect 20772 10180 20778 10192
rect 21450 10180 21456 10192
rect 20772 10152 21456 10180
rect 20772 10140 20778 10152
rect 21008 10121 21036 10152
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 21545 10183 21603 10189
rect 21545 10149 21557 10183
rect 21591 10180 21603 10183
rect 21591 10152 22968 10180
rect 21591 10149 21603 10152
rect 21545 10143 21603 10149
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 17696 10084 18061 10112
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 21085 10115 21143 10121
rect 21085 10081 21097 10115
rect 21131 10112 21143 10115
rect 22094 10112 22100 10124
rect 21131 10084 22100 10112
rect 21131 10081 21143 10084
rect 21085 10075 21143 10081
rect 22066 10072 22100 10084
rect 22152 10072 22158 10124
rect 22940 10121 22968 10152
rect 22925 10115 22983 10121
rect 22925 10081 22937 10115
rect 22971 10081 22983 10115
rect 22925 10075 22983 10081
rect 14507 10016 15424 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 8904 9948 9413 9976
rect 8904 9936 8910 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 10042 9976 10048 9988
rect 9401 9939 9459 9945
rect 9600 9948 10048 9976
rect 9600 9908 9628 9948
rect 10042 9936 10048 9948
rect 10100 9976 10106 9988
rect 10321 9979 10379 9985
rect 10321 9976 10333 9979
rect 10100 9948 10333 9976
rect 10100 9936 10106 9948
rect 10321 9945 10333 9948
rect 10367 9976 10379 9979
rect 13814 9976 13820 9988
rect 10367 9948 13820 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 13814 9936 13820 9948
rect 13872 9976 13878 9988
rect 15286 9976 15292 9988
rect 13872 9948 15292 9976
rect 13872 9936 13878 9948
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 15344 9948 15393 9976
rect 15344 9936 15350 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 17236 9976 17264 10072
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17604 10044 17632 10072
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 17451 10016 17632 10044
rect 17696 10016 18889 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17696 9976 17724 10016
rect 18877 10013 18889 10016
rect 18923 10013 18935 10047
rect 21450 10044 21456 10056
rect 18877 10007 18935 10013
rect 20640 10016 21456 10044
rect 17236 9948 17724 9976
rect 15381 9939 15439 9945
rect 17770 9936 17776 9988
rect 17828 9936 17834 9988
rect 20640 9985 20668 10016
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 17865 9979 17923 9985
rect 17865 9945 17877 9979
rect 17911 9976 17923 9979
rect 18325 9979 18383 9985
rect 18325 9976 18337 9979
rect 17911 9948 18337 9976
rect 17911 9945 17923 9948
rect 17865 9939 17923 9945
rect 18325 9945 18337 9948
rect 18371 9945 18383 9979
rect 18325 9939 18383 9945
rect 20625 9979 20683 9985
rect 20625 9945 20637 9979
rect 20671 9945 20683 9979
rect 20625 9939 20683 9945
rect 21177 9979 21235 9985
rect 21177 9945 21189 9979
rect 21223 9976 21235 9979
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21223 9948 21649 9976
rect 21223 9945 21235 9948
rect 21177 9939 21235 9945
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 22066 9976 22094 10072
rect 22278 10004 22284 10056
rect 22336 10004 22342 10056
rect 23032 10044 23060 10208
rect 25222 10180 25228 10192
rect 23952 10152 25228 10180
rect 23952 10121 23980 10152
rect 25222 10140 25228 10152
rect 25280 10140 25286 10192
rect 25317 10183 25375 10189
rect 25317 10149 25329 10183
rect 25363 10180 25375 10183
rect 26878 10180 26884 10192
rect 25363 10152 26884 10180
rect 25363 10149 25375 10152
rect 25317 10143 25375 10149
rect 26878 10140 26884 10152
rect 26936 10140 26942 10192
rect 27982 10140 27988 10192
rect 28040 10180 28046 10192
rect 28040 10152 29132 10180
rect 28040 10140 28046 10152
rect 29104 10124 29132 10152
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10112 24823 10115
rect 24854 10112 24860 10124
rect 24811 10084 24860 10112
rect 24811 10081 24823 10084
rect 24765 10075 24823 10081
rect 24854 10072 24860 10084
rect 24912 10112 24918 10124
rect 25593 10115 25651 10121
rect 25593 10112 25605 10115
rect 24912 10084 25605 10112
rect 24912 10072 24918 10084
rect 25593 10081 25605 10084
rect 25639 10112 25651 10115
rect 25639 10084 29040 10112
rect 25639 10081 25651 10084
rect 25593 10075 25651 10081
rect 24949 10047 25007 10053
rect 24949 10044 24961 10047
rect 23032 10016 24961 10044
rect 24949 10013 24961 10016
rect 24995 10013 25007 10047
rect 24949 10007 25007 10013
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10044 26755 10047
rect 27062 10044 27068 10056
rect 26743 10016 27068 10044
rect 26743 10013 26755 10016
rect 26697 10007 26755 10013
rect 27062 10004 27068 10016
rect 27120 10004 27126 10056
rect 29012 10044 29040 10084
rect 29086 10072 29092 10124
rect 29144 10072 29150 10124
rect 29288 10112 29316 10208
rect 31726 10124 31754 10220
rect 30101 10115 30159 10121
rect 30101 10112 30113 10115
rect 29288 10084 30113 10112
rect 30101 10081 30113 10084
rect 30147 10112 30159 10115
rect 30926 10112 30932 10124
rect 30147 10084 30932 10112
rect 30147 10081 30159 10084
rect 30101 10075 30159 10081
rect 30926 10072 30932 10084
rect 30984 10072 30990 10124
rect 31726 10072 31760 10124
rect 31812 10072 31818 10124
rect 31726 10044 31754 10072
rect 33321 10047 33379 10053
rect 33321 10044 33333 10047
rect 29012 10016 31754 10044
rect 31864 10016 33333 10044
rect 23661 9979 23719 9985
rect 23661 9976 23673 9979
rect 22066 9948 23673 9976
rect 21637 9939 21695 9945
rect 23661 9945 23673 9948
rect 23707 9976 23719 9979
rect 24302 9976 24308 9988
rect 23707 9948 24308 9976
rect 23707 9945 23719 9948
rect 23661 9939 23719 9945
rect 24302 9936 24308 9948
rect 24360 9976 24366 9988
rect 25682 9976 25688 9988
rect 24360 9948 25688 9976
rect 24360 9936 24366 9948
rect 25682 9936 25688 9948
rect 25740 9936 25746 9988
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 29549 9979 29607 9985
rect 29549 9976 29561 9979
rect 28951 9948 29561 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 29549 9945 29561 9948
rect 29595 9945 29607 9979
rect 29549 9939 29607 9945
rect 8352 9880 9628 9908
rect 8352 9868 8358 9880
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9732 9880 9965 9908
rect 9732 9868 9738 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 9953 9871 10011 9877
rect 12250 9868 12256 9920
rect 12308 9868 12314 9920
rect 15565 9911 15623 9917
rect 15565 9877 15577 9911
rect 15611 9908 15623 9911
rect 17034 9908 17040 9920
rect 15611 9880 17040 9908
rect 15611 9877 15623 9880
rect 15565 9871 15623 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 17494 9868 17500 9920
rect 17552 9868 17558 9920
rect 17788 9908 17816 9936
rect 31864 9920 31892 10016
rect 33321 10013 33333 10016
rect 33367 10044 33379 10047
rect 33410 10044 33416 10056
rect 33367 10016 33416 10044
rect 33367 10013 33379 10016
rect 33321 10007 33379 10013
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33502 10004 33508 10056
rect 33560 10044 33566 10056
rect 33965 10047 34023 10053
rect 33965 10044 33977 10047
rect 33560 10016 33977 10044
rect 33560 10004 33566 10016
rect 33965 10013 33977 10016
rect 34011 10013 34023 10047
rect 33965 10007 34023 10013
rect 33076 9979 33134 9985
rect 33076 9945 33088 9979
rect 33122 9976 33134 9979
rect 34164 9976 34192 10220
rect 35802 10208 35808 10260
rect 35860 10208 35866 10260
rect 36541 10251 36599 10257
rect 36541 10217 36553 10251
rect 36587 10248 36599 10251
rect 36814 10248 36820 10260
rect 36587 10220 36820 10248
rect 36587 10217 36599 10220
rect 36541 10211 36599 10217
rect 36814 10208 36820 10220
rect 36872 10208 36878 10260
rect 37458 10208 37464 10260
rect 37516 10248 37522 10260
rect 39393 10251 39451 10257
rect 39393 10248 39405 10251
rect 37516 10220 39405 10248
rect 37516 10208 37522 10220
rect 39393 10217 39405 10220
rect 39439 10217 39451 10251
rect 44450 10248 44456 10260
rect 39393 10211 39451 10217
rect 42352 10220 44456 10248
rect 37642 10140 37648 10192
rect 37700 10140 37706 10192
rect 38381 10183 38439 10189
rect 38381 10149 38393 10183
rect 38427 10149 38439 10183
rect 38381 10143 38439 10149
rect 36354 10072 36360 10124
rect 36412 10072 36418 10124
rect 36722 10072 36728 10124
rect 36780 10112 36786 10124
rect 37093 10115 37151 10121
rect 37093 10112 37105 10115
rect 36780 10084 37105 10112
rect 36780 10072 36786 10084
rect 37093 10081 37105 10084
rect 37139 10081 37151 10115
rect 37093 10075 37151 10081
rect 38289 10115 38347 10121
rect 38289 10081 38301 10115
rect 38335 10112 38347 10115
rect 38396 10112 38424 10143
rect 39850 10140 39856 10192
rect 39908 10140 39914 10192
rect 41248 10152 41368 10180
rect 41248 10124 41276 10152
rect 38335 10084 38424 10112
rect 38335 10081 38347 10084
rect 38289 10075 38347 10081
rect 38838 10072 38844 10124
rect 38896 10112 38902 10124
rect 38933 10115 38991 10121
rect 38933 10112 38945 10115
rect 38896 10084 38945 10112
rect 38896 10072 38902 10084
rect 38933 10081 38945 10084
rect 38979 10081 38991 10115
rect 38933 10075 38991 10081
rect 41230 10072 41236 10124
rect 41288 10072 41294 10124
rect 41340 10121 41368 10152
rect 41325 10115 41383 10121
rect 41325 10081 41337 10115
rect 41371 10081 41383 10115
rect 41325 10075 41383 10081
rect 38746 10004 38752 10056
rect 38804 10004 38810 10056
rect 42352 10044 42380 10220
rect 44450 10208 44456 10220
rect 44508 10208 44514 10260
rect 46198 10248 46204 10260
rect 45940 10220 46204 10248
rect 42705 10183 42763 10189
rect 42705 10149 42717 10183
rect 42751 10149 42763 10183
rect 42705 10143 42763 10149
rect 42720 10112 42748 10143
rect 43438 10112 43444 10124
rect 42720 10084 43444 10112
rect 43438 10072 43444 10084
rect 43496 10112 43502 10124
rect 43763 10115 43821 10121
rect 43763 10112 43775 10115
rect 43496 10084 43775 10112
rect 43496 10072 43502 10084
rect 43763 10081 43775 10084
rect 43809 10081 43821 10115
rect 43763 10075 43821 10081
rect 43898 10072 43904 10124
rect 43956 10072 43962 10124
rect 44174 10072 44180 10124
rect 44232 10072 44238 10124
rect 44821 10115 44879 10121
rect 44821 10081 44833 10115
rect 44867 10112 44879 10115
rect 45646 10112 45652 10124
rect 44867 10084 45652 10112
rect 44867 10081 44879 10084
rect 44821 10075 44879 10081
rect 45646 10072 45652 10084
rect 45704 10072 45710 10124
rect 40880 10016 42380 10044
rect 40880 9976 40908 10016
rect 43622 10004 43628 10056
rect 43680 10004 43686 10056
rect 44634 10004 44640 10056
rect 44692 10004 44698 10056
rect 45940 10053 45968 10220
rect 46198 10208 46204 10220
rect 46256 10208 46262 10260
rect 49602 10208 49608 10260
rect 49660 10208 49666 10260
rect 49970 10208 49976 10260
rect 50028 10208 50034 10260
rect 51350 10208 51356 10260
rect 51408 10248 51414 10260
rect 51629 10251 51687 10257
rect 51629 10248 51641 10251
rect 51408 10220 51641 10248
rect 51408 10208 51414 10220
rect 51629 10217 51641 10220
rect 51675 10217 51687 10251
rect 51629 10211 51687 10217
rect 53285 10251 53343 10257
rect 53285 10217 53297 10251
rect 53331 10248 53343 10251
rect 53834 10248 53840 10260
rect 53331 10220 53840 10248
rect 53331 10217 53343 10220
rect 53285 10211 53343 10217
rect 53834 10208 53840 10220
rect 53892 10208 53898 10260
rect 54849 10251 54907 10257
rect 54849 10217 54861 10251
rect 54895 10248 54907 10251
rect 55030 10248 55036 10260
rect 54895 10220 55036 10248
rect 54895 10217 54907 10220
rect 54849 10211 54907 10217
rect 55030 10208 55036 10220
rect 55088 10208 55094 10260
rect 56686 10208 56692 10260
rect 56744 10248 56750 10260
rect 57701 10251 57759 10257
rect 57701 10248 57713 10251
rect 56744 10220 57713 10248
rect 56744 10208 56750 10220
rect 57701 10217 57713 10220
rect 57747 10217 57759 10251
rect 57701 10211 57759 10217
rect 57882 10208 57888 10260
rect 57940 10208 57946 10260
rect 47857 10183 47915 10189
rect 47857 10149 47869 10183
rect 47903 10180 47915 10183
rect 48406 10180 48412 10192
rect 47903 10152 48412 10180
rect 47903 10149 47915 10152
rect 47857 10143 47915 10149
rect 48406 10140 48412 10152
rect 48464 10180 48470 10192
rect 49620 10180 49648 10208
rect 48464 10152 49648 10180
rect 48464 10140 48470 10152
rect 48961 10115 49019 10121
rect 48961 10081 48973 10115
rect 49007 10112 49019 10115
rect 49988 10112 50016 10208
rect 52270 10140 52276 10192
rect 52328 10180 52334 10192
rect 52825 10183 52883 10189
rect 52825 10180 52837 10183
rect 52328 10152 52837 10180
rect 52328 10140 52334 10152
rect 52825 10149 52837 10152
rect 52871 10180 52883 10183
rect 52871 10152 54340 10180
rect 52871 10149 52883 10152
rect 52825 10143 52883 10149
rect 49007 10084 50016 10112
rect 51537 10115 51595 10121
rect 49007 10081 49019 10084
rect 48961 10075 49019 10081
rect 51537 10081 51549 10115
rect 51583 10112 51595 10115
rect 52454 10112 52460 10124
rect 51583 10084 52460 10112
rect 51583 10081 51595 10084
rect 51537 10075 51595 10081
rect 45925 10047 45983 10053
rect 45925 10013 45937 10047
rect 45971 10013 45983 10047
rect 45925 10007 45983 10013
rect 46477 10047 46535 10053
rect 46477 10013 46489 10047
rect 46523 10013 46535 10047
rect 46477 10007 46535 10013
rect 33122 9948 33456 9976
rect 34164 9948 40908 9976
rect 40988 9979 41046 9985
rect 33122 9945 33134 9948
rect 33076 9939 33134 9945
rect 17957 9911 18015 9917
rect 17957 9908 17969 9911
rect 17788 9880 17969 9908
rect 17957 9877 17969 9880
rect 18003 9877 18015 9911
rect 17957 9871 18015 9877
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 22373 9911 22431 9917
rect 22373 9908 22385 9911
rect 21416 9880 22385 9908
rect 21416 9868 21422 9880
rect 22373 9877 22385 9880
rect 22419 9877 22431 9911
rect 22373 9871 22431 9877
rect 23293 9911 23351 9917
rect 23293 9877 23305 9911
rect 23339 9908 23351 9911
rect 23566 9908 23572 9920
rect 23339 9880 23572 9908
rect 23339 9877 23351 9880
rect 23293 9871 23351 9877
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 23750 9868 23756 9920
rect 23808 9868 23814 9920
rect 24394 9868 24400 9920
rect 24452 9908 24458 9920
rect 24857 9911 24915 9917
rect 24857 9908 24869 9911
rect 24452 9880 24869 9908
rect 24452 9868 24458 9880
rect 24857 9877 24869 9880
rect 24903 9877 24915 9911
rect 24857 9871 24915 9877
rect 27706 9868 27712 9920
rect 27764 9908 27770 9920
rect 27985 9911 28043 9917
rect 27985 9908 27997 9911
rect 27764 9880 27997 9908
rect 27764 9868 27770 9880
rect 27985 9877 27997 9880
rect 28031 9908 28043 9911
rect 28074 9908 28080 9920
rect 28031 9880 28080 9908
rect 28031 9877 28043 9880
rect 27985 9871 28043 9877
rect 28074 9868 28080 9880
rect 28132 9868 28138 9920
rect 28810 9868 28816 9920
rect 28868 9908 28874 9920
rect 28997 9911 29055 9917
rect 28997 9908 29009 9911
rect 28868 9880 29009 9908
rect 28868 9868 28874 9880
rect 28997 9877 29009 9880
rect 29043 9877 29055 9911
rect 28997 9871 29055 9877
rect 29086 9868 29092 9920
rect 29144 9908 29150 9920
rect 30469 9911 30527 9917
rect 30469 9908 30481 9911
rect 29144 9880 30481 9908
rect 29144 9868 29150 9880
rect 30469 9877 30481 9880
rect 30515 9877 30527 9911
rect 30469 9871 30527 9877
rect 30558 9868 30564 9920
rect 30616 9908 30622 9920
rect 31389 9911 31447 9917
rect 31389 9908 31401 9911
rect 30616 9880 31401 9908
rect 30616 9868 30622 9880
rect 31389 9877 31401 9880
rect 31435 9877 31447 9911
rect 31389 9871 31447 9877
rect 31846 9868 31852 9920
rect 31904 9868 31910 9920
rect 31938 9868 31944 9920
rect 31996 9908 32002 9920
rect 33226 9908 33232 9920
rect 31996 9880 33232 9908
rect 31996 9868 32002 9880
rect 33226 9868 33232 9880
rect 33284 9868 33290 9920
rect 33428 9917 33456 9948
rect 40988 9945 41000 9979
rect 41034 9976 41046 9979
rect 41138 9976 41144 9988
rect 41034 9948 41144 9976
rect 41034 9945 41046 9948
rect 40988 9939 41046 9945
rect 41138 9936 41144 9948
rect 41196 9936 41202 9988
rect 41598 9985 41604 9988
rect 41592 9939 41604 9985
rect 41598 9936 41604 9939
rect 41656 9936 41662 9988
rect 44818 9936 44824 9988
rect 44876 9976 44882 9988
rect 45097 9979 45155 9985
rect 45097 9976 45109 9979
rect 44876 9948 45109 9976
rect 44876 9936 44882 9948
rect 45097 9945 45109 9948
rect 45143 9945 45155 9979
rect 45097 9939 45155 9945
rect 45830 9936 45836 9988
rect 45888 9976 45894 9988
rect 46492 9976 46520 10007
rect 48314 10004 48320 10056
rect 48372 10044 48378 10056
rect 48501 10047 48559 10053
rect 48501 10044 48513 10047
rect 48372 10016 48513 10044
rect 48372 10004 48378 10016
rect 48501 10013 48513 10016
rect 48547 10013 48559 10047
rect 48501 10007 48559 10013
rect 49605 10047 49663 10053
rect 49605 10013 49617 10047
rect 49651 10044 49663 10047
rect 49878 10044 49884 10056
rect 49651 10016 49884 10044
rect 49651 10013 49663 10016
rect 49605 10007 49663 10013
rect 49878 10004 49884 10016
rect 49936 10004 49942 10056
rect 51552 10044 51580 10075
rect 52454 10072 52460 10084
rect 52512 10072 52518 10124
rect 54312 10121 54340 10152
rect 53837 10115 53895 10121
rect 53837 10112 53849 10115
rect 53116 10084 53849 10112
rect 49988 10016 51580 10044
rect 52181 10047 52239 10053
rect 45888 9948 46520 9976
rect 45888 9936 45894 9948
rect 33413 9911 33471 9917
rect 33413 9877 33425 9911
rect 33459 9877 33471 9911
rect 33413 9871 33471 9877
rect 38841 9911 38899 9917
rect 38841 9877 38853 9911
rect 38887 9908 38899 9911
rect 38930 9908 38936 9920
rect 38887 9880 38936 9908
rect 38887 9877 38899 9880
rect 38841 9871 38899 9877
rect 38930 9868 38936 9880
rect 38988 9908 38994 9920
rect 39298 9908 39304 9920
rect 38988 9880 39304 9908
rect 38988 9868 38994 9880
rect 39298 9868 39304 9880
rect 39356 9868 39362 9920
rect 42981 9911 43039 9917
rect 42981 9877 42993 9911
rect 43027 9908 43039 9911
rect 45462 9908 45468 9920
rect 43027 9880 45468 9908
rect 43027 9877 43039 9880
rect 42981 9871 43039 9877
rect 45462 9868 45468 9880
rect 45520 9868 45526 9920
rect 46492 9908 46520 9948
rect 46744 9979 46802 9985
rect 46744 9945 46756 9979
rect 46790 9976 46802 9979
rect 47949 9979 48007 9985
rect 47949 9976 47961 9979
rect 46790 9948 47961 9976
rect 46790 9945 46802 9948
rect 46744 9939 46802 9945
rect 47949 9945 47961 9948
rect 47995 9945 48007 9979
rect 47949 9939 48007 9945
rect 49418 9936 49424 9988
rect 49476 9936 49482 9988
rect 49988 9920 50016 10016
rect 52181 10013 52193 10047
rect 52227 10013 52239 10047
rect 52181 10007 52239 10013
rect 51292 9979 51350 9985
rect 51292 9945 51304 9979
rect 51338 9976 51350 9979
rect 51810 9976 51816 9988
rect 51338 9948 51816 9976
rect 51338 9945 51350 9948
rect 51292 9939 51350 9945
rect 51810 9936 51816 9948
rect 51868 9936 51874 9988
rect 49970 9908 49976 9920
rect 46492 9880 49976 9908
rect 49970 9868 49976 9880
rect 50028 9868 50034 9920
rect 50157 9911 50215 9917
rect 50157 9877 50169 9911
rect 50203 9908 50215 9911
rect 50522 9908 50528 9920
rect 50203 9880 50528 9908
rect 50203 9877 50215 9880
rect 50157 9871 50215 9877
rect 50522 9868 50528 9880
rect 50580 9908 50586 9920
rect 52196 9908 52224 10007
rect 50580 9880 52224 9908
rect 50580 9868 50586 9880
rect 52638 9868 52644 9920
rect 52696 9908 52702 9920
rect 53116 9917 53144 10084
rect 53837 10081 53849 10084
rect 53883 10081 53895 10115
rect 53837 10075 53895 10081
rect 54297 10115 54355 10121
rect 54297 10081 54309 10115
rect 54343 10112 54355 10115
rect 54386 10112 54392 10124
rect 54343 10084 54392 10112
rect 54343 10081 54355 10084
rect 54297 10075 54355 10081
rect 54386 10072 54392 10084
rect 54444 10072 54450 10124
rect 55398 10072 55404 10124
rect 55456 10112 55462 10124
rect 55861 10115 55919 10121
rect 55861 10112 55873 10115
rect 55456 10084 55873 10112
rect 55456 10072 55462 10084
rect 55861 10081 55873 10084
rect 55907 10081 55919 10115
rect 57900 10112 57928 10208
rect 55861 10075 55919 10081
rect 57532 10084 57928 10112
rect 57353 10047 57411 10053
rect 57353 10013 57365 10047
rect 57399 10044 57411 10047
rect 57532 10044 57560 10084
rect 57399 10016 57560 10044
rect 57609 10047 57667 10053
rect 57399 10013 57411 10016
rect 57353 10007 57411 10013
rect 57609 10013 57621 10047
rect 57655 10044 57667 10047
rect 57698 10044 57704 10056
rect 57655 10016 57704 10044
rect 57655 10013 57667 10016
rect 57609 10007 57667 10013
rect 57698 10004 57704 10016
rect 57756 10004 57762 10056
rect 58253 10047 58311 10053
rect 58253 10013 58265 10047
rect 58299 10013 58311 10047
rect 58253 10007 58311 10013
rect 53653 9979 53711 9985
rect 53653 9945 53665 9979
rect 53699 9976 53711 9979
rect 54018 9976 54024 9988
rect 53699 9948 54024 9976
rect 53699 9945 53711 9948
rect 53653 9939 53711 9945
rect 54018 9936 54024 9948
rect 54076 9936 54082 9988
rect 54389 9979 54447 9985
rect 54389 9945 54401 9979
rect 54435 9976 54447 9979
rect 55309 9979 55367 9985
rect 55309 9976 55321 9979
rect 54435 9948 55321 9976
rect 54435 9945 54447 9948
rect 54389 9939 54447 9945
rect 55309 9945 55321 9948
rect 55355 9945 55367 9979
rect 55309 9939 55367 9945
rect 53101 9911 53159 9917
rect 53101 9908 53113 9911
rect 52696 9880 53113 9908
rect 52696 9868 52702 9880
rect 53101 9877 53113 9880
rect 53147 9877 53159 9911
rect 53101 9871 53159 9877
rect 53745 9911 53803 9917
rect 53745 9877 53757 9911
rect 53791 9908 53803 9911
rect 54110 9908 54116 9920
rect 53791 9880 54116 9908
rect 53791 9877 53803 9880
rect 53745 9871 53803 9877
rect 54110 9868 54116 9880
rect 54168 9908 54174 9920
rect 54481 9911 54539 9917
rect 54481 9908 54493 9911
rect 54168 9880 54493 9908
rect 54168 9868 54174 9880
rect 54481 9877 54493 9880
rect 54527 9877 54539 9911
rect 54481 9871 54539 9877
rect 56229 9911 56287 9917
rect 56229 9877 56241 9911
rect 56275 9908 56287 9911
rect 56318 9908 56324 9920
rect 56275 9880 56324 9908
rect 56275 9877 56287 9880
rect 56229 9871 56287 9877
rect 56318 9868 56324 9880
rect 56376 9908 56382 9920
rect 58268 9908 58296 10007
rect 56376 9880 58296 9908
rect 56376 9868 56382 9880
rect 1104 9818 59040 9840
rect 1104 9766 15394 9818
rect 15446 9766 15458 9818
rect 15510 9766 15522 9818
rect 15574 9766 15586 9818
rect 15638 9766 15650 9818
rect 15702 9766 29838 9818
rect 29890 9766 29902 9818
rect 29954 9766 29966 9818
rect 30018 9766 30030 9818
rect 30082 9766 30094 9818
rect 30146 9766 44282 9818
rect 44334 9766 44346 9818
rect 44398 9766 44410 9818
rect 44462 9766 44474 9818
rect 44526 9766 44538 9818
rect 44590 9766 58726 9818
rect 58778 9766 58790 9818
rect 58842 9766 58854 9818
rect 58906 9766 58918 9818
rect 58970 9766 58982 9818
rect 59034 9766 59040 9818
rect 1104 9744 59040 9766
rect 3050 9664 3056 9716
rect 3108 9664 3114 9716
rect 8662 9704 8668 9716
rect 8220 9676 8668 9704
rect 2222 9596 2228 9648
rect 2280 9636 2286 9648
rect 3234 9636 3240 9648
rect 2280 9608 3240 9636
rect 2280 9596 2286 9608
rect 3234 9596 3240 9608
rect 3292 9636 3298 9648
rect 3292 9608 4016 9636
rect 3292 9596 3298 9608
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 3878 9568 3884 9580
rect 3835 9540 3884 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 3988 9577 4016 9608
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4120 9608 4629 9636
rect 4120 9596 4126 9608
rect 4617 9605 4629 9608
rect 4663 9605 4675 9639
rect 4617 9599 4675 9605
rect 4908 9608 5488 9636
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4908 9568 4936 9608
rect 5460 9580 5488 9608
rect 6730 9596 6736 9648
rect 6788 9596 6794 9648
rect 7650 9596 7656 9648
rect 7708 9636 7714 9648
rect 8220 9645 8248 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 9122 9664 9128 9716
rect 9180 9664 9186 9716
rect 12253 9707 12311 9713
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 12802 9704 12808 9716
rect 12299 9676 12808 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 19610 9664 19616 9716
rect 19668 9664 19674 9716
rect 22094 9664 22100 9716
rect 22152 9664 22158 9716
rect 32953 9707 33011 9713
rect 32953 9673 32965 9707
rect 32999 9704 33011 9707
rect 33502 9704 33508 9716
rect 32999 9676 33508 9704
rect 32999 9673 33011 9676
rect 32953 9667 33011 9673
rect 33502 9664 33508 9676
rect 33560 9664 33566 9716
rect 33686 9664 33692 9716
rect 33744 9664 33750 9716
rect 41138 9664 41144 9716
rect 41196 9664 41202 9716
rect 41598 9664 41604 9716
rect 41656 9664 41662 9716
rect 42426 9664 42432 9716
rect 42484 9704 42490 9716
rect 43441 9707 43499 9713
rect 43441 9704 43453 9707
rect 42484 9676 43453 9704
rect 42484 9664 42490 9676
rect 43441 9673 43453 9676
rect 43487 9704 43499 9707
rect 43530 9704 43536 9716
rect 43487 9676 43536 9704
rect 43487 9673 43499 9676
rect 43441 9667 43499 9673
rect 43530 9664 43536 9676
rect 43588 9664 43594 9716
rect 45462 9664 45468 9716
rect 45520 9664 45526 9716
rect 48774 9704 48780 9716
rect 46768 9676 48780 9704
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7708 9608 7849 9636
rect 7708 9596 7714 9608
rect 7837 9605 7849 9608
rect 7883 9636 7895 9639
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7883 9608 8217 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 9140 9636 9168 9664
rect 8588 9608 9168 9636
rect 9217 9639 9275 9645
rect 4387 9540 4936 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 3988 9432 4016 9531
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5368 9500 5396 9531
rect 5442 9528 5448 9580
rect 5500 9528 5506 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5684 9540 6561 9568
rect 5684 9528 5690 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 7926 9528 7932 9580
rect 7984 9528 7990 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8312 9568 8340 9596
rect 8588 9577 8616 9608
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 9490 9636 9496 9648
rect 9263 9608 9496 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 12621 9639 12679 9645
rect 12621 9605 12633 9639
rect 12667 9636 12679 9639
rect 14185 9639 14243 9645
rect 14185 9636 14197 9639
rect 12667 9608 14197 9636
rect 12667 9605 12679 9608
rect 12621 9599 12679 9605
rect 14185 9605 14197 9608
rect 14231 9605 14243 9639
rect 14185 9599 14243 9605
rect 15378 9596 15384 9648
rect 15436 9636 15442 9648
rect 16206 9636 16212 9648
rect 15436 9608 16212 9636
rect 15436 9596 15442 9608
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18141 9639 18199 9645
rect 18141 9636 18153 9639
rect 18104 9608 18153 9636
rect 18104 9596 18110 9608
rect 18141 9605 18153 9608
rect 18187 9605 18199 9639
rect 18141 9599 18199 9605
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9636 18567 9639
rect 19628 9636 19656 9664
rect 20432 9639 20490 9645
rect 18555 9608 20208 9636
rect 18555 9605 18567 9608
rect 18509 9599 18567 9605
rect 8021 9531 8079 9537
rect 8128 9540 8340 9568
rect 8573 9571 8631 9577
rect 5534 9500 5540 9512
rect 5368 9472 5540 9500
rect 5534 9460 5540 9472
rect 5592 9500 5598 9512
rect 7116 9500 7144 9528
rect 7742 9500 7748 9512
rect 5592 9472 6132 9500
rect 7116 9472 7748 9500
rect 5592 9460 5598 9472
rect 6104 9441 6132 9472
rect 7742 9460 7748 9472
rect 7800 9500 7806 9512
rect 8036 9500 8064 9531
rect 7800 9472 8064 9500
rect 7800 9460 7806 9472
rect 6089 9435 6147 9441
rect 3988 9404 4568 9432
rect 4540 9376 4568 9404
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6178 9432 6184 9444
rect 6135 9404 6184 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 6178 9392 6184 9404
rect 6236 9432 6242 9444
rect 8128 9432 8156 9540
rect 8573 9537 8585 9571
rect 8619 9537 8631 9571
rect 10606 9571 10664 9577
rect 10606 9568 10618 9571
rect 8573 9531 8631 9537
rect 8772 9540 10618 9568
rect 6236 9404 8156 9432
rect 8205 9435 8263 9441
rect 6236 9392 6242 9404
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8665 9435 8723 9441
rect 8665 9432 8677 9435
rect 8251 9404 8677 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8665 9401 8677 9404
rect 8711 9401 8723 9435
rect 8665 9395 8723 9401
rect 4522 9324 4528 9376
rect 4580 9324 4586 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 8772 9373 8800 9540
rect 10606 9537 10618 9540
rect 10652 9537 10664 9571
rect 10606 9531 10664 9537
rect 12084 9540 12848 9568
rect 12084 9512 12112 9540
rect 8846 9460 8852 9512
rect 8904 9460 8910 9512
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 9272 9472 9536 9500
rect 9272 9460 9278 9472
rect 9508 9441 9536 9472
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11882 9500 11888 9512
rect 10928 9472 11888 9500
rect 10928 9460 10934 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 12066 9460 12072 9512
rect 12124 9460 12130 9512
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 12820 9509 12848 9540
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 13044 9540 13093 9568
rect 13044 9528 13050 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16080 9540 16804 9568
rect 16080 9528 16086 9540
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 12851 9472 13461 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16666 9500 16672 9512
rect 15344 9472 16672 9500
rect 15344 9460 15350 9472
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16776 9509 16804 9540
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 20180 9577 20208 9608
rect 20432 9605 20444 9639
rect 20478 9636 20490 9639
rect 21358 9636 21364 9648
rect 20478 9608 21364 9636
rect 20478 9605 20490 9608
rect 20432 9599 20490 9605
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 22112 9636 22140 9664
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 22112 9608 22201 9636
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 22189 9599 22247 9605
rect 28074 9596 28080 9648
rect 28132 9596 28138 9648
rect 28537 9639 28595 9645
rect 28537 9605 28549 9639
rect 28583 9636 28595 9639
rect 28810 9636 28816 9648
rect 28583 9608 28816 9636
rect 28583 9605 28595 9608
rect 28537 9599 28595 9605
rect 28810 9596 28816 9608
rect 28868 9596 28874 9648
rect 30834 9636 30840 9648
rect 29656 9608 30840 9636
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 23474 9528 23480 9580
rect 23532 9528 23538 9580
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9568 24547 9571
rect 24535 9540 24992 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 16942 9460 16948 9512
rect 17000 9460 17006 9512
rect 21910 9500 21916 9512
rect 21468 9472 21916 9500
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9401 9551 9435
rect 9493 9395 9551 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11793 9435 11851 9441
rect 11793 9432 11805 9435
rect 11112 9404 11805 9432
rect 11112 9392 11118 9404
rect 11793 9401 11805 9404
rect 11839 9432 11851 9435
rect 19242 9432 19248 9444
rect 11839 9404 19248 9432
rect 11839 9401 11851 9404
rect 11793 9395 11851 9401
rect 19242 9392 19248 9404
rect 19300 9392 19306 9444
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6880 9336 7021 9364
rect 6880 9324 6886 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 8757 9367 8815 9373
rect 8757 9333 8769 9367
rect 8803 9333 8815 9367
rect 8757 9327 8815 9333
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 13630 9364 13636 9376
rect 12400 9336 13636 9364
rect 12400 9324 12406 9336
rect 13630 9324 13636 9336
rect 13688 9364 13694 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 13688 9336 15577 9364
rect 13688 9324 13694 9336
rect 15565 9333 15577 9336
rect 15611 9364 15623 9367
rect 15930 9364 15936 9376
rect 15611 9336 15936 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16022 9324 16028 9376
rect 16080 9324 16086 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16393 9327 16451 9333
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17092 9336 17417 9364
rect 17092 9324 17098 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17405 9327 17463 9333
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 18656 9336 20085 9364
rect 18656 9324 18662 9336
rect 20073 9333 20085 9336
rect 20119 9364 20131 9367
rect 21468 9364 21496 9472
rect 21910 9460 21916 9472
rect 21968 9460 21974 9512
rect 22094 9460 22100 9512
rect 22152 9460 22158 9512
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 23615 9503 23673 9509
rect 23615 9500 23627 9503
rect 22336 9472 23627 9500
rect 22336 9460 22342 9472
rect 23615 9469 23627 9472
rect 23661 9469 23673 9503
rect 23615 9463 23673 9469
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9500 23811 9503
rect 23934 9500 23940 9512
rect 23799 9472 23940 9500
rect 23799 9469 23811 9472
rect 23753 9463 23811 9469
rect 23934 9460 23940 9472
rect 23992 9460 23998 9512
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9500 24087 9503
rect 24118 9500 24124 9512
rect 24075 9472 24124 9500
rect 24075 9469 24087 9472
rect 24029 9463 24087 9469
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 24394 9460 24400 9512
rect 24452 9460 24458 9512
rect 24673 9503 24731 9509
rect 24673 9469 24685 9503
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 21545 9435 21603 9441
rect 21545 9401 21557 9435
rect 21591 9432 21603 9435
rect 22296 9432 22324 9460
rect 21591 9404 22324 9432
rect 21591 9401 21603 9404
rect 21545 9395 21603 9401
rect 20119 9336 21496 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 22557 9367 22615 9373
rect 22557 9364 22569 9367
rect 22520 9336 22569 9364
rect 22520 9324 22526 9336
rect 22557 9333 22569 9336
rect 22603 9333 22615 9367
rect 22557 9327 22615 9333
rect 22833 9367 22891 9373
rect 22833 9333 22845 9367
rect 22879 9364 22891 9367
rect 24412 9364 24440 9460
rect 24688 9376 24716 9463
rect 22879 9336 24440 9364
rect 22879 9333 22891 9336
rect 22833 9327 22891 9333
rect 24670 9324 24676 9376
rect 24728 9324 24734 9376
rect 24964 9373 24992 9540
rect 26050 9528 26056 9580
rect 26108 9577 26114 9580
rect 26108 9531 26120 9577
rect 28092 9568 28120 9596
rect 29656 9577 29684 9608
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 31294 9596 31300 9648
rect 31352 9596 31358 9648
rect 32490 9596 32496 9648
rect 32548 9636 32554 9648
rect 33704 9636 33732 9664
rect 32548 9608 33732 9636
rect 32548 9596 32554 9608
rect 35894 9596 35900 9648
rect 35952 9636 35958 9648
rect 36357 9639 36415 9645
rect 36357 9636 36369 9639
rect 35952 9608 36369 9636
rect 35952 9596 35958 9608
rect 36357 9605 36369 9608
rect 36403 9605 36415 9639
rect 36357 9599 36415 9605
rect 36464 9608 38240 9636
rect 28629 9571 28687 9577
rect 28092 9540 28580 9568
rect 26108 9528 26114 9531
rect 28552 9512 28580 9540
rect 28629 9537 28641 9571
rect 28675 9568 28687 9571
rect 28997 9571 29055 9577
rect 28997 9568 29009 9571
rect 28675 9540 29009 9568
rect 28675 9537 28687 9540
rect 28629 9531 28687 9537
rect 28997 9537 29009 9540
rect 29043 9537 29055 9571
rect 28997 9531 29055 9537
rect 29641 9571 29699 9577
rect 29641 9537 29653 9571
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 30561 9571 30619 9577
rect 30561 9537 30573 9571
rect 30607 9568 30619 9571
rect 30742 9568 30748 9580
rect 30607 9540 30748 9568
rect 30607 9537 30619 9540
rect 30561 9531 30619 9537
rect 30742 9528 30748 9540
rect 30800 9528 30806 9580
rect 31846 9568 31852 9580
rect 30852 9540 31852 9568
rect 26329 9503 26387 9509
rect 26329 9469 26341 9503
rect 26375 9469 26387 9503
rect 26329 9463 26387 9469
rect 27433 9503 27491 9509
rect 27433 9469 27445 9503
rect 27479 9500 27491 9503
rect 27706 9500 27712 9512
rect 27479 9472 27712 9500
rect 27479 9469 27491 9472
rect 27433 9463 27491 9469
rect 26344 9432 26372 9463
rect 27706 9460 27712 9472
rect 27764 9460 27770 9512
rect 28077 9503 28135 9509
rect 28077 9469 28089 9503
rect 28123 9500 28135 9503
rect 28123 9472 28212 9500
rect 28123 9469 28135 9472
rect 28077 9463 28135 9469
rect 28184 9441 28212 9472
rect 28534 9460 28540 9512
rect 28592 9500 28598 9512
rect 28721 9503 28779 9509
rect 28721 9500 28733 9503
rect 28592 9472 28733 9500
rect 28592 9460 28598 9472
rect 28721 9469 28733 9472
rect 28767 9469 28779 9503
rect 28721 9463 28779 9469
rect 26697 9435 26755 9441
rect 26697 9432 26709 9435
rect 26344 9404 26709 9432
rect 26697 9401 26709 9404
rect 26743 9401 26755 9435
rect 26697 9395 26755 9401
rect 28169 9435 28227 9441
rect 28169 9401 28181 9435
rect 28215 9401 28227 9435
rect 30852 9432 30880 9540
rect 31846 9528 31852 9540
rect 31904 9528 31910 9580
rect 32585 9571 32643 9577
rect 32585 9537 32597 9571
rect 32631 9568 32643 9571
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32631 9540 33057 9568
rect 32631 9537 32643 9540
rect 32585 9531 32643 9537
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 33226 9528 33232 9580
rect 33284 9568 33290 9580
rect 33597 9571 33655 9577
rect 33597 9568 33609 9571
rect 33284 9540 33609 9568
rect 33284 9528 33290 9540
rect 33597 9537 33609 9540
rect 33643 9537 33655 9571
rect 33597 9531 33655 9537
rect 34057 9571 34115 9577
rect 34057 9537 34069 9571
rect 34103 9568 34115 9571
rect 34146 9568 34152 9580
rect 34103 9540 34152 9568
rect 34103 9537 34115 9540
rect 34057 9531 34115 9537
rect 32401 9503 32459 9509
rect 32401 9469 32413 9503
rect 32447 9500 32459 9503
rect 34072 9500 34100 9531
rect 34146 9528 34152 9540
rect 34204 9568 34210 9580
rect 36464 9568 36492 9608
rect 38212 9580 38240 9608
rect 39298 9596 39304 9648
rect 39356 9636 39362 9648
rect 39758 9636 39764 9648
rect 39356 9608 39764 9636
rect 39356 9596 39362 9608
rect 39758 9596 39764 9608
rect 39816 9596 39822 9648
rect 43622 9596 43628 9648
rect 43680 9636 43686 9648
rect 43680 9608 44128 9636
rect 43680 9596 43686 9608
rect 34204 9540 36492 9568
rect 36541 9571 36599 9577
rect 34204 9528 34210 9540
rect 36541 9537 36553 9571
rect 36587 9568 36599 9571
rect 36630 9568 36636 9580
rect 36587 9540 36636 9568
rect 36587 9537 36599 9540
rect 36541 9531 36599 9537
rect 36630 9528 36636 9540
rect 36688 9528 36694 9580
rect 38194 9528 38200 9580
rect 38252 9568 38258 9580
rect 38746 9568 38752 9580
rect 38252 9540 38752 9568
rect 38252 9528 38258 9540
rect 38746 9528 38752 9540
rect 38804 9528 38810 9580
rect 38838 9528 38844 9580
rect 38896 9528 38902 9580
rect 39850 9528 39856 9580
rect 39908 9568 39914 9580
rect 40313 9571 40371 9577
rect 40313 9568 40325 9571
rect 39908 9540 40325 9568
rect 39908 9528 39914 9540
rect 40313 9537 40325 9540
rect 40359 9537 40371 9571
rect 40313 9531 40371 9537
rect 42794 9528 42800 9580
rect 42852 9528 42858 9580
rect 42886 9528 42892 9580
rect 42944 9568 42950 9580
rect 42944 9540 43300 9568
rect 42944 9528 42950 9540
rect 32447 9472 34100 9500
rect 35345 9503 35403 9509
rect 32447 9469 32459 9472
rect 32401 9463 32459 9469
rect 35345 9469 35357 9503
rect 35391 9500 35403 9503
rect 36078 9500 36084 9512
rect 35391 9472 36084 9500
rect 35391 9469 35403 9472
rect 35345 9463 35403 9469
rect 36078 9460 36084 9472
rect 36136 9460 36142 9512
rect 37734 9460 37740 9512
rect 37792 9500 37798 9512
rect 39025 9503 39083 9509
rect 39025 9500 39037 9503
rect 37792 9472 39037 9500
rect 37792 9460 37798 9472
rect 28169 9395 28227 9401
rect 29932 9404 30880 9432
rect 24949 9367 25007 9373
rect 24949 9333 24961 9367
rect 24995 9364 25007 9367
rect 26602 9364 26608 9376
rect 24995 9336 26608 9364
rect 24995 9333 25007 9336
rect 24949 9327 25007 9333
rect 26602 9324 26608 9336
rect 26660 9324 26666 9376
rect 26712 9364 26740 9395
rect 27614 9364 27620 9376
rect 26712 9336 27620 9364
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 29454 9324 29460 9376
rect 29512 9364 29518 9376
rect 29932 9373 29960 9404
rect 29917 9367 29975 9373
rect 29917 9364 29929 9367
rect 29512 9336 29929 9364
rect 29512 9324 29518 9336
rect 29917 9333 29929 9336
rect 29963 9333 29975 9367
rect 29917 9327 29975 9333
rect 31846 9324 31852 9376
rect 31904 9364 31910 9376
rect 32398 9364 32404 9376
rect 31904 9336 32404 9364
rect 31904 9324 31910 9336
rect 32398 9324 32404 9336
rect 32456 9324 32462 9376
rect 34238 9324 34244 9376
rect 34296 9364 34302 9376
rect 34333 9367 34391 9373
rect 34333 9364 34345 9367
rect 34296 9336 34345 9364
rect 34296 9324 34302 9336
rect 34333 9333 34345 9336
rect 34379 9333 34391 9367
rect 34333 9327 34391 9333
rect 35894 9324 35900 9376
rect 35952 9324 35958 9376
rect 37458 9324 37464 9376
rect 37516 9364 37522 9376
rect 37844 9373 37872 9472
rect 39025 9469 39037 9472
rect 39071 9469 39083 9503
rect 39025 9463 39083 9469
rect 39209 9503 39267 9509
rect 39209 9469 39221 9503
rect 39255 9500 39267 9503
rect 39761 9503 39819 9509
rect 39761 9500 39773 9503
rect 39255 9472 39773 9500
rect 39255 9469 39267 9472
rect 39209 9463 39267 9469
rect 39761 9469 39773 9472
rect 39807 9469 39819 9503
rect 39761 9463 39819 9469
rect 40497 9503 40555 9509
rect 40497 9469 40509 9503
rect 40543 9469 40555 9503
rect 40497 9463 40555 9469
rect 42245 9503 42303 9509
rect 42245 9469 42257 9503
rect 42291 9500 42303 9503
rect 42981 9503 43039 9509
rect 42981 9500 42993 9503
rect 42291 9472 42472 9500
rect 42291 9469 42303 9472
rect 42245 9463 42303 9469
rect 38654 9392 38660 9444
rect 38712 9392 38718 9444
rect 39669 9435 39727 9441
rect 39669 9401 39681 9435
rect 39715 9432 39727 9435
rect 40512 9432 40540 9463
rect 42444 9441 42472 9472
rect 42904 9472 42993 9500
rect 39715 9404 40540 9432
rect 42429 9435 42487 9441
rect 39715 9401 39727 9404
rect 39669 9395 39727 9401
rect 42429 9401 42441 9435
rect 42475 9401 42487 9435
rect 42429 9395 42487 9401
rect 37829 9367 37887 9373
rect 37829 9364 37841 9367
rect 37516 9336 37841 9364
rect 37516 9324 37522 9336
rect 37829 9333 37841 9336
rect 37875 9333 37887 9367
rect 37829 9327 37887 9333
rect 38194 9324 38200 9376
rect 38252 9324 38258 9376
rect 38286 9324 38292 9376
rect 38344 9364 38350 9376
rect 39114 9364 39120 9376
rect 38344 9336 39120 9364
rect 38344 9324 38350 9336
rect 39114 9324 39120 9336
rect 39172 9324 39178 9376
rect 42334 9324 42340 9376
rect 42392 9364 42398 9376
rect 42904 9364 42932 9472
rect 42981 9469 42993 9472
rect 43027 9469 43039 9503
rect 43272 9500 43300 9540
rect 43346 9528 43352 9580
rect 43404 9568 43410 9580
rect 43993 9571 44051 9577
rect 43993 9568 44005 9571
rect 43404 9540 44005 9568
rect 43404 9528 43410 9540
rect 43993 9537 44005 9540
rect 44039 9537 44051 9571
rect 44100 9568 44128 9608
rect 44174 9596 44180 9648
rect 44232 9636 44238 9648
rect 44358 9636 44364 9648
rect 44232 9608 44364 9636
rect 44232 9596 44238 9608
rect 44358 9596 44364 9608
rect 44416 9596 44422 9648
rect 44726 9596 44732 9648
rect 44784 9636 44790 9648
rect 45373 9639 45431 9645
rect 45373 9636 45385 9639
rect 44784 9608 45385 9636
rect 44784 9596 44790 9608
rect 45373 9605 45385 9608
rect 45419 9605 45431 9639
rect 45373 9599 45431 9605
rect 46768 9580 46796 9676
rect 48774 9664 48780 9676
rect 48832 9704 48838 9716
rect 49050 9704 49056 9716
rect 48832 9676 49056 9704
rect 48832 9664 48838 9676
rect 49050 9664 49056 9676
rect 49108 9664 49114 9716
rect 49970 9664 49976 9716
rect 50028 9704 50034 9716
rect 50617 9707 50675 9713
rect 50617 9704 50629 9707
rect 50028 9676 50629 9704
rect 50028 9664 50034 9676
rect 50617 9673 50629 9676
rect 50663 9673 50675 9707
rect 50617 9667 50675 9673
rect 51810 9664 51816 9716
rect 51868 9664 51874 9716
rect 53190 9664 53196 9716
rect 53248 9704 53254 9716
rect 53285 9707 53343 9713
rect 53285 9704 53297 9707
rect 53248 9676 53297 9704
rect 53248 9664 53254 9676
rect 53285 9673 53297 9676
rect 53331 9673 53343 9707
rect 53285 9667 53343 9673
rect 47486 9596 47492 9648
rect 47544 9636 47550 9648
rect 47765 9639 47823 9645
rect 47765 9636 47777 9639
rect 47544 9608 47777 9636
rect 47544 9596 47550 9608
rect 47765 9605 47777 9608
rect 47811 9605 47823 9639
rect 56226 9636 56232 9648
rect 47765 9599 47823 9605
rect 55600 9608 56232 9636
rect 44818 9568 44824 9580
rect 44100 9540 44824 9568
rect 43993 9531 44051 9537
rect 44818 9528 44824 9540
rect 44876 9528 44882 9580
rect 46750 9528 46756 9580
rect 46808 9528 46814 9580
rect 48406 9528 48412 9580
rect 48464 9528 48470 9580
rect 51166 9528 51172 9580
rect 51224 9528 51230 9580
rect 53834 9528 53840 9580
rect 53892 9528 53898 9580
rect 54018 9528 54024 9580
rect 54076 9528 54082 9580
rect 54570 9528 54576 9580
rect 54628 9528 54634 9580
rect 44174 9500 44180 9512
rect 43272 9472 44180 9500
rect 42981 9463 43039 9469
rect 44174 9460 44180 9472
rect 44232 9460 44238 9512
rect 45002 9460 45008 9512
rect 45060 9500 45066 9512
rect 45557 9503 45615 9509
rect 45557 9500 45569 9503
rect 45060 9472 45569 9500
rect 45060 9460 45066 9472
rect 45557 9469 45569 9472
rect 45603 9469 45615 9503
rect 45557 9463 45615 9469
rect 46934 9460 46940 9512
rect 46992 9460 46998 9512
rect 55600 9509 55628 9608
rect 56226 9596 56232 9608
rect 56284 9636 56290 9648
rect 56686 9636 56692 9648
rect 56284 9608 56692 9636
rect 56284 9596 56290 9608
rect 56686 9596 56692 9608
rect 56744 9596 56750 9648
rect 56873 9639 56931 9645
rect 56873 9605 56885 9639
rect 56919 9636 56931 9639
rect 57790 9636 57796 9648
rect 56919 9608 57796 9636
rect 56919 9605 56931 9608
rect 56873 9599 56931 9605
rect 57790 9596 57796 9608
rect 57848 9596 57854 9648
rect 58250 9596 58256 9648
rect 58308 9596 58314 9648
rect 57514 9568 57520 9580
rect 56704 9540 57520 9568
rect 55585 9503 55643 9509
rect 55585 9500 55597 9503
rect 51184 9472 55597 9500
rect 51184 9444 51212 9472
rect 55585 9469 55597 9472
rect 55631 9469 55643 9503
rect 55585 9463 55643 9469
rect 55858 9460 55864 9512
rect 55916 9460 55922 9512
rect 47762 9392 47768 9444
rect 47820 9432 47826 9444
rect 47820 9404 51074 9432
rect 47820 9392 47826 9404
rect 42392 9336 42932 9364
rect 45005 9367 45063 9373
rect 42392 9324 42398 9336
rect 45005 9333 45017 9367
rect 45051 9364 45063 9367
rect 45094 9364 45100 9376
rect 45051 9336 45100 9364
rect 45051 9333 45063 9336
rect 45005 9327 45063 9333
rect 45094 9324 45100 9336
rect 45152 9324 45158 9376
rect 45830 9324 45836 9376
rect 45888 9364 45894 9376
rect 46017 9367 46075 9373
rect 46017 9364 46029 9367
rect 45888 9336 46029 9364
rect 45888 9324 45894 9336
rect 46017 9333 46029 9336
rect 46063 9333 46075 9367
rect 46017 9327 46075 9333
rect 46198 9324 46204 9376
rect 46256 9364 46262 9376
rect 46385 9367 46443 9373
rect 46385 9364 46397 9367
rect 46256 9336 46397 9364
rect 46256 9324 46262 9336
rect 46385 9333 46397 9336
rect 46431 9333 46443 9367
rect 46385 9327 46443 9333
rect 47118 9324 47124 9376
rect 47176 9364 47182 9376
rect 47305 9367 47363 9373
rect 47305 9364 47317 9367
rect 47176 9336 47317 9364
rect 47176 9324 47182 9336
rect 47305 9333 47317 9336
rect 47351 9333 47363 9367
rect 47305 9327 47363 9333
rect 48682 9324 48688 9376
rect 48740 9324 48746 9376
rect 49786 9324 49792 9376
rect 49844 9364 49850 9376
rect 49973 9367 50031 9373
rect 49973 9364 49985 9367
rect 49844 9336 49985 9364
rect 49844 9324 49850 9336
rect 49973 9333 49985 9336
rect 50019 9333 50031 9367
rect 51046 9364 51074 9404
rect 51166 9392 51172 9444
rect 51224 9392 51230 9444
rect 52270 9392 52276 9444
rect 52328 9432 52334 9444
rect 56704 9432 56732 9540
rect 57514 9528 57520 9540
rect 57572 9568 57578 9580
rect 58069 9571 58127 9577
rect 58069 9568 58081 9571
rect 57572 9540 58081 9568
rect 57572 9528 57578 9540
rect 58069 9537 58081 9540
rect 58115 9537 58127 9571
rect 58069 9531 58127 9537
rect 58434 9528 58440 9580
rect 58492 9528 58498 9580
rect 56778 9460 56784 9512
rect 56836 9460 56842 9512
rect 56962 9460 56968 9512
rect 57020 9460 57026 9512
rect 57054 9460 57060 9512
rect 57112 9460 57118 9512
rect 52328 9404 56732 9432
rect 56796 9432 56824 9460
rect 57072 9432 57100 9460
rect 56796 9404 57100 9432
rect 52328 9392 52334 9404
rect 53006 9364 53012 9376
rect 51046 9336 53012 9364
rect 49973 9327 50031 9333
rect 53006 9324 53012 9336
rect 53064 9324 53070 9376
rect 53466 9324 53472 9376
rect 53524 9364 53530 9376
rect 55125 9367 55183 9373
rect 55125 9364 55137 9367
rect 53524 9336 55137 9364
rect 53524 9324 53530 9336
rect 55125 9333 55137 9336
rect 55171 9333 55183 9367
rect 55125 9327 55183 9333
rect 56318 9324 56324 9376
rect 56376 9364 56382 9376
rect 56413 9367 56471 9373
rect 56413 9364 56425 9367
rect 56376 9336 56425 9364
rect 56376 9324 56382 9336
rect 56413 9333 56425 9336
rect 56459 9333 56471 9367
rect 56413 9327 56471 9333
rect 56505 9367 56563 9373
rect 56505 9333 56517 9367
rect 56551 9364 56563 9367
rect 57146 9364 57152 9376
rect 56551 9336 57152 9364
rect 56551 9333 56563 9336
rect 56505 9327 56563 9333
rect 57146 9324 57152 9336
rect 57204 9324 57210 9376
rect 1104 9274 58880 9296
rect 1104 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 22616 9274
rect 22668 9222 22680 9274
rect 22732 9222 22744 9274
rect 22796 9222 22808 9274
rect 22860 9222 22872 9274
rect 22924 9222 37060 9274
rect 37112 9222 37124 9274
rect 37176 9222 37188 9274
rect 37240 9222 37252 9274
rect 37304 9222 37316 9274
rect 37368 9222 51504 9274
rect 51556 9222 51568 9274
rect 51620 9222 51632 9274
rect 51684 9222 51696 9274
rect 51748 9222 51760 9274
rect 51812 9222 58880 9274
rect 1104 9200 58880 9222
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4801 9163 4859 9169
rect 4801 9160 4813 9163
rect 4396 9132 4813 9160
rect 4396 9120 4402 9132
rect 4801 9129 4813 9132
rect 4847 9129 4859 9163
rect 4801 9123 4859 9129
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5534 9120 5540 9172
rect 5592 9120 5598 9172
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8662 9160 8668 9172
rect 8435 9132 8668 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8662 9120 8668 9132
rect 8720 9160 8726 9172
rect 9122 9160 9128 9172
rect 8720 9132 9128 9160
rect 8720 9120 8726 9132
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 12342 9160 12348 9172
rect 9180 9132 12348 9160
rect 9180 9120 9186 9132
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 14734 9160 14740 9172
rect 13403 9132 14740 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 14884 9132 15884 9160
rect 14884 9120 14890 9132
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9061 3387 9095
rect 3329 9055 3387 9061
rect 4893 9095 4951 9101
rect 4893 9061 4905 9095
rect 4939 9092 4951 9095
rect 5000 9092 5028 9120
rect 4939 9064 7512 9092
rect 4939 9061 4951 9064
rect 4893 9055 4951 9061
rect 3344 9024 3372 9055
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 3344 8996 4353 9024
rect 4341 8993 4353 8996
rect 4387 9024 4399 9027
rect 6270 9024 6276 9036
rect 4387 8996 6276 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 7484 9033 7512 9064
rect 13814 9052 13820 9104
rect 13872 9052 13878 9104
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 7742 9024 7748 9036
rect 7515 8996 7748 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7742 8984 7748 8996
rect 7800 9024 7806 9036
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 7800 8996 9045 9024
rect 7800 8984 7806 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 14752 9024 14780 9120
rect 15519 9027 15577 9033
rect 15519 9024 15531 9027
rect 14752 8996 15531 9024
rect 9033 8987 9091 8993
rect 15519 8993 15531 8996
rect 15565 8993 15577 9027
rect 15519 8987 15577 8993
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 15856 9024 15884 9132
rect 15930 9120 15936 9172
rect 15988 9120 15994 9172
rect 18785 9163 18843 9169
rect 18785 9129 18797 9163
rect 18831 9160 18843 9163
rect 19610 9160 19616 9172
rect 18831 9132 19616 9160
rect 18831 9129 18843 9132
rect 18785 9123 18843 9129
rect 15948 9033 15976 9120
rect 15703 8996 15884 9024
rect 15933 9027 15991 9033
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15933 8993 15945 9027
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 9024 18475 9027
rect 18800 9024 18828 9123
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 22005 9163 22063 9169
rect 22005 9129 22017 9163
rect 22051 9160 22063 9163
rect 22094 9160 22100 9172
rect 22051 9132 22100 9160
rect 22051 9129 22063 9132
rect 22005 9123 22063 9129
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22756 9132 23704 9160
rect 21729 9095 21787 9101
rect 21729 9061 21741 9095
rect 21775 9092 21787 9095
rect 22756 9092 22784 9132
rect 21775 9064 22784 9092
rect 23676 9092 23704 9132
rect 23750 9120 23756 9172
rect 23808 9160 23814 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 23808 9132 24409 9160
rect 23808 9120 23814 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 24397 9123 24455 9129
rect 28813 9163 28871 9169
rect 28813 9129 28825 9163
rect 28859 9160 28871 9163
rect 30834 9160 30840 9172
rect 28859 9132 30840 9160
rect 28859 9129 28871 9132
rect 28813 9123 28871 9129
rect 30834 9120 30840 9132
rect 30892 9120 30898 9172
rect 30926 9120 30932 9172
rect 30984 9160 30990 9172
rect 31386 9160 31392 9172
rect 30984 9132 31392 9160
rect 30984 9120 30990 9132
rect 31386 9120 31392 9132
rect 31444 9160 31450 9172
rect 36446 9160 36452 9172
rect 31444 9132 36452 9160
rect 31444 9120 31450 9132
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 37553 9163 37611 9169
rect 37553 9129 37565 9163
rect 37599 9160 37611 9163
rect 37642 9160 37648 9172
rect 37599 9132 37648 9160
rect 37599 9129 37611 9132
rect 37553 9123 37611 9129
rect 37642 9120 37648 9132
rect 37700 9160 37706 9172
rect 37700 9132 39068 9160
rect 37700 9120 37706 9132
rect 23934 9092 23940 9104
rect 23676 9064 23940 9092
rect 21775 9061 21787 9064
rect 21729 9055 21787 9061
rect 18463 8996 18828 9024
rect 22649 9027 22707 9033
rect 18463 8993 18475 8996
rect 18417 8987 18475 8993
rect 22649 8993 22661 9027
rect 22695 9024 22707 9027
rect 22756 9024 22784 9064
rect 23934 9052 23940 9064
rect 23992 9052 23998 9104
rect 24121 9095 24179 9101
rect 24121 9061 24133 9095
rect 24167 9092 24179 9095
rect 24670 9092 24676 9104
rect 24167 9064 24676 9092
rect 24167 9061 24179 9064
rect 24121 9055 24179 9061
rect 24670 9052 24676 9064
rect 24728 9092 24734 9104
rect 24728 9064 24992 9092
rect 24728 9052 24734 9064
rect 24964 9033 24992 9064
rect 28994 9052 29000 9104
rect 29052 9092 29058 9104
rect 29273 9095 29331 9101
rect 29273 9092 29285 9095
rect 29052 9064 29285 9092
rect 29052 9052 29058 9064
rect 29273 9061 29285 9064
rect 29319 9061 29331 9095
rect 29273 9055 29331 9061
rect 31128 9064 32628 9092
rect 22695 8996 22784 9024
rect 24949 9027 25007 9033
rect 22695 8993 22707 8996
rect 22649 8987 22707 8993
rect 24949 8993 24961 9027
rect 24995 8993 25007 9027
rect 25682 9024 25688 9036
rect 24949 8987 25007 8993
rect 25056 8996 25688 9024
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 3326 8956 3332 8968
rect 1995 8928 3332 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5534 8956 5540 8968
rect 5307 8928 5540 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 2216 8891 2274 8897
rect 2216 8857 2228 8891
rect 2262 8888 2274 8891
rect 2406 8888 2412 8900
rect 2262 8860 2412 8888
rect 2262 8857 2274 8860
rect 2216 8851 2274 8857
rect 2406 8848 2412 8860
rect 2464 8848 2470 8900
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 8846 8888 8852 8900
rect 5408 8860 8852 8888
rect 5408 8848 5414 8860
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 9125 8891 9183 8897
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9214 8888 9220 8900
rect 9171 8860 9220 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 9214 8848 9220 8860
rect 9272 8848 9278 8900
rect 9508 8832 9536 8919
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9824 8928 9873 8956
rect 9824 8916 9830 8928
rect 9861 8925 9873 8928
rect 9907 8956 9919 8959
rect 11054 8956 11060 8968
rect 9907 8928 11060 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11882 8956 11888 8968
rect 11655 8928 11888 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 11882 8916 11888 8928
rect 11940 8956 11946 8968
rect 12250 8965 12256 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11940 8928 11989 8956
rect 11940 8916 11946 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 12244 8956 12256 8965
rect 12211 8928 12256 8956
rect 11977 8919 12035 8925
rect 12244 8919 12256 8928
rect 9582 8848 9588 8900
rect 9640 8848 9646 8900
rect 11992 8888 12020 8919
rect 12250 8916 12256 8919
rect 12308 8916 12314 8968
rect 15378 8916 15384 8968
rect 15436 8916 15442 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 12342 8888 12348 8900
rect 11992 8860 12348 8888
rect 12342 8848 12348 8860
rect 12400 8888 12406 8900
rect 16408 8888 16436 8919
rect 16574 8916 16580 8968
rect 16632 8916 16638 8968
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 20349 8959 20407 8965
rect 16724 8928 18828 8956
rect 16724 8916 16730 8928
rect 12400 8860 13492 8888
rect 16408 8860 17080 8888
rect 12400 8848 12406 8860
rect 13464 8832 13492 8860
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 6144 8792 6929 8820
rect 6144 8780 6150 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 6917 8783 6975 8789
rect 9490 8780 9496 8832
rect 9548 8780 9554 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 14642 8820 14648 8832
rect 14332 8792 14648 8820
rect 14332 8780 14338 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 16942 8820 16948 8832
rect 14783 8792 16948 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17052 8829 17080 8860
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18150 8891 18208 8897
rect 18150 8888 18162 8891
rect 18012 8860 18162 8888
rect 18012 8848 18018 8860
rect 18150 8857 18162 8860
rect 18196 8857 18208 8891
rect 18150 8851 18208 8857
rect 17037 8823 17095 8829
rect 17037 8789 17049 8823
rect 17083 8820 17095 8823
rect 18690 8820 18696 8832
rect 17083 8792 18696 8820
rect 17083 8789 17095 8792
rect 17037 8783 17095 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18800 8820 18828 8928
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20438 8956 20444 8968
rect 20395 8928 20444 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 24026 8956 24032 8968
rect 22787 8928 24032 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 25056 8956 25084 8996
rect 25682 8984 25688 8996
rect 25740 8984 25746 9036
rect 25866 8984 25872 9036
rect 25924 8984 25930 9036
rect 26602 8984 26608 9036
rect 26660 8984 26666 9036
rect 27706 8965 27712 8968
rect 24872 8928 25084 8956
rect 27433 8959 27491 8965
rect 24872 8900 24900 8928
rect 27433 8925 27445 8959
rect 27479 8925 27491 8959
rect 27700 8956 27712 8965
rect 27667 8928 27712 8956
rect 27433 8919 27491 8925
rect 27700 8919 27712 8928
rect 20616 8891 20674 8897
rect 20616 8857 20628 8891
rect 20662 8888 20674 8891
rect 21818 8888 21824 8900
rect 20662 8860 21824 8888
rect 20662 8857 20674 8860
rect 20616 8851 20674 8857
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 23008 8891 23066 8897
rect 23008 8857 23020 8891
rect 23054 8888 23066 8891
rect 23198 8888 23204 8900
rect 23054 8860 23204 8888
rect 23054 8857 23066 8860
rect 23008 8851 23066 8857
rect 23198 8848 23204 8860
rect 23256 8848 23262 8900
rect 24854 8848 24860 8900
rect 24912 8848 24918 8900
rect 25593 8891 25651 8897
rect 25148 8860 25544 8888
rect 25148 8820 25176 8860
rect 18800 8792 25176 8820
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 25516 8820 25544 8860
rect 25593 8857 25605 8891
rect 25639 8888 25651 8891
rect 26053 8891 26111 8897
rect 26053 8888 26065 8891
rect 25639 8860 26065 8888
rect 25639 8857 25651 8860
rect 25593 8851 25651 8857
rect 26053 8857 26065 8860
rect 26099 8857 26111 8891
rect 27448 8888 27476 8919
rect 27706 8916 27712 8919
rect 27764 8916 27770 8968
rect 29288 8956 29316 9055
rect 31128 9033 31156 9064
rect 31113 9027 31171 9033
rect 31113 8993 31125 9027
rect 31159 8993 31171 9027
rect 31113 8987 31171 8993
rect 31202 8984 31208 9036
rect 31260 8984 31266 9036
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29288 8928 29561 8956
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 31754 8916 31760 8968
rect 31812 8916 31818 8968
rect 27614 8888 27620 8900
rect 27448 8860 27620 8888
rect 26053 8851 26111 8857
rect 27614 8848 27620 8860
rect 27672 8848 27678 8900
rect 30190 8848 30196 8900
rect 30248 8888 30254 8900
rect 32600 8897 32628 9064
rect 39040 9033 39068 9132
rect 42794 9120 42800 9172
rect 42852 9120 42858 9172
rect 43346 9120 43352 9172
rect 43404 9160 43410 9172
rect 43717 9163 43775 9169
rect 43717 9160 43729 9163
rect 43404 9132 43729 9160
rect 43404 9120 43410 9132
rect 43717 9129 43729 9132
rect 43763 9129 43775 9163
rect 43717 9123 43775 9129
rect 44358 9120 44364 9172
rect 44416 9120 44422 9172
rect 44545 9163 44603 9169
rect 44545 9129 44557 9163
rect 44591 9160 44603 9163
rect 45370 9160 45376 9172
rect 44591 9132 45376 9160
rect 44591 9129 44603 9132
rect 44545 9123 44603 9129
rect 45370 9120 45376 9132
rect 45428 9120 45434 9172
rect 46569 9163 46627 9169
rect 46569 9129 46581 9163
rect 46615 9160 46627 9163
rect 46934 9160 46940 9172
rect 46615 9132 46940 9160
rect 46615 9129 46627 9132
rect 46569 9123 46627 9129
rect 46934 9120 46940 9132
rect 46992 9120 46998 9172
rect 51074 9120 51080 9172
rect 51132 9160 51138 9172
rect 51445 9163 51503 9169
rect 51445 9160 51457 9163
rect 51132 9132 51457 9160
rect 51132 9120 51138 9132
rect 51445 9129 51457 9132
rect 51491 9129 51503 9163
rect 53837 9163 53895 9169
rect 51445 9123 51503 9129
rect 52932 9132 53788 9160
rect 39114 9052 39120 9104
rect 39172 9092 39178 9104
rect 43364 9092 43392 9120
rect 39172 9064 43392 9092
rect 44376 9092 44404 9120
rect 45557 9095 45615 9101
rect 45557 9092 45569 9095
rect 44376 9064 45569 9092
rect 39172 9052 39178 9064
rect 45557 9061 45569 9064
rect 45603 9092 45615 9095
rect 46658 9092 46664 9104
rect 45603 9064 46664 9092
rect 45603 9061 45615 9064
rect 45557 9055 45615 9061
rect 46658 9052 46664 9064
rect 46716 9092 46722 9104
rect 49602 9092 49608 9104
rect 46716 9064 49608 9092
rect 46716 9052 46722 9064
rect 49602 9052 49608 9064
rect 49660 9092 49666 9104
rect 49697 9095 49755 9101
rect 49697 9092 49709 9095
rect 49660 9064 49709 9092
rect 49660 9052 49666 9064
rect 49697 9061 49709 9064
rect 49743 9061 49755 9095
rect 49697 9055 49755 9061
rect 51258 9052 51264 9104
rect 51316 9092 51322 9104
rect 52932 9092 52960 9132
rect 51316 9064 52960 9092
rect 53009 9095 53067 9101
rect 51316 9052 51322 9064
rect 53009 9061 53021 9095
rect 53055 9061 53067 9095
rect 53009 9055 53067 9061
rect 39025 9027 39083 9033
rect 39025 8993 39037 9027
rect 39071 8993 39083 9027
rect 39025 8987 39083 8993
rect 43438 8984 43444 9036
rect 43496 8984 43502 9036
rect 44818 8984 44824 9036
rect 44876 9024 44882 9036
rect 45189 9027 45247 9033
rect 45189 9024 45201 9027
rect 44876 8996 45201 9024
rect 44876 8984 44882 8996
rect 45189 8993 45201 8996
rect 45235 9024 45247 9027
rect 46750 9024 46756 9036
rect 45235 8996 46756 9024
rect 45235 8993 45247 8996
rect 45189 8987 45247 8993
rect 46750 8984 46756 8996
rect 46808 8984 46814 9036
rect 47118 8984 47124 9036
rect 47176 8984 47182 9036
rect 48682 9024 48688 9036
rect 47964 8996 48688 9024
rect 32858 8916 32864 8968
rect 32916 8916 32922 8968
rect 33410 8916 33416 8968
rect 33468 8916 33474 8968
rect 34701 8959 34759 8965
rect 34701 8956 34713 8959
rect 34440 8928 34713 8956
rect 30377 8891 30435 8897
rect 30377 8888 30389 8891
rect 30248 8860 30389 8888
rect 30248 8848 30254 8860
rect 30377 8857 30389 8860
rect 30423 8857 30435 8891
rect 30377 8851 30435 8857
rect 32585 8891 32643 8897
rect 32585 8857 32597 8891
rect 32631 8888 32643 8891
rect 32631 8860 33824 8888
rect 32631 8857 32643 8860
rect 32585 8851 32643 8857
rect 33796 8832 33824 8860
rect 30742 8820 30748 8832
rect 25516 8792 30748 8820
rect 30742 8780 30748 8792
rect 30800 8780 30806 8832
rect 31294 8780 31300 8832
rect 31352 8780 31358 8832
rect 31662 8780 31668 8832
rect 31720 8780 31726 8832
rect 33778 8780 33784 8832
rect 33836 8780 33842 8832
rect 34238 8780 34244 8832
rect 34296 8820 34302 8832
rect 34440 8829 34468 8928
rect 34701 8925 34713 8928
rect 34747 8925 34759 8959
rect 34701 8919 34759 8925
rect 36722 8916 36728 8968
rect 36780 8916 36786 8968
rect 38930 8916 38936 8968
rect 38988 8916 38994 8968
rect 40402 8916 40408 8968
rect 40460 8916 40466 8968
rect 47964 8956 47992 8996
rect 48682 8984 48688 8996
rect 48740 9024 48746 9036
rect 49237 9027 49295 9033
rect 49237 9024 49249 9027
rect 48740 8996 49249 9024
rect 48740 8984 48746 8996
rect 49237 8993 49249 8996
rect 49283 9024 49295 9027
rect 49283 8996 49464 9024
rect 49283 8993 49295 8996
rect 49237 8987 49295 8993
rect 41386 8928 47992 8956
rect 34968 8891 35026 8897
rect 34968 8857 34980 8891
rect 35014 8888 35026 8891
rect 36173 8891 36231 8897
rect 36173 8888 36185 8891
rect 35014 8860 36185 8888
rect 35014 8857 35026 8860
rect 34968 8851 35026 8857
rect 36173 8857 36185 8860
rect 36219 8857 36231 8891
rect 36173 8851 36231 8857
rect 38688 8891 38746 8897
rect 38688 8857 38700 8891
rect 38734 8888 38746 8891
rect 39853 8891 39911 8897
rect 39853 8888 39865 8891
rect 38734 8860 39865 8888
rect 38734 8857 38746 8860
rect 38688 8851 38746 8857
rect 39853 8857 39865 8860
rect 39899 8857 39911 8891
rect 39853 8851 39911 8857
rect 40310 8848 40316 8900
rect 40368 8888 40374 8900
rect 41386 8888 41414 8928
rect 48038 8916 48044 8968
rect 48096 8956 48102 8968
rect 49326 8956 49332 8968
rect 48096 8928 49332 8956
rect 48096 8916 48102 8928
rect 49326 8916 49332 8928
rect 49384 8916 49390 8968
rect 49436 8956 49464 8996
rect 49786 8984 49792 9036
rect 49844 9024 49850 9036
rect 50249 9027 50307 9033
rect 50249 9024 50261 9027
rect 49844 8996 50261 9024
rect 49844 8984 49850 8996
rect 50249 8993 50261 8996
rect 50295 9024 50307 9027
rect 52270 9024 52276 9036
rect 50295 8996 52276 9024
rect 50295 8993 50307 8996
rect 50249 8987 50307 8993
rect 52270 8984 52276 8996
rect 52328 8984 52334 9036
rect 52365 9027 52423 9033
rect 52365 8993 52377 9027
rect 52411 9024 52423 9027
rect 53024 9024 53052 9055
rect 52411 8996 53052 9024
rect 53561 9027 53619 9033
rect 52411 8993 52423 8996
rect 52365 8987 52423 8993
rect 53561 8993 53573 9027
rect 53607 8993 53619 9027
rect 53760 9024 53788 9132
rect 53837 9129 53849 9163
rect 53883 9160 53895 9163
rect 53883 9132 53972 9160
rect 53883 9129 53895 9132
rect 53837 9123 53895 9129
rect 53944 9104 53972 9132
rect 55858 9120 55864 9172
rect 55916 9160 55922 9172
rect 56505 9163 56563 9169
rect 56505 9160 56517 9163
rect 55916 9132 56517 9160
rect 55916 9120 55922 9132
rect 56505 9129 56517 9132
rect 56551 9129 56563 9163
rect 56505 9123 56563 9129
rect 56686 9120 56692 9172
rect 56744 9160 56750 9172
rect 56744 9132 57100 9160
rect 56744 9120 56750 9132
rect 53926 9052 53932 9104
rect 53984 9052 53990 9104
rect 56321 9095 56379 9101
rect 56321 9092 56333 9095
rect 54128 9064 56333 9092
rect 54128 9024 54156 9064
rect 56321 9061 56333 9064
rect 56367 9092 56379 9095
rect 56778 9092 56784 9104
rect 56367 9064 56784 9092
rect 56367 9061 56379 9064
rect 56321 9055 56379 9061
rect 56778 9052 56784 9064
rect 56836 9052 56842 9104
rect 57072 9092 57100 9132
rect 58345 9095 58403 9101
rect 58345 9092 58357 9095
rect 57072 9064 58357 9092
rect 53760 8996 54156 9024
rect 53561 8987 53619 8993
rect 51074 8956 51080 8968
rect 49436 8928 51080 8956
rect 51074 8916 51080 8928
rect 51132 8916 51138 8968
rect 53006 8916 53012 8968
rect 53064 8956 53070 8968
rect 53576 8956 53604 8987
rect 54386 8984 54392 9036
rect 54444 9024 54450 9036
rect 57072 9033 57100 9064
rect 58345 9061 58357 9064
rect 58391 9061 58403 9095
rect 58345 9055 58403 9061
rect 54849 9027 54907 9033
rect 54849 9024 54861 9027
rect 54444 8996 54861 9024
rect 54444 8984 54450 8996
rect 54849 8993 54861 8996
rect 54895 8993 54907 9027
rect 54849 8987 54907 8993
rect 57057 9027 57115 9033
rect 57057 8993 57069 9027
rect 57103 8993 57115 9027
rect 57057 8987 57115 8993
rect 57238 8984 57244 9036
rect 57296 9024 57302 9036
rect 57514 9024 57520 9036
rect 57296 8996 57520 9024
rect 57296 8984 57302 8996
rect 57514 8984 57520 8996
rect 57572 8984 57578 9036
rect 53064 8928 53604 8956
rect 53064 8916 53070 8928
rect 54018 8916 54024 8968
rect 54076 8956 54082 8968
rect 54297 8959 54355 8965
rect 54297 8956 54309 8959
rect 54076 8928 54309 8956
rect 54076 8916 54082 8928
rect 54297 8925 54309 8928
rect 54343 8925 54355 8959
rect 54297 8919 54355 8925
rect 54662 8916 54668 8968
rect 54720 8956 54726 8968
rect 55861 8959 55919 8965
rect 55861 8956 55873 8959
rect 54720 8928 55873 8956
rect 54720 8916 54726 8928
rect 55861 8925 55873 8928
rect 55907 8925 55919 8959
rect 55861 8919 55919 8925
rect 40368 8860 41414 8888
rect 44453 8891 44511 8897
rect 40368 8848 40374 8860
rect 44453 8857 44465 8891
rect 44499 8888 44511 8891
rect 44726 8888 44732 8900
rect 44499 8860 44732 8888
rect 44499 8857 44511 8860
rect 44453 8851 44511 8857
rect 44726 8848 44732 8860
rect 44784 8848 44790 8900
rect 46937 8891 46995 8897
rect 46937 8857 46949 8891
rect 46983 8888 46995 8891
rect 48222 8888 48228 8900
rect 46983 8860 48228 8888
rect 46983 8857 46995 8860
rect 46937 8851 46995 8857
rect 48222 8848 48228 8860
rect 48280 8888 48286 8900
rect 49053 8891 49111 8897
rect 49053 8888 49065 8891
rect 48280 8860 49065 8888
rect 48280 8848 48286 8860
rect 49053 8857 49065 8860
rect 49099 8888 49111 8891
rect 50338 8888 50344 8900
rect 49099 8860 50344 8888
rect 49099 8857 49111 8860
rect 49053 8851 49111 8857
rect 50338 8848 50344 8860
rect 50396 8888 50402 8900
rect 50433 8891 50491 8897
rect 50433 8888 50445 8891
rect 50396 8860 50445 8888
rect 50396 8848 50402 8860
rect 50433 8857 50445 8860
rect 50479 8857 50491 8891
rect 50433 8851 50491 8857
rect 50525 8891 50583 8897
rect 50525 8857 50537 8891
rect 50571 8888 50583 8891
rect 51166 8888 51172 8900
rect 50571 8860 51172 8888
rect 50571 8857 50583 8860
rect 50525 8851 50583 8857
rect 51166 8848 51172 8860
rect 51224 8848 51230 8900
rect 51350 8848 51356 8900
rect 51408 8888 51414 8900
rect 51537 8891 51595 8897
rect 51537 8888 51549 8891
rect 51408 8860 51549 8888
rect 51408 8848 51414 8860
rect 51537 8857 51549 8860
rect 51583 8857 51595 8891
rect 51537 8851 51595 8857
rect 53377 8891 53435 8897
rect 53377 8857 53389 8891
rect 53423 8888 53435 8891
rect 55309 8891 55367 8897
rect 55309 8888 55321 8891
rect 53423 8860 55321 8888
rect 53423 8857 53435 8860
rect 53377 8851 53435 8857
rect 55309 8857 55321 8860
rect 55355 8857 55367 8891
rect 55309 8851 55367 8857
rect 56965 8891 57023 8897
rect 56965 8857 56977 8891
rect 57011 8888 57023 8891
rect 57790 8888 57796 8900
rect 57011 8860 57796 8888
rect 57011 8857 57023 8860
rect 56965 8851 57023 8857
rect 57790 8848 57796 8860
rect 57848 8848 57854 8900
rect 34425 8823 34483 8829
rect 34425 8820 34437 8823
rect 34296 8792 34437 8820
rect 34296 8780 34302 8792
rect 34425 8789 34437 8792
rect 34471 8789 34483 8823
rect 34425 8783 34483 8789
rect 36078 8780 36084 8832
rect 36136 8820 36142 8832
rect 36906 8820 36912 8832
rect 36136 8792 36912 8820
rect 36136 8780 36142 8792
rect 36906 8780 36912 8792
rect 36964 8780 36970 8832
rect 39666 8780 39672 8832
rect 39724 8780 39730 8832
rect 40494 8780 40500 8832
rect 40552 8820 40558 8832
rect 40773 8823 40831 8829
rect 40773 8820 40785 8823
rect 40552 8792 40785 8820
rect 40552 8780 40558 8792
rect 40773 8789 40785 8792
rect 40819 8820 40831 8823
rect 41141 8823 41199 8829
rect 41141 8820 41153 8823
rect 40819 8792 41153 8820
rect 40819 8789 40831 8792
rect 40773 8783 40831 8789
rect 41141 8789 41153 8792
rect 41187 8789 41199 8823
rect 41141 8783 41199 8789
rect 42334 8780 42340 8832
rect 42392 8780 42398 8832
rect 44269 8823 44327 8829
rect 44269 8789 44281 8823
rect 44315 8820 44327 8823
rect 45002 8820 45008 8832
rect 44315 8792 45008 8820
rect 44315 8789 44327 8792
rect 44269 8783 44327 8789
rect 45002 8780 45008 8792
rect 45060 8780 45066 8832
rect 45370 8780 45376 8832
rect 45428 8820 45434 8832
rect 45830 8820 45836 8832
rect 45428 8792 45836 8820
rect 45428 8780 45434 8792
rect 45830 8780 45836 8792
rect 45888 8820 45894 8832
rect 45925 8823 45983 8829
rect 45925 8820 45937 8823
rect 45888 8792 45937 8820
rect 45888 8780 45894 8792
rect 45925 8789 45937 8792
rect 45971 8820 45983 8823
rect 46293 8823 46351 8829
rect 46293 8820 46305 8823
rect 45971 8792 46305 8820
rect 45971 8789 45983 8792
rect 45925 8783 45983 8789
rect 46293 8789 46305 8792
rect 46339 8789 46351 8823
rect 46293 8783 46351 8789
rect 47029 8823 47087 8829
rect 47029 8789 47041 8823
rect 47075 8820 47087 8823
rect 47397 8823 47455 8829
rect 47397 8820 47409 8823
rect 47075 8792 47409 8820
rect 47075 8789 47087 8792
rect 47029 8783 47087 8789
rect 47397 8789 47409 8792
rect 47443 8789 47455 8823
rect 47397 8783 47455 8789
rect 47762 8780 47768 8832
rect 47820 8820 47826 8832
rect 48317 8823 48375 8829
rect 48317 8820 48329 8823
rect 47820 8792 48329 8820
rect 47820 8780 47826 8792
rect 48317 8789 48329 8792
rect 48363 8789 48375 8823
rect 48317 8783 48375 8789
rect 48682 8780 48688 8832
rect 48740 8780 48746 8832
rect 49142 8780 49148 8832
rect 49200 8780 49206 8832
rect 50890 8780 50896 8832
rect 50948 8780 50954 8832
rect 52914 8780 52920 8832
rect 52972 8780 52978 8832
rect 53469 8823 53527 8829
rect 53469 8789 53481 8823
rect 53515 8820 53527 8823
rect 53742 8820 53748 8832
rect 53515 8792 53748 8820
rect 53515 8789 53527 8792
rect 53469 8783 53527 8789
rect 53742 8780 53748 8792
rect 53800 8820 53806 8832
rect 54205 8823 54263 8829
rect 54205 8820 54217 8823
rect 53800 8792 54217 8820
rect 53800 8780 53806 8792
rect 54205 8789 54217 8792
rect 54251 8789 54263 8823
rect 54205 8783 54263 8789
rect 56870 8780 56876 8832
rect 56928 8820 56934 8832
rect 57609 8823 57667 8829
rect 57609 8820 57621 8823
rect 56928 8792 57621 8820
rect 56928 8780 56934 8792
rect 57609 8789 57621 8792
rect 57655 8789 57667 8823
rect 57609 8783 57667 8789
rect 57701 8823 57759 8829
rect 57701 8789 57713 8823
rect 57747 8820 57759 8823
rect 57882 8820 57888 8832
rect 57747 8792 57888 8820
rect 57747 8789 57759 8792
rect 57701 8783 57759 8789
rect 57882 8780 57888 8792
rect 57940 8780 57946 8832
rect 58066 8780 58072 8832
rect 58124 8780 58130 8832
rect 1104 8730 59040 8752
rect 1104 8678 15394 8730
rect 15446 8678 15458 8730
rect 15510 8678 15522 8730
rect 15574 8678 15586 8730
rect 15638 8678 15650 8730
rect 15702 8678 29838 8730
rect 29890 8678 29902 8730
rect 29954 8678 29966 8730
rect 30018 8678 30030 8730
rect 30082 8678 30094 8730
rect 30146 8678 44282 8730
rect 44334 8678 44346 8730
rect 44398 8678 44410 8730
rect 44462 8678 44474 8730
rect 44526 8678 44538 8730
rect 44590 8678 58726 8730
rect 58778 8678 58790 8730
rect 58842 8678 58854 8730
rect 58906 8678 58918 8730
rect 58970 8678 58982 8730
rect 59034 8678 59040 8730
rect 1104 8656 59040 8678
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 3878 8616 3884 8628
rect 2746 8588 3884 8616
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 2746 8548 2774 8588
rect 3878 8576 3884 8588
rect 3936 8616 3942 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3936 8588 3985 8616
rect 3936 8576 3942 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 5721 8619 5779 8625
rect 3973 8579 4031 8585
rect 4264 8588 5672 8616
rect 2271 8520 2774 8548
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 4157 8551 4215 8557
rect 4157 8548 4169 8551
rect 3844 8520 4169 8548
rect 3844 8508 3850 8520
rect 4157 8517 4169 8520
rect 4203 8517 4215 8551
rect 4157 8511 4215 8517
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 2363 8452 3249 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 2056 8412 2084 8443
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 4264 8480 4292 8588
rect 5534 8508 5540 8560
rect 5592 8508 5598 8560
rect 3384 8452 4292 8480
rect 3384 8440 3390 8452
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 4396 8452 5580 8480
rect 4396 8440 4402 8452
rect 2222 8412 2228 8424
rect 2056 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2746 8384 2973 8412
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2746 8344 2774 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3878 8372 3884 8424
rect 3936 8372 3942 8424
rect 2087 8316 2774 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 5169 8347 5227 8353
rect 5169 8344 5181 8347
rect 4580 8316 5181 8344
rect 4580 8304 4586 8316
rect 5169 8313 5181 8316
rect 5215 8344 5227 8347
rect 5350 8344 5356 8356
rect 5215 8316 5356 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5552 8285 5580 8452
rect 5644 8412 5672 8588
rect 5721 8585 5733 8619
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 5736 8548 5764 8579
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 9582 8616 9588 8628
rect 8680 8588 9588 8616
rect 5736 8520 6224 8548
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6086 8480 6092 8492
rect 6043 8452 6092 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6196 8480 6224 8520
rect 6196 8452 6684 8480
rect 6656 8421 6684 8452
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5644 8384 6377 8412
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8381 6699 8415
rect 7760 8412 7788 8576
rect 8680 8492 8708 8588
rect 9582 8576 9588 8588
rect 9640 8616 9646 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9640 8588 9873 8616
rect 9640 8576 9646 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 12986 8616 12992 8628
rect 10091 8588 12992 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 16025 8619 16083 8625
rect 13311 8588 14872 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 14844 8560 14872 8588
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16574 8616 16580 8628
rect 16071 8588 16580 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 17770 8576 17776 8628
rect 17828 8576 17834 8628
rect 21818 8576 21824 8628
rect 21876 8576 21882 8628
rect 22462 8576 22468 8628
rect 22520 8576 22526 8628
rect 23198 8576 23204 8628
rect 23256 8576 23262 8628
rect 25222 8576 25228 8628
rect 25280 8576 25286 8628
rect 25869 8619 25927 8625
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 26050 8616 26056 8628
rect 25915 8588 26056 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 29917 8619 29975 8625
rect 29917 8585 29929 8619
rect 29963 8616 29975 8619
rect 31294 8616 31300 8628
rect 29963 8588 31300 8616
rect 29963 8585 29975 8588
rect 29917 8579 29975 8585
rect 31294 8576 31300 8588
rect 31352 8576 31358 8628
rect 32125 8619 32183 8625
rect 32125 8616 32137 8619
rect 31726 8588 32137 8616
rect 9490 8548 9496 8560
rect 8772 8520 9496 8548
rect 8772 8492 8800 8520
rect 9490 8508 9496 8520
rect 9548 8548 9554 8560
rect 9677 8551 9735 8557
rect 9677 8548 9689 8551
rect 9548 8520 9689 8548
rect 9548 8508 9554 8520
rect 9677 8517 9689 8520
rect 9723 8517 9735 8551
rect 9677 8511 9735 8517
rect 14826 8508 14832 8560
rect 14884 8508 14890 8560
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8662 8480 8668 8492
rect 8343 8452 8668 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 10134 8480 10140 8492
rect 9631 8452 10140 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 8956 8412 8984 8443
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 11882 8440 11888 8492
rect 11940 8489 11946 8492
rect 12158 8489 12164 8492
rect 11940 8480 11950 8489
rect 11940 8452 11985 8480
rect 11940 8443 11950 8452
rect 12152 8443 12164 8489
rect 11940 8440 11946 8443
rect 12158 8440 12164 8443
rect 12216 8440 12222 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 14918 8489 14924 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13504 8452 14657 8480
rect 13504 8440 13510 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14912 8443 14924 8489
rect 14918 8440 14924 8443
rect 14976 8440 14982 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 17727 8452 18153 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 21174 8480 21180 8492
rect 19076 8452 21180 8480
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 7760 8384 8984 8412
rect 6641 8375 6699 8381
rect 5537 8279 5595 8285
rect 5537 8245 5549 8279
rect 5583 8276 5595 8279
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5583 8248 5917 8276
rect 5583 8245 5595 8248
rect 5537 8239 5595 8245
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 6380 8276 6408 8375
rect 8570 8344 8576 8356
rect 7300 8316 8576 8344
rect 7300 8276 7328 8316
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 6380 8248 7328 8276
rect 8956 8276 8984 8384
rect 13004 8384 13737 8412
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 9456 8316 10425 8344
rect 9456 8304 9462 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11422 8344 11428 8356
rect 11379 8316 11428 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 13004 8288 13032 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 17865 8415 17923 8421
rect 17865 8412 17877 8415
rect 13725 8375 13783 8381
rect 17144 8384 17877 8412
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 13814 8344 13820 8356
rect 13596 8316 13820 8344
rect 13596 8304 13602 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 16850 8304 16856 8356
rect 16908 8344 16914 8356
rect 17144 8353 17172 8384
rect 17865 8381 17877 8384
rect 17911 8412 17923 8415
rect 19076 8412 19104 8452
rect 21174 8440 21180 8452
rect 21232 8480 21238 8492
rect 22480 8489 22508 8576
rect 22572 8520 25176 8548
rect 22465 8483 22523 8489
rect 21232 8452 21956 8480
rect 21232 8440 21238 8452
rect 17911 8384 19104 8412
rect 17911 8381 17923 8384
rect 17865 8375 17923 8381
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 19208 8384 19441 8412
rect 19208 8372 19214 8384
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 21928 8412 21956 8452
rect 22465 8449 22477 8483
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 22572 8412 22600 8520
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23753 8483 23811 8489
rect 23753 8480 23765 8483
rect 23624 8452 23765 8480
rect 23624 8440 23630 8452
rect 23753 8449 23765 8452
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 21928 8384 22600 8412
rect 22833 8415 22891 8421
rect 19429 8375 19487 8381
rect 22833 8381 22845 8415
rect 22879 8412 22891 8415
rect 23474 8412 23480 8424
rect 22879 8384 23480 8412
rect 22879 8381 22891 8384
rect 22833 8375 22891 8381
rect 23474 8372 23480 8384
rect 23532 8412 23538 8424
rect 23658 8412 23664 8424
rect 23532 8384 23664 8412
rect 23532 8372 23538 8384
rect 23658 8372 23664 8384
rect 23716 8372 23722 8424
rect 25148 8421 25176 8520
rect 25240 8489 25268 8576
rect 27709 8551 27767 8557
rect 27709 8517 27721 8551
rect 27755 8548 27767 8551
rect 28046 8551 28104 8557
rect 28046 8548 28058 8551
rect 27755 8520 28058 8548
rect 27755 8517 27767 8520
rect 27709 8511 27767 8517
rect 28046 8517 28058 8520
rect 28092 8517 28104 8551
rect 28046 8511 28104 8517
rect 25225 8483 25283 8489
rect 25225 8449 25237 8483
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8480 27215 8483
rect 28442 8480 28448 8492
rect 27203 8452 28448 8480
rect 27203 8449 27215 8452
rect 27157 8443 27215 8449
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 30558 8440 30564 8492
rect 30616 8440 30622 8492
rect 30834 8440 30840 8492
rect 30892 8440 30898 8492
rect 31573 8483 31631 8489
rect 31573 8449 31585 8483
rect 31619 8480 31631 8483
rect 31726 8480 31754 8588
rect 32125 8585 32137 8588
rect 32171 8616 32183 8619
rect 33410 8616 33416 8628
rect 32171 8588 33416 8616
rect 32171 8585 32183 8588
rect 32125 8579 32183 8585
rect 33410 8576 33416 8588
rect 33468 8576 33474 8628
rect 35894 8576 35900 8628
rect 35952 8616 35958 8628
rect 35989 8619 36047 8625
rect 35989 8616 36001 8619
rect 35952 8588 36001 8616
rect 35952 8576 35958 8588
rect 35989 8585 36001 8588
rect 36035 8585 36047 8619
rect 35989 8579 36047 8585
rect 36449 8619 36507 8625
rect 36449 8585 36461 8619
rect 36495 8616 36507 8619
rect 36722 8616 36728 8628
rect 36495 8588 36728 8616
rect 36495 8585 36507 8588
rect 36449 8579 36507 8585
rect 36722 8576 36728 8588
rect 36780 8576 36786 8628
rect 38930 8576 38936 8628
rect 38988 8576 38994 8628
rect 39117 8619 39175 8625
rect 39117 8585 39129 8619
rect 39163 8616 39175 8619
rect 39666 8616 39672 8628
rect 39163 8588 39672 8616
rect 39163 8585 39175 8588
rect 39117 8579 39175 8585
rect 39666 8576 39672 8588
rect 39724 8576 39730 8628
rect 39758 8576 39764 8628
rect 39816 8576 39822 8628
rect 44634 8576 44640 8628
rect 44692 8616 44698 8628
rect 44821 8619 44879 8625
rect 44821 8616 44833 8619
rect 44692 8588 44833 8616
rect 44692 8576 44698 8588
rect 44821 8585 44833 8588
rect 44867 8585 44879 8619
rect 44821 8579 44879 8585
rect 46198 8576 46204 8628
rect 46256 8576 46262 8628
rect 47213 8619 47271 8625
rect 47213 8585 47225 8619
rect 47259 8616 47271 8619
rect 48038 8616 48044 8628
rect 47259 8588 48044 8616
rect 47259 8585 47271 8588
rect 47213 8579 47271 8585
rect 48038 8576 48044 8588
rect 48096 8576 48102 8628
rect 48222 8576 48228 8628
rect 48280 8576 48286 8628
rect 48409 8619 48467 8625
rect 48409 8585 48421 8619
rect 48455 8616 48467 8619
rect 50617 8619 50675 8625
rect 50617 8616 50629 8619
rect 48455 8588 50629 8616
rect 48455 8585 48467 8588
rect 48409 8579 48467 8585
rect 50617 8585 50629 8588
rect 50663 8585 50675 8619
rect 50617 8579 50675 8585
rect 50890 8576 50896 8628
rect 50948 8616 50954 8628
rect 50948 8588 51074 8616
rect 50948 8576 50954 8588
rect 38948 8548 38976 8576
rect 40494 8548 40500 8560
rect 31619 8452 31754 8480
rect 32416 8520 33548 8548
rect 31619 8449 31631 8452
rect 31573 8443 31631 8449
rect 32416 8424 32444 8520
rect 33249 8483 33307 8489
rect 33249 8449 33261 8483
rect 33295 8480 33307 8483
rect 33410 8480 33416 8492
rect 33295 8452 33416 8480
rect 33295 8449 33307 8452
rect 33249 8443 33307 8449
rect 33410 8440 33416 8452
rect 33468 8440 33474 8492
rect 33520 8489 33548 8520
rect 36096 8520 38608 8548
rect 33505 8483 33563 8489
rect 33505 8449 33517 8483
rect 33551 8480 33563 8483
rect 34238 8480 34244 8492
rect 33551 8452 34244 8480
rect 33551 8449 33563 8452
rect 33505 8443 33563 8449
rect 34238 8440 34244 8452
rect 34296 8440 34302 8492
rect 34514 8489 34520 8492
rect 34508 8443 34520 8489
rect 34514 8440 34520 8443
rect 34572 8440 34578 8492
rect 35986 8440 35992 8492
rect 36044 8480 36050 8492
rect 36096 8489 36124 8520
rect 36081 8483 36139 8489
rect 36081 8480 36093 8483
rect 36044 8452 36093 8480
rect 36044 8440 36050 8452
rect 36081 8449 36093 8452
rect 36127 8449 36139 8483
rect 36081 8443 36139 8449
rect 36446 8440 36452 8492
rect 36504 8480 36510 8492
rect 36725 8483 36783 8489
rect 36725 8480 36737 8483
rect 36504 8452 36737 8480
rect 36504 8440 36510 8452
rect 36725 8449 36737 8452
rect 36771 8449 36783 8483
rect 36725 8443 36783 8449
rect 38378 8440 38384 8492
rect 38436 8489 38442 8492
rect 38436 8443 38448 8489
rect 38436 8440 38442 8443
rect 25133 8415 25191 8421
rect 25133 8381 25145 8415
rect 25179 8412 25191 8415
rect 25866 8412 25872 8424
rect 25179 8384 25872 8412
rect 25179 8381 25191 8384
rect 25133 8375 25191 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 27614 8372 27620 8424
rect 27672 8412 27678 8424
rect 27801 8415 27859 8421
rect 27801 8412 27813 8415
rect 27672 8384 27813 8412
rect 27672 8372 27678 8384
rect 27801 8381 27813 8384
rect 27847 8381 27859 8415
rect 29362 8412 29368 8424
rect 27801 8375 27859 8381
rect 29196 8384 29368 8412
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 16908 8316 17141 8344
rect 16908 8304 16914 8316
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17129 8307 17187 8313
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 26694 8344 26700 8356
rect 19300 8316 26700 8344
rect 19300 8304 19306 8316
rect 26694 8304 26700 8316
rect 26752 8304 26758 8356
rect 29196 8353 29224 8384
rect 29362 8372 29368 8384
rect 29420 8412 29426 8424
rect 30699 8415 30757 8421
rect 30699 8412 30711 8415
rect 29420 8384 30711 8412
rect 29420 8372 29426 8384
rect 30699 8381 30711 8384
rect 30745 8381 30757 8415
rect 30699 8375 30757 8381
rect 31757 8415 31815 8421
rect 31757 8381 31769 8415
rect 31803 8412 31815 8415
rect 31846 8412 31852 8424
rect 31803 8384 31852 8412
rect 31803 8381 31815 8384
rect 31757 8375 31815 8381
rect 31846 8372 31852 8384
rect 31904 8372 31910 8424
rect 32398 8372 32404 8424
rect 32456 8372 32462 8424
rect 35897 8415 35955 8421
rect 35897 8381 35909 8415
rect 35943 8412 35955 8415
rect 36464 8412 36492 8440
rect 35943 8384 36492 8412
rect 38580 8412 38608 8520
rect 38672 8520 40500 8548
rect 38672 8489 38700 8520
rect 40494 8508 40500 8520
rect 40552 8508 40558 8560
rect 45370 8548 45376 8560
rect 43548 8520 45376 8548
rect 43548 8492 43576 8520
rect 45370 8508 45376 8520
rect 45428 8508 45434 8560
rect 46100 8551 46158 8557
rect 46100 8517 46112 8551
rect 46146 8548 46158 8551
rect 46216 8548 46244 8576
rect 46146 8520 46244 8548
rect 47857 8551 47915 8557
rect 46146 8517 46158 8520
rect 46100 8511 46158 8517
rect 47857 8517 47869 8551
rect 47903 8548 47915 8551
rect 48240 8548 48268 8576
rect 47903 8520 48268 8548
rect 47903 8517 47915 8520
rect 47857 8511 47915 8517
rect 50154 8508 50160 8560
rect 50212 8548 50218 8560
rect 50709 8551 50767 8557
rect 50709 8548 50721 8551
rect 50212 8520 50721 8548
rect 50212 8508 50218 8520
rect 50709 8517 50721 8520
rect 50755 8517 50767 8551
rect 50709 8511 50767 8517
rect 38657 8483 38715 8489
rect 38657 8449 38669 8483
rect 38703 8449 38715 8483
rect 38657 8443 38715 8449
rect 38948 8452 39160 8480
rect 38948 8421 38976 8452
rect 38933 8415 38991 8421
rect 38580 8384 38700 8412
rect 35943 8381 35955 8384
rect 35897 8375 35955 8381
rect 29181 8347 29239 8353
rect 29181 8313 29193 8347
rect 29227 8313 29239 8347
rect 29181 8307 29239 8313
rect 29454 8304 29460 8356
rect 29512 8344 29518 8356
rect 29549 8347 29607 8353
rect 29549 8344 29561 8347
rect 29512 8316 29561 8344
rect 29512 8304 29518 8316
rect 29549 8313 29561 8316
rect 29595 8313 29607 8347
rect 29549 8307 29607 8313
rect 31113 8347 31171 8353
rect 31113 8313 31125 8347
rect 31159 8344 31171 8347
rect 31386 8344 31392 8356
rect 31159 8316 31392 8344
rect 31159 8313 31171 8316
rect 31113 8307 31171 8313
rect 31386 8304 31392 8316
rect 31444 8344 31450 8356
rect 32122 8344 32128 8356
rect 31444 8316 32128 8344
rect 31444 8304 31450 8316
rect 32122 8304 32128 8316
rect 32180 8344 32186 8356
rect 33781 8347 33839 8353
rect 33781 8344 33793 8347
rect 32180 8316 32628 8344
rect 32180 8304 32186 8316
rect 9861 8279 9919 8285
rect 9861 8276 9873 8279
rect 8956 8248 9873 8276
rect 5905 8239 5963 8245
rect 9861 8245 9873 8248
rect 9907 8245 9919 8279
rect 9861 8239 9919 8245
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12986 8276 12992 8288
rect 11848 8248 12992 8276
rect 11848 8236 11854 8248
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 17310 8236 17316 8288
rect 17368 8236 17374 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 20073 8279 20131 8285
rect 20073 8276 20085 8279
rect 19484 8248 20085 8276
rect 19484 8236 19490 8248
rect 20073 8245 20085 8248
rect 20119 8245 20131 8279
rect 20073 8239 20131 8245
rect 21634 8236 21640 8288
rect 21692 8236 21698 8288
rect 24026 8236 24032 8288
rect 24084 8276 24090 8288
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 24084 8248 24225 8276
rect 24084 8236 24090 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 32600 8276 32628 8316
rect 33520 8316 33793 8344
rect 33520 8276 33548 8316
rect 33781 8313 33793 8316
rect 33827 8313 33839 8347
rect 33781 8307 33839 8313
rect 38672 8344 38700 8384
rect 38933 8381 38945 8415
rect 38979 8381 38991 8415
rect 38933 8375 38991 8381
rect 39025 8415 39083 8421
rect 39025 8381 39037 8415
rect 39071 8381 39083 8415
rect 39132 8412 39160 8452
rect 39666 8440 39672 8492
rect 39724 8440 39730 8492
rect 40402 8440 40408 8492
rect 40460 8440 40466 8492
rect 43441 8483 43499 8489
rect 43441 8449 43453 8483
rect 43487 8480 43499 8483
rect 43530 8480 43536 8492
rect 43487 8452 43536 8480
rect 43487 8449 43499 8452
rect 43441 8443 43499 8449
rect 43530 8440 43536 8452
rect 43588 8440 43594 8492
rect 43708 8483 43766 8489
rect 43708 8449 43720 8483
rect 43754 8480 43766 8483
rect 44913 8483 44971 8489
rect 44913 8480 44925 8483
rect 43754 8452 44925 8480
rect 43754 8449 43766 8452
rect 43708 8443 43766 8449
rect 44913 8449 44925 8452
rect 44959 8449 44971 8483
rect 45388 8480 45416 8508
rect 45388 8452 45692 8480
rect 44913 8443 44971 8449
rect 40218 8412 40224 8424
rect 39132 8384 40224 8412
rect 39025 8375 39083 8381
rect 39040 8344 39068 8375
rect 40218 8372 40224 8384
rect 40276 8372 40282 8424
rect 38672 8316 39068 8344
rect 39485 8347 39543 8353
rect 32600 8248 33548 8276
rect 35621 8279 35679 8285
rect 24213 8239 24271 8245
rect 35621 8245 35633 8279
rect 35667 8276 35679 8279
rect 36078 8276 36084 8288
rect 35667 8248 36084 8276
rect 35667 8245 35679 8248
rect 35621 8239 35679 8245
rect 36078 8236 36084 8248
rect 36136 8276 36142 8288
rect 36722 8276 36728 8288
rect 36136 8248 36728 8276
rect 36136 8236 36142 8248
rect 36722 8236 36728 8248
rect 36780 8236 36786 8288
rect 37277 8279 37335 8285
rect 37277 8245 37289 8279
rect 37323 8276 37335 8279
rect 37734 8276 37740 8288
rect 37323 8248 37740 8276
rect 37323 8245 37335 8248
rect 37277 8239 37335 8245
rect 37734 8236 37740 8248
rect 37792 8236 37798 8288
rect 38286 8236 38292 8288
rect 38344 8276 38350 8288
rect 38672 8276 38700 8316
rect 39485 8313 39497 8347
rect 39531 8344 39543 8347
rect 40420 8344 40448 8440
rect 41414 8372 41420 8424
rect 41472 8372 41478 8424
rect 42242 8372 42248 8424
rect 42300 8372 42306 8424
rect 42518 8372 42524 8424
rect 42576 8412 42582 8424
rect 42981 8415 43039 8421
rect 42981 8412 42993 8415
rect 42576 8384 42993 8412
rect 42576 8372 42582 8384
rect 42981 8381 42993 8384
rect 43027 8381 43039 8415
rect 42981 8375 43039 8381
rect 45554 8372 45560 8424
rect 45612 8372 45618 8424
rect 45664 8412 45692 8452
rect 47946 8440 47952 8492
rect 48004 8440 48010 8492
rect 49050 8440 49056 8492
rect 49108 8440 49114 8492
rect 49326 8440 49332 8492
rect 49384 8440 49390 8492
rect 51046 8480 51074 8588
rect 51166 8576 51172 8628
rect 51224 8576 51230 8628
rect 52914 8576 52920 8628
rect 52972 8576 52978 8628
rect 54205 8619 54263 8625
rect 54205 8585 54217 8619
rect 54251 8616 54263 8619
rect 55214 8616 55220 8628
rect 54251 8588 55220 8616
rect 54251 8585 54263 8588
rect 54205 8579 54263 8585
rect 55214 8576 55220 8588
rect 55272 8576 55278 8628
rect 57609 8619 57667 8625
rect 57609 8585 57621 8619
rect 57655 8585 57667 8619
rect 57609 8579 57667 8585
rect 52457 8483 52515 8489
rect 52457 8480 52469 8483
rect 49896 8452 50476 8480
rect 51046 8452 52469 8480
rect 49896 8424 49924 8452
rect 45833 8415 45891 8421
rect 45833 8412 45845 8415
rect 45664 8384 45845 8412
rect 45833 8381 45845 8384
rect 45879 8381 45891 8415
rect 45833 8375 45891 8381
rect 47762 8372 47768 8424
rect 47820 8372 47826 8424
rect 49234 8421 49240 8424
rect 49212 8415 49240 8421
rect 49212 8381 49224 8415
rect 49212 8375 49240 8381
rect 49234 8372 49240 8375
rect 49292 8372 49298 8424
rect 49602 8372 49608 8424
rect 49660 8372 49666 8424
rect 49878 8372 49884 8424
rect 49936 8372 49942 8424
rect 50065 8415 50123 8421
rect 50065 8381 50077 8415
rect 50111 8381 50123 8415
rect 50065 8375 50123 8381
rect 39531 8316 40448 8344
rect 39531 8313 39543 8316
rect 39485 8307 39543 8313
rect 41506 8304 41512 8356
rect 41564 8344 41570 8356
rect 42429 8347 42487 8353
rect 42429 8344 42441 8347
rect 41564 8316 42441 8344
rect 41564 8304 41570 8316
rect 42429 8313 42441 8316
rect 42475 8313 42487 8347
rect 42429 8307 42487 8313
rect 38344 8248 38700 8276
rect 38344 8236 38350 8248
rect 40862 8236 40868 8288
rect 40920 8236 40926 8288
rect 41601 8279 41659 8285
rect 41601 8245 41613 8279
rect 41647 8276 41659 8279
rect 42150 8276 42156 8288
rect 41647 8248 42156 8276
rect 41647 8245 41659 8248
rect 41601 8239 41659 8245
rect 42150 8236 42156 8248
rect 42208 8236 42214 8288
rect 42334 8236 42340 8288
rect 42392 8276 42398 8288
rect 45370 8276 45376 8288
rect 42392 8248 45376 8276
rect 42392 8236 42398 8248
rect 45370 8236 45376 8248
rect 45428 8276 45434 8288
rect 47780 8276 47808 8372
rect 49620 8344 49648 8372
rect 50080 8344 50108 8375
rect 50246 8372 50252 8424
rect 50304 8372 50310 8424
rect 50448 8421 50476 8452
rect 52457 8449 52469 8452
rect 52503 8449 52515 8483
rect 52457 8443 52515 8449
rect 52733 8483 52791 8489
rect 52733 8449 52745 8483
rect 52779 8480 52791 8483
rect 52822 8480 52828 8492
rect 52779 8452 52828 8480
rect 52779 8449 52791 8452
rect 52733 8443 52791 8449
rect 52822 8440 52828 8452
rect 52880 8440 52886 8492
rect 52932 8480 52960 8576
rect 57624 8548 57652 8579
rect 57790 8576 57796 8628
rect 57848 8616 57854 8628
rect 57885 8619 57943 8625
rect 57885 8616 57897 8619
rect 57848 8588 57897 8616
rect 57848 8576 57854 8588
rect 57885 8585 57897 8588
rect 57931 8585 57943 8619
rect 57885 8579 57943 8585
rect 56060 8520 57652 8548
rect 52989 8483 53047 8489
rect 52989 8480 53001 8483
rect 52932 8452 53001 8480
rect 52989 8449 53001 8452
rect 53035 8449 53047 8483
rect 52989 8443 53047 8449
rect 54846 8440 54852 8492
rect 54904 8440 54910 8492
rect 56060 8489 56088 8520
rect 56045 8483 56103 8489
rect 56045 8449 56057 8483
rect 56091 8449 56103 8483
rect 56045 8443 56103 8449
rect 56318 8440 56324 8492
rect 56376 8480 56382 8492
rect 56485 8483 56543 8489
rect 56485 8480 56497 8483
rect 56376 8452 56497 8480
rect 56376 8440 56382 8452
rect 56485 8449 56497 8452
rect 56531 8449 56543 8483
rect 57624 8480 57652 8520
rect 58437 8483 58495 8489
rect 58437 8480 58449 8483
rect 57624 8452 58449 8480
rect 56485 8443 56543 8449
rect 58437 8449 58449 8452
rect 58483 8449 58495 8483
rect 58437 8443 58495 8449
rect 50433 8415 50491 8421
rect 50433 8381 50445 8415
rect 50479 8381 50491 8415
rect 51721 8415 51779 8421
rect 51721 8412 51733 8415
rect 50433 8375 50491 8381
rect 50724 8384 51733 8412
rect 50154 8344 50160 8356
rect 49620 8316 50016 8344
rect 50080 8316 50160 8344
rect 45428 8248 47808 8276
rect 45428 8236 45434 8248
rect 48314 8236 48320 8288
rect 48372 8236 48378 8288
rect 49988 8276 50016 8316
rect 50154 8304 50160 8316
rect 50212 8344 50218 8356
rect 50724 8344 50752 8384
rect 51721 8381 51733 8384
rect 51767 8381 51779 8415
rect 54662 8412 54668 8424
rect 51721 8375 51779 8381
rect 54128 8384 54668 8412
rect 50212 8316 50752 8344
rect 51077 8347 51135 8353
rect 50212 8304 50218 8316
rect 51077 8313 51089 8347
rect 51123 8344 51135 8347
rect 51258 8344 51264 8356
rect 51123 8316 51264 8344
rect 51123 8313 51135 8316
rect 51077 8307 51135 8313
rect 51258 8304 51264 8316
rect 51316 8304 51322 8356
rect 54128 8353 54156 8384
rect 54662 8372 54668 8384
rect 54720 8412 54726 8424
rect 54987 8415 55045 8421
rect 54987 8412 54999 8415
rect 54720 8384 54999 8412
rect 54720 8372 54726 8384
rect 54987 8381 54999 8384
rect 55033 8381 55045 8415
rect 54987 8375 55045 8381
rect 55122 8372 55128 8424
rect 55180 8372 55186 8424
rect 55306 8372 55312 8424
rect 55364 8412 55370 8424
rect 55401 8415 55459 8421
rect 55401 8412 55413 8415
rect 55364 8384 55413 8412
rect 55364 8372 55370 8384
rect 55401 8381 55413 8384
rect 55447 8381 55459 8415
rect 55401 8375 55459 8381
rect 55861 8415 55919 8421
rect 55861 8381 55873 8415
rect 55907 8412 55919 8415
rect 56134 8412 56140 8424
rect 55907 8384 56140 8412
rect 55907 8381 55919 8384
rect 55861 8375 55919 8381
rect 56134 8372 56140 8384
rect 56192 8372 56198 8424
rect 56229 8415 56287 8421
rect 56229 8381 56241 8415
rect 56275 8381 56287 8415
rect 56229 8375 56287 8381
rect 54113 8347 54171 8353
rect 51828 8316 52040 8344
rect 51828 8276 51856 8316
rect 49988 8248 51856 8276
rect 51902 8236 51908 8288
rect 51960 8236 51966 8288
rect 52012 8276 52040 8316
rect 54113 8313 54125 8347
rect 54159 8313 54171 8347
rect 54113 8307 54171 8313
rect 54018 8276 54024 8288
rect 52012 8248 54024 8276
rect 54018 8236 54024 8248
rect 54076 8276 54082 8288
rect 55324 8276 55352 8372
rect 54076 8248 55352 8276
rect 56244 8276 56272 8375
rect 57532 8316 57744 8344
rect 57532 8276 57560 8316
rect 57716 8288 57744 8316
rect 56244 8248 57560 8276
rect 54076 8236 54082 8248
rect 57698 8236 57704 8288
rect 57756 8236 57762 8288
rect 1104 8186 58880 8208
rect 1104 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 22616 8186
rect 22668 8134 22680 8186
rect 22732 8134 22744 8186
rect 22796 8134 22808 8186
rect 22860 8134 22872 8186
rect 22924 8134 37060 8186
rect 37112 8134 37124 8186
rect 37176 8134 37188 8186
rect 37240 8134 37252 8186
rect 37304 8134 37316 8186
rect 37368 8134 51504 8186
rect 51556 8134 51568 8186
rect 51620 8134 51632 8186
rect 51684 8134 51696 8186
rect 51748 8134 51760 8186
rect 51812 8134 58880 8186
rect 1104 8112 58880 8134
rect 3878 8032 3884 8084
rect 3936 8032 3942 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4028 8044 4445 8072
rect 4028 8032 4034 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 8754 8072 8760 8084
rect 6328 8044 8760 8072
rect 6328 8032 6334 8044
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 4663 7976 5212 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3694 7868 3700 7880
rect 2832 7840 3700 7868
rect 2832 7828 2838 7840
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4338 7868 4344 7880
rect 4019 7840 4344 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 5184 7877 5212 7976
rect 7742 7964 7748 8016
rect 7800 7964 7806 8016
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5810 7868 5816 7880
rect 5215 7840 5816 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 7760 7868 7788 7964
rect 7852 7945 7880 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10836 8044 10885 8072
rect 10836 8032 10842 8044
rect 10873 8041 10885 8044
rect 10919 8072 10931 8075
rect 11790 8072 11796 8084
rect 10919 8044 11796 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12158 8072 12164 8084
rect 11931 8044 12164 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 13354 8072 13360 8084
rect 12452 8044 13360 8072
rect 8297 8007 8355 8013
rect 8297 7973 8309 8007
rect 8343 7973 8355 8007
rect 8846 8004 8852 8016
rect 8297 7967 8355 7973
rect 8404 7976 8852 8004
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 8312 7880 8340 7967
rect 8404 7945 8432 7976
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 12452 8004 12480 8044
rect 13354 8032 13360 8044
rect 13412 8072 13418 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13412 8044 13645 8072
rect 13412 8032 13418 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 13740 8044 17908 8072
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 12406 7976 12480 8004
rect 12544 7976 12633 8004
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 12406 7936 12434 7976
rect 12544 7945 12572 7976
rect 12621 7973 12633 7976
rect 12667 7973 12679 8007
rect 13740 8004 13768 8044
rect 17880 8004 17908 8044
rect 17954 8032 17960 8084
rect 18012 8032 18018 8084
rect 18064 8044 33364 8072
rect 18064 8004 18092 8044
rect 12621 7967 12679 7973
rect 12728 7976 13768 8004
rect 15120 7976 17448 8004
rect 17880 7976 18092 8004
rect 18693 8007 18751 8013
rect 8803 7908 12434 7936
rect 12529 7939 12587 7945
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12728 7936 12756 7976
rect 15120 7948 15148 7976
rect 12529 7899 12587 7905
rect 12616 7908 12756 7936
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7760 7840 7941 7868
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 3421 7803 3479 7809
rect 3421 7769 3433 7803
rect 3467 7800 3479 7803
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 3467 7772 4261 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 4249 7769 4261 7772
rect 4295 7800 4307 7803
rect 4706 7800 4712 7812
rect 4295 7772 4712 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 5353 7803 5411 7809
rect 5353 7769 5365 7803
rect 5399 7800 5411 7803
rect 6104 7800 6132 7828
rect 7944 7800 7972 7831
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8404 7868 8432 7899
rect 8478 7868 8484 7880
rect 8404 7840 8484 7868
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 8720 7840 9229 7868
rect 8720 7828 8726 7840
rect 9217 7837 9229 7840
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9548 7840 9689 7868
rect 9548 7828 9554 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 12616 7868 12644 7908
rect 13078 7896 13084 7948
rect 13136 7936 13142 7948
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 13136 7908 13185 7936
rect 13136 7896 13142 7908
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 14826 7936 14832 7948
rect 14783 7908 14832 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15194 7896 15200 7948
rect 15252 7896 15258 7948
rect 16574 7896 16580 7948
rect 16632 7896 16638 7948
rect 17310 7896 17316 7948
rect 17368 7896 17374 7948
rect 17420 7936 17448 7976
rect 18693 7973 18705 8007
rect 18739 8004 18751 8007
rect 19334 8004 19340 8016
rect 18739 7976 19340 8004
rect 18739 7973 18751 7976
rect 18693 7967 18751 7973
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 22278 7964 22284 8016
rect 22336 8004 22342 8016
rect 22557 8007 22615 8013
rect 22557 8004 22569 8007
rect 22336 7976 22569 8004
rect 22336 7964 22342 7976
rect 22557 7973 22569 7976
rect 22603 8004 22615 8007
rect 24118 8004 24124 8016
rect 22603 7976 24124 8004
rect 22603 7973 22615 7976
rect 22557 7967 22615 7973
rect 24118 7964 24124 7976
rect 24176 7964 24182 8016
rect 25314 7964 25320 8016
rect 25372 8004 25378 8016
rect 25774 8004 25780 8016
rect 25372 7976 25780 8004
rect 25372 7964 25378 7976
rect 25774 7964 25780 7976
rect 25832 7964 25838 8016
rect 32769 8007 32827 8013
rect 31036 7976 32720 8004
rect 18966 7936 18972 7948
rect 17420 7908 18972 7936
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 29362 7896 29368 7948
rect 29420 7896 29426 7948
rect 29748 7908 30144 7936
rect 12406 7840 12644 7868
rect 9125 7803 9183 7809
rect 9125 7800 9137 7803
rect 5399 7772 6132 7800
rect 6196 7772 7696 7800
rect 7944 7772 9137 7800
rect 5399 7769 5411 7772
rect 5353 7763 5411 7769
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 4459 7735 4517 7741
rect 4459 7732 4471 7735
rect 4120 7704 4471 7732
rect 4120 7692 4126 7704
rect 4459 7701 4471 7704
rect 4505 7701 4517 7735
rect 4459 7695 4517 7701
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 6196 7732 6224 7772
rect 5500 7704 6224 7732
rect 7285 7735 7343 7741
rect 5500 7692 5506 7704
rect 7285 7701 7297 7735
rect 7331 7732 7343 7735
rect 7374 7732 7380 7744
rect 7331 7704 7380 7732
rect 7331 7701 7343 7704
rect 7285 7695 7343 7701
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7524 7704 7573 7732
rect 7524 7692 7530 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7668 7732 7696 7772
rect 9125 7769 9137 7772
rect 9171 7769 9183 7803
rect 9125 7763 9183 7769
rect 9582 7760 9588 7812
rect 9640 7760 9646 7812
rect 12406 7800 12434 7840
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12768 7840 13001 7868
rect 12768 7828 12774 7840
rect 12989 7837 13001 7840
rect 13035 7868 13047 7871
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 13035 7840 15485 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 15473 7837 15485 7840
rect 15519 7868 15531 7871
rect 17770 7868 17776 7880
rect 15519 7840 17776 7868
rect 15519 7837 15531 7840
rect 15473 7831 15531 7837
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 20588 7840 20637 7868
rect 20588 7828 20594 7840
rect 20625 7837 20637 7840
rect 20671 7868 20683 7871
rect 20806 7868 20812 7880
rect 20671 7840 20812 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 26510 7828 26516 7880
rect 26568 7828 26574 7880
rect 26694 7828 26700 7880
rect 26752 7868 26758 7880
rect 26881 7871 26939 7877
rect 26881 7868 26893 7871
rect 26752 7840 26893 7868
rect 26752 7828 26758 7840
rect 26881 7837 26893 7840
rect 26927 7837 26939 7871
rect 26881 7831 26939 7837
rect 9692 7772 12434 7800
rect 13081 7803 13139 7809
rect 9692 7732 9720 7772
rect 13081 7769 13093 7803
rect 13127 7800 13139 7803
rect 14093 7803 14151 7809
rect 14093 7800 14105 7803
rect 13127 7772 14105 7800
rect 13127 7769 13139 7772
rect 13081 7763 13139 7769
rect 14093 7769 14105 7772
rect 14139 7769 14151 7803
rect 14093 7763 14151 7769
rect 15381 7803 15439 7809
rect 15381 7769 15393 7803
rect 15427 7800 15439 7803
rect 15933 7803 15991 7809
rect 15933 7800 15945 7803
rect 15427 7772 15945 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 15933 7769 15945 7772
rect 15979 7769 15991 7803
rect 15933 7763 15991 7769
rect 18138 7760 18144 7812
rect 18196 7800 18202 7812
rect 18509 7803 18567 7809
rect 18509 7800 18521 7803
rect 18196 7772 18521 7800
rect 18196 7760 18202 7772
rect 18509 7769 18521 7772
rect 18555 7769 18567 7803
rect 18509 7763 18567 7769
rect 20380 7803 20438 7809
rect 20380 7769 20392 7803
rect 20426 7800 20438 7803
rect 20717 7803 20775 7809
rect 20717 7800 20729 7803
rect 20426 7772 20729 7800
rect 20426 7769 20438 7772
rect 20380 7763 20438 7769
rect 20717 7769 20729 7772
rect 20763 7769 20775 7803
rect 29748 7800 29776 7908
rect 30009 7871 30067 7877
rect 30009 7868 30021 7871
rect 20717 7763 20775 7769
rect 20824 7772 29776 7800
rect 29840 7840 30021 7868
rect 7668 7704 9720 7732
rect 7561 7695 7619 7701
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 11054 7692 11060 7744
rect 11112 7692 11118 7744
rect 15838 7692 15844 7744
rect 15896 7692 15902 7744
rect 19150 7692 19156 7744
rect 19208 7732 19214 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 19208 7704 19257 7732
rect 19208 7692 19214 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 20622 7692 20628 7744
rect 20680 7732 20686 7744
rect 20824 7732 20852 7772
rect 20680 7704 20852 7732
rect 20680 7692 20686 7704
rect 23014 7692 23020 7744
rect 23072 7692 23078 7744
rect 24026 7692 24032 7744
rect 24084 7692 24090 7744
rect 25958 7692 25964 7744
rect 26016 7692 26022 7744
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 28169 7735 28227 7741
rect 28169 7732 28181 7735
rect 27672 7704 28181 7732
rect 27672 7692 27678 7704
rect 28169 7701 28181 7704
rect 28215 7701 28227 7735
rect 28169 7695 28227 7701
rect 28718 7692 28724 7744
rect 28776 7692 28782 7744
rect 29454 7692 29460 7744
rect 29512 7732 29518 7744
rect 29840 7741 29868 7840
rect 30009 7837 30021 7840
rect 30055 7837 30067 7871
rect 30116 7868 30144 7908
rect 31036 7868 31064 7976
rect 32692 7948 32720 7976
rect 32769 7973 32781 8007
rect 32815 7973 32827 8007
rect 33336 8004 33364 8044
rect 33410 8032 33416 8084
rect 33468 8072 33474 8084
rect 33597 8075 33655 8081
rect 33597 8072 33609 8075
rect 33468 8044 33609 8072
rect 33468 8032 33474 8044
rect 33597 8041 33609 8044
rect 33643 8041 33655 8075
rect 38470 8072 38476 8084
rect 33597 8035 33655 8041
rect 36280 8044 38476 8072
rect 36280 8004 36308 8044
rect 38470 8032 38476 8044
rect 38528 8032 38534 8084
rect 41690 8072 41696 8084
rect 38626 8044 41696 8072
rect 38626 8004 38654 8044
rect 41690 8032 41696 8044
rect 41748 8032 41754 8084
rect 41785 8075 41843 8081
rect 41785 8041 41797 8075
rect 41831 8072 41843 8075
rect 42518 8072 42524 8084
rect 41831 8044 42524 8072
rect 41831 8041 41843 8044
rect 41785 8035 41843 8041
rect 42518 8032 42524 8044
rect 42576 8032 42582 8084
rect 44729 8075 44787 8081
rect 44729 8041 44741 8075
rect 44775 8072 44787 8075
rect 45554 8072 45560 8084
rect 44775 8044 45560 8072
rect 44775 8041 44787 8044
rect 44729 8035 44787 8041
rect 45554 8032 45560 8044
rect 45612 8032 45618 8084
rect 47946 8032 47952 8084
rect 48004 8032 48010 8084
rect 49513 8075 49571 8081
rect 49513 8041 49525 8075
rect 49559 8072 49571 8075
rect 50246 8072 50252 8084
rect 49559 8044 50252 8072
rect 49559 8041 49571 8044
rect 49513 8035 49571 8041
rect 50246 8032 50252 8044
rect 50304 8032 50310 8084
rect 52822 8072 52828 8084
rect 52564 8044 52828 8072
rect 44818 8004 44824 8016
rect 33336 7976 36308 8004
rect 38488 7976 38654 8004
rect 44192 7976 44824 8004
rect 32769 7967 32827 7973
rect 31754 7896 31760 7948
rect 31812 7896 31818 7948
rect 32214 7896 32220 7948
rect 32272 7896 32278 7948
rect 32309 7939 32367 7945
rect 32309 7905 32321 7939
rect 32355 7936 32367 7939
rect 32490 7936 32496 7948
rect 32355 7908 32496 7936
rect 32355 7905 32367 7908
rect 32309 7899 32367 7905
rect 32490 7896 32496 7908
rect 32548 7896 32554 7948
rect 32674 7896 32680 7948
rect 32732 7896 32738 7948
rect 32784 7936 32812 7967
rect 34149 7939 34207 7945
rect 34149 7936 34161 7939
rect 32784 7908 34161 7936
rect 34149 7905 34161 7908
rect 34195 7905 34207 7939
rect 34149 7899 34207 7905
rect 35529 7939 35587 7945
rect 35529 7905 35541 7939
rect 35575 7936 35587 7939
rect 35710 7936 35716 7948
rect 35575 7908 35716 7936
rect 35575 7905 35587 7908
rect 35529 7899 35587 7905
rect 35710 7896 35716 7908
rect 35768 7896 35774 7948
rect 35986 7896 35992 7948
rect 36044 7896 36050 7948
rect 36446 7896 36452 7948
rect 36504 7936 36510 7948
rect 36504 7908 36676 7936
rect 36504 7896 36510 7908
rect 30116 7840 31064 7868
rect 32401 7871 32459 7877
rect 30009 7831 30067 7837
rect 32401 7837 32413 7871
rect 32447 7868 32459 7871
rect 32858 7868 32864 7880
rect 32447 7840 32864 7868
rect 32447 7837 32459 7840
rect 32401 7831 32459 7837
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 33413 7871 33471 7877
rect 33413 7837 33425 7871
rect 33459 7837 33471 7871
rect 33413 7831 33471 7837
rect 35345 7871 35403 7877
rect 35345 7837 35357 7871
rect 35391 7868 35403 7871
rect 36004 7868 36032 7896
rect 36648 7877 36676 7908
rect 36906 7896 36912 7948
rect 36964 7896 36970 7948
rect 37182 7896 37188 7948
rect 37240 7896 37246 7948
rect 37642 7896 37648 7948
rect 37700 7896 37706 7948
rect 37734 7896 37740 7948
rect 37792 7936 37798 7948
rect 37829 7939 37887 7945
rect 37829 7936 37841 7939
rect 37792 7908 37841 7936
rect 37792 7896 37798 7908
rect 37829 7905 37841 7908
rect 37875 7905 37887 7939
rect 37829 7899 37887 7905
rect 35391 7840 36032 7868
rect 36633 7871 36691 7877
rect 35391 7837 35403 7840
rect 35345 7831 35403 7837
rect 36633 7837 36645 7871
rect 36679 7837 36691 7871
rect 36633 7831 36691 7837
rect 30276 7803 30334 7809
rect 30276 7769 30288 7803
rect 30322 7800 30334 7803
rect 30466 7800 30472 7812
rect 30322 7772 30472 7800
rect 30322 7769 30334 7772
rect 30276 7763 30334 7769
rect 30466 7760 30472 7772
rect 30524 7760 30530 7812
rect 31846 7800 31852 7812
rect 31726 7772 31852 7800
rect 29825 7735 29883 7741
rect 29825 7732 29837 7735
rect 29512 7704 29837 7732
rect 29512 7692 29518 7704
rect 29825 7701 29837 7704
rect 29871 7701 29883 7735
rect 29825 7695 29883 7701
rect 31389 7735 31447 7741
rect 31389 7701 31401 7735
rect 31435 7732 31447 7735
rect 31726 7732 31754 7772
rect 31846 7760 31852 7772
rect 31904 7800 31910 7812
rect 33428 7800 33456 7831
rect 36722 7828 36728 7880
rect 36780 7877 36786 7880
rect 36780 7871 36829 7877
rect 36780 7837 36783 7871
rect 36817 7837 36829 7871
rect 37844 7868 37872 7899
rect 38010 7896 38016 7948
rect 38068 7936 38074 7948
rect 38488 7945 38516 7976
rect 44192 7945 44220 7976
rect 44818 7964 44824 7976
rect 44876 8004 44882 8016
rect 45186 8004 45192 8016
rect 44876 7976 45192 8004
rect 44876 7964 44882 7976
rect 45186 7964 45192 7976
rect 45244 7964 45250 8016
rect 50154 7964 50160 8016
rect 50212 7964 50218 8016
rect 38473 7939 38531 7945
rect 38473 7936 38485 7939
rect 38068 7908 38485 7936
rect 38068 7896 38074 7908
rect 38473 7905 38485 7908
rect 38519 7905 38531 7939
rect 38473 7899 38531 7905
rect 44177 7939 44235 7945
rect 44177 7905 44189 7939
rect 44223 7905 44235 7939
rect 44177 7899 44235 7905
rect 44634 7896 44640 7948
rect 44692 7936 44698 7948
rect 52564 7945 52592 8044
rect 52822 8032 52828 8044
rect 52880 8032 52886 8084
rect 53929 8075 53987 8081
rect 53929 8041 53941 8075
rect 53975 8072 53987 8075
rect 55122 8072 55128 8084
rect 53975 8044 55128 8072
rect 53975 8041 53987 8044
rect 53929 8035 53987 8041
rect 55122 8032 55128 8044
rect 55180 8032 55186 8084
rect 54938 8004 54944 8016
rect 53760 7976 54944 8004
rect 45557 7939 45615 7945
rect 45557 7936 45569 7939
rect 44692 7908 45569 7936
rect 44692 7896 44698 7908
rect 45557 7905 45569 7908
rect 45603 7905 45615 7939
rect 45557 7899 45615 7905
rect 47213 7939 47271 7945
rect 47213 7905 47225 7939
rect 47259 7936 47271 7939
rect 51537 7939 51595 7945
rect 47259 7908 48176 7936
rect 47259 7905 47271 7908
rect 47213 7899 47271 7905
rect 39301 7871 39359 7877
rect 39301 7868 39313 7871
rect 37844 7840 39313 7868
rect 36780 7831 36829 7837
rect 39301 7837 39313 7840
rect 39347 7837 39359 7871
rect 39301 7831 39359 7837
rect 40405 7871 40463 7877
rect 40405 7837 40417 7871
rect 40451 7868 40463 7871
rect 40494 7868 40500 7880
rect 40451 7840 40500 7868
rect 40451 7837 40463 7840
rect 40405 7831 40463 7837
rect 36780 7828 36786 7831
rect 40494 7828 40500 7840
rect 40552 7868 40558 7880
rect 41877 7871 41935 7877
rect 41877 7868 41889 7871
rect 40552 7840 41889 7868
rect 40552 7828 40558 7840
rect 41877 7837 41889 7840
rect 41923 7868 41935 7871
rect 41966 7868 41972 7880
rect 41923 7840 41972 7868
rect 41923 7837 41935 7840
rect 41877 7831 41935 7837
rect 41966 7828 41972 7840
rect 42024 7828 42030 7880
rect 42150 7877 42156 7880
rect 42144 7868 42156 7877
rect 42111 7840 42156 7868
rect 42144 7831 42156 7840
rect 42150 7828 42156 7831
rect 42208 7828 42214 7880
rect 48148 7877 48176 7908
rect 51537 7905 51549 7939
rect 51583 7936 51595 7939
rect 52549 7939 52607 7945
rect 52549 7936 52561 7939
rect 51583 7908 52561 7936
rect 51583 7905 51595 7908
rect 51537 7899 51595 7905
rect 52549 7905 52561 7908
rect 52595 7905 52607 7939
rect 52549 7899 52607 7905
rect 47397 7871 47455 7877
rect 43180 7840 46520 7868
rect 31904 7772 33456 7800
rect 31904 7760 31910 7772
rect 38286 7760 38292 7812
rect 38344 7760 38350 7812
rect 40037 7803 40095 7809
rect 40037 7769 40049 7803
rect 40083 7800 40095 7803
rect 40310 7800 40316 7812
rect 40083 7772 40316 7800
rect 40083 7769 40095 7772
rect 40037 7763 40095 7769
rect 40310 7760 40316 7772
rect 40368 7760 40374 7812
rect 40672 7803 40730 7809
rect 40672 7769 40684 7803
rect 40718 7800 40730 7803
rect 40862 7800 40868 7812
rect 40718 7772 40868 7800
rect 40718 7769 40730 7772
rect 40672 7763 40730 7769
rect 40862 7760 40868 7772
rect 40920 7760 40926 7812
rect 31435 7704 31754 7732
rect 31435 7701 31447 7704
rect 31389 7695 31447 7701
rect 32306 7692 32312 7744
rect 32364 7732 32370 7744
rect 32861 7735 32919 7741
rect 32861 7732 32873 7735
rect 32364 7704 32873 7732
rect 32364 7692 32370 7704
rect 32861 7701 32873 7704
rect 32907 7701 32919 7735
rect 32861 7695 32919 7701
rect 34882 7692 34888 7744
rect 34940 7692 34946 7744
rect 35250 7692 35256 7744
rect 35308 7692 35314 7744
rect 35989 7735 36047 7741
rect 35989 7701 36001 7735
rect 36035 7732 36047 7735
rect 37642 7732 37648 7744
rect 36035 7704 37648 7732
rect 36035 7701 36047 7704
rect 35989 7695 36047 7701
rect 37642 7692 37648 7704
rect 37700 7692 37706 7744
rect 37918 7692 37924 7744
rect 37976 7692 37982 7744
rect 38381 7735 38439 7741
rect 38381 7701 38393 7735
rect 38427 7732 38439 7735
rect 38749 7735 38807 7741
rect 38749 7732 38761 7735
rect 38427 7704 38761 7732
rect 38427 7701 38439 7704
rect 38381 7695 38439 7701
rect 38749 7701 38761 7704
rect 38795 7701 38807 7735
rect 38749 7695 38807 7701
rect 39022 7692 39028 7744
rect 39080 7732 39086 7744
rect 43180 7732 43208 7840
rect 46492 7812 46520 7840
rect 47397 7837 47409 7871
rect 47443 7868 47455 7871
rect 48133 7871 48191 7877
rect 47443 7840 47716 7868
rect 47443 7837 47455 7840
rect 47397 7831 47455 7837
rect 44361 7803 44419 7809
rect 44361 7769 44373 7803
rect 44407 7800 44419 7803
rect 45005 7803 45063 7809
rect 45005 7800 45017 7803
rect 44407 7772 45017 7800
rect 44407 7769 44419 7772
rect 44361 7763 44419 7769
rect 45005 7769 45017 7772
rect 45051 7769 45063 7803
rect 45005 7763 45063 7769
rect 46474 7760 46480 7812
rect 46532 7760 46538 7812
rect 46968 7803 47026 7809
rect 46968 7769 46980 7803
rect 47014 7800 47026 7803
rect 47578 7800 47584 7812
rect 47014 7772 47584 7800
rect 47014 7769 47026 7772
rect 46968 7763 47026 7769
rect 47578 7760 47584 7772
rect 47636 7760 47642 7812
rect 39080 7704 43208 7732
rect 39080 7692 39086 7704
rect 43254 7692 43260 7744
rect 43312 7692 43318 7744
rect 43625 7735 43683 7741
rect 43625 7701 43637 7735
rect 43671 7732 43683 7735
rect 43990 7732 43996 7744
rect 43671 7704 43996 7732
rect 43671 7701 43683 7704
rect 43625 7695 43683 7701
rect 43990 7692 43996 7704
rect 44048 7692 44054 7744
rect 44174 7692 44180 7744
rect 44232 7732 44238 7744
rect 44269 7735 44327 7741
rect 44269 7732 44281 7735
rect 44232 7704 44281 7732
rect 44232 7692 44238 7704
rect 44269 7701 44281 7704
rect 44315 7732 44327 7735
rect 45462 7732 45468 7744
rect 44315 7704 45468 7732
rect 44315 7701 44327 7704
rect 44269 7695 44327 7701
rect 45462 7692 45468 7704
rect 45520 7692 45526 7744
rect 45833 7735 45891 7741
rect 45833 7701 45845 7735
rect 45879 7732 45891 7735
rect 47688 7732 47716 7840
rect 48133 7837 48145 7871
rect 48179 7868 48191 7871
rect 51552 7868 51580 7899
rect 48179 7840 51580 7868
rect 48179 7837 48191 7840
rect 48133 7831 48191 7837
rect 51902 7828 51908 7880
rect 51960 7828 51966 7880
rect 52457 7871 52515 7877
rect 52457 7837 52469 7871
rect 52503 7868 52515 7871
rect 53760 7868 53788 7976
rect 54938 7964 54944 7976
rect 54996 7964 55002 8016
rect 53926 7896 53932 7948
rect 53984 7936 53990 7948
rect 54573 7939 54631 7945
rect 54573 7936 54585 7939
rect 53984 7908 54585 7936
rect 53984 7896 53990 7908
rect 54573 7905 54585 7908
rect 54619 7905 54631 7939
rect 54573 7899 54631 7905
rect 55214 7896 55220 7948
rect 55272 7936 55278 7948
rect 55769 7939 55827 7945
rect 55769 7936 55781 7939
rect 55272 7908 55781 7936
rect 55272 7896 55278 7908
rect 55769 7905 55781 7908
rect 55815 7905 55827 7939
rect 55769 7899 55827 7905
rect 55858 7896 55864 7948
rect 55916 7896 55922 7948
rect 57698 7896 57704 7948
rect 57756 7896 57762 7948
rect 58066 7896 58072 7948
rect 58124 7936 58130 7948
rect 58345 7939 58403 7945
rect 58345 7936 58357 7939
rect 58124 7908 58357 7936
rect 58124 7896 58130 7908
rect 58345 7905 58357 7908
rect 58391 7905 58403 7939
rect 58345 7899 58403 7905
rect 52503 7840 53788 7868
rect 52503 7837 52515 7840
rect 52457 7831 52515 7837
rect 54478 7828 54484 7880
rect 54536 7868 54542 7880
rect 55677 7871 55735 7877
rect 55677 7868 55689 7871
rect 54536 7840 55689 7868
rect 54536 7828 54542 7840
rect 55677 7837 55689 7840
rect 55723 7837 55735 7871
rect 55677 7831 55735 7837
rect 48400 7803 48458 7809
rect 48400 7769 48412 7803
rect 48446 7800 48458 7803
rect 48590 7800 48596 7812
rect 48446 7772 48596 7800
rect 48446 7769 48458 7772
rect 48400 7763 48458 7769
rect 48590 7760 48596 7772
rect 48648 7760 48654 7812
rect 49234 7760 49240 7812
rect 49292 7760 49298 7812
rect 51292 7803 51350 7809
rect 51292 7769 51304 7803
rect 51338 7800 51350 7803
rect 51920 7800 51948 7828
rect 51338 7772 51948 7800
rect 52816 7803 52874 7809
rect 51338 7769 51350 7772
rect 51292 7763 51350 7769
rect 52816 7769 52828 7803
rect 52862 7800 52874 7803
rect 54021 7803 54079 7809
rect 54021 7800 54033 7803
rect 52862 7772 54033 7800
rect 52862 7769 52874 7772
rect 52816 7763 52874 7769
rect 54021 7769 54033 7772
rect 54067 7769 54079 7803
rect 54021 7763 54079 7769
rect 57456 7803 57514 7809
rect 57456 7769 57468 7803
rect 57502 7800 57514 7803
rect 57793 7803 57851 7809
rect 57793 7800 57805 7803
rect 57502 7772 57805 7800
rect 57502 7769 57514 7772
rect 57456 7763 57514 7769
rect 57793 7769 57805 7772
rect 57839 7769 57851 7803
rect 57793 7763 57851 7769
rect 49252 7732 49280 7760
rect 45879 7704 49280 7732
rect 45879 7701 45891 7704
rect 45833 7695 45891 7701
rect 49878 7692 49884 7744
rect 49936 7692 49942 7744
rect 51994 7692 52000 7744
rect 52052 7692 52058 7744
rect 55306 7692 55312 7744
rect 55364 7692 55370 7744
rect 56134 7692 56140 7744
rect 56192 7732 56198 7744
rect 56321 7735 56379 7741
rect 56321 7732 56333 7735
rect 56192 7704 56333 7732
rect 56192 7692 56198 7704
rect 56321 7701 56333 7704
rect 56367 7732 56379 7735
rect 56502 7732 56508 7744
rect 56367 7704 56508 7732
rect 56367 7701 56379 7704
rect 56321 7695 56379 7701
rect 56502 7692 56508 7704
rect 56560 7692 56566 7744
rect 1104 7642 59040 7664
rect 1104 7590 15394 7642
rect 15446 7590 15458 7642
rect 15510 7590 15522 7642
rect 15574 7590 15586 7642
rect 15638 7590 15650 7642
rect 15702 7590 29838 7642
rect 29890 7590 29902 7642
rect 29954 7590 29966 7642
rect 30018 7590 30030 7642
rect 30082 7590 30094 7642
rect 30146 7590 44282 7642
rect 44334 7590 44346 7642
rect 44398 7590 44410 7642
rect 44462 7590 44474 7642
rect 44526 7590 44538 7642
rect 44590 7590 58726 7642
rect 58778 7590 58790 7642
rect 58842 7590 58854 7642
rect 58906 7590 58918 7642
rect 58970 7590 58982 7642
rect 59034 7590 59040 7642
rect 1104 7568 59040 7590
rect 5813 7531 5871 7537
rect 3712 7500 5212 7528
rect 2593 7463 2651 7469
rect 2593 7429 2605 7463
rect 2639 7460 2651 7463
rect 3418 7460 3424 7472
rect 2639 7432 3424 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 3712 7460 3740 7500
rect 3528 7432 3740 7460
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 3528 7401 3556 7432
rect 3712 7401 3740 7432
rect 4522 7420 4528 7472
rect 4580 7420 4586 7472
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3620 7324 3648 7355
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4724 7324 4752 7352
rect 3620 7296 4752 7324
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4948 7296 4997 7324
rect 4948 7284 4954 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5074 7284 5080 7336
rect 5132 7284 5138 7336
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 2608 7228 2881 7256
rect 2608 7197 2636 7228
rect 2869 7225 2881 7228
rect 2915 7225 2927 7259
rect 4338 7256 4344 7268
rect 2869 7219 2927 7225
rect 3620 7228 4344 7256
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7157 2651 7191
rect 2593 7151 2651 7157
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3620 7188 3648 7228
rect 4338 7216 4344 7228
rect 4396 7216 4402 7268
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7225 4583 7259
rect 5184 7256 5212 7500
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 5994 7528 6000 7540
rect 5859 7500 6000 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9640 7488 9674 7528
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 11296 7500 12817 7528
rect 11296 7488 11302 7500
rect 12805 7497 12817 7500
rect 12851 7528 12863 7531
rect 14274 7528 14280 7540
rect 12851 7500 14280 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 14274 7488 14280 7500
rect 14332 7528 14338 7540
rect 14826 7528 14832 7540
rect 14332 7500 14832 7528
rect 14332 7488 14338 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14976 7500 15025 7528
rect 14976 7488 14982 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 20622 7528 20628 7540
rect 16632 7500 20628 7528
rect 16632 7488 16638 7500
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 20732 7500 25452 7528
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 8662 7460 8668 7472
rect 5307 7432 8668 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 9646 7460 9674 7488
rect 10597 7463 10655 7469
rect 10597 7460 10609 7463
rect 8772 7432 8984 7460
rect 9646 7432 10609 7460
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 6687 7364 7328 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7300 7336 7328 7364
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8772 7392 8800 7432
rect 7800 7364 8800 7392
rect 8849 7395 8907 7401
rect 7800 7352 7806 7364
rect 7190 7284 7196 7336
rect 7248 7284 7254 7336
rect 7282 7284 7288 7336
rect 7340 7284 7346 7336
rect 8110 7284 8116 7336
rect 8168 7284 8174 7336
rect 8220 7333 8248 7364
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8956 7392 8984 7432
rect 10597 7429 10609 7432
rect 10643 7460 10655 7463
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10643 7432 11529 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 11517 7429 11529 7432
rect 11563 7460 11575 7463
rect 11563 7432 14596 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 9079 7395 9137 7401
rect 9079 7392 9091 7395
rect 8956 7364 9091 7392
rect 8849 7355 8907 7361
rect 9079 7361 9091 7364
rect 9125 7361 9137 7395
rect 9079 7355 9137 7361
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8864 7324 8892 7355
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9640 7364 9965 7392
rect 9640 7352 9646 7364
rect 9953 7361 9965 7364
rect 9999 7392 10011 7395
rect 9999 7364 13492 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 8352 7296 8892 7324
rect 8956 7296 9229 7324
rect 8352 7284 8358 7296
rect 8404 7265 8432 7296
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 5184 7228 8401 7256
rect 4525 7219 4583 7225
rect 8389 7225 8401 7228
rect 8435 7225 8447 7259
rect 8389 7219 8447 7225
rect 2823 7160 3648 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 4540 7188 4568 7219
rect 8754 7216 8760 7268
rect 8812 7256 8818 7268
rect 8956 7256 8984 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 10827 7296 12434 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 8812 7228 8984 7256
rect 12406 7256 12434 7296
rect 13357 7259 13415 7265
rect 13357 7256 13369 7259
rect 12406 7228 13369 7256
rect 8812 7216 8818 7228
rect 13357 7225 13369 7228
rect 13403 7225 13415 7259
rect 13464 7256 13492 7364
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 14568 7392 14596 7432
rect 15396 7432 20576 7460
rect 15396 7392 15424 7432
rect 14568 7364 15424 7392
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 15838 7392 15844 7404
rect 15703 7364 15844 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16574 7352 16580 7404
rect 16632 7352 16638 7404
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17770 7392 17776 7404
rect 17635 7364 17776 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17770 7352 17776 7364
rect 17828 7352 17834 7404
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19518 7352 19524 7404
rect 19576 7352 19582 7404
rect 20548 7392 20576 7432
rect 20732 7392 20760 7500
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 21358 7460 21364 7472
rect 20864 7432 21364 7460
rect 20864 7420 20870 7432
rect 21358 7420 21364 7432
rect 21416 7460 21422 7472
rect 21634 7460 21640 7472
rect 21416 7432 21640 7460
rect 21416 7420 21422 7432
rect 21634 7420 21640 7432
rect 21692 7460 21698 7472
rect 21692 7432 24072 7460
rect 21692 7420 21698 7432
rect 22204 7401 22232 7432
rect 24044 7404 24072 7432
rect 24118 7420 24124 7472
rect 24176 7460 24182 7472
rect 24670 7460 24676 7472
rect 24176 7432 24676 7460
rect 24176 7420 24182 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 20548 7364 20760 7392
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22456 7395 22514 7401
rect 22235 7364 22269 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22456 7361 22468 7395
rect 22502 7392 22514 7395
rect 23014 7392 23020 7404
rect 22502 7364 23020 7392
rect 22502 7361 22514 7364
rect 22456 7355 22514 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 25225 7395 25283 7401
rect 25225 7392 25237 7395
rect 24084 7364 25237 7392
rect 24084 7352 24090 7364
rect 25225 7361 25237 7364
rect 25271 7361 25283 7395
rect 25424 7392 25452 7500
rect 25958 7488 25964 7540
rect 26016 7488 26022 7540
rect 28442 7488 28448 7540
rect 28500 7488 28506 7540
rect 28718 7488 28724 7540
rect 28776 7528 28782 7540
rect 28813 7531 28871 7537
rect 28813 7528 28825 7531
rect 28776 7500 28825 7528
rect 28776 7488 28782 7500
rect 28813 7497 28825 7500
rect 28859 7497 28871 7531
rect 28813 7491 28871 7497
rect 29638 7488 29644 7540
rect 29696 7528 29702 7540
rect 29733 7531 29791 7537
rect 29733 7528 29745 7531
rect 29696 7500 29745 7528
rect 29696 7488 29702 7500
rect 29733 7497 29745 7500
rect 29779 7497 29791 7531
rect 29733 7491 29791 7497
rect 30558 7488 30564 7540
rect 30616 7528 30622 7540
rect 31570 7528 31576 7540
rect 30616 7500 31576 7528
rect 30616 7488 30622 7500
rect 31570 7488 31576 7500
rect 31628 7528 31634 7540
rect 31849 7531 31907 7537
rect 31849 7528 31861 7531
rect 31628 7500 31861 7528
rect 31628 7488 31634 7500
rect 31849 7497 31861 7500
rect 31895 7497 31907 7531
rect 31849 7491 31907 7497
rect 32398 7488 32404 7540
rect 32456 7488 32462 7540
rect 34238 7488 34244 7540
rect 34296 7488 34302 7540
rect 34514 7488 34520 7540
rect 34572 7528 34578 7540
rect 34701 7531 34759 7537
rect 34701 7528 34713 7531
rect 34572 7500 34713 7528
rect 34572 7488 34578 7500
rect 34701 7497 34713 7500
rect 34747 7497 34759 7531
rect 34701 7491 34759 7497
rect 35250 7488 35256 7540
rect 35308 7528 35314 7540
rect 35529 7531 35587 7537
rect 35529 7528 35541 7531
rect 35308 7500 35541 7528
rect 35308 7488 35314 7500
rect 35529 7497 35541 7500
rect 35575 7497 35587 7531
rect 35529 7491 35587 7497
rect 35802 7488 35808 7540
rect 35860 7528 35866 7540
rect 36446 7528 36452 7540
rect 35860 7500 36452 7528
rect 35860 7488 35866 7500
rect 36446 7488 36452 7500
rect 36504 7528 36510 7540
rect 36814 7528 36820 7540
rect 36504 7500 36820 7528
rect 36504 7488 36510 7500
rect 36814 7488 36820 7500
rect 36872 7488 36878 7540
rect 38378 7488 38384 7540
rect 38436 7488 38442 7540
rect 38470 7488 38476 7540
rect 38528 7528 38534 7540
rect 40865 7531 40923 7537
rect 40865 7528 40877 7531
rect 38528 7500 40877 7528
rect 38528 7488 38534 7500
rect 40865 7497 40877 7500
rect 40911 7497 40923 7531
rect 40865 7491 40923 7497
rect 41049 7531 41107 7537
rect 41049 7497 41061 7531
rect 41095 7528 41107 7531
rect 41414 7528 41420 7540
rect 41095 7500 41420 7528
rect 41095 7497 41107 7500
rect 41049 7491 41107 7497
rect 25492 7463 25550 7469
rect 25492 7429 25504 7463
rect 25538 7460 25550 7463
rect 25976 7460 26004 7488
rect 37734 7460 37740 7472
rect 25538 7432 26004 7460
rect 26068 7432 37740 7460
rect 25538 7429 25550 7432
rect 25492 7423 25550 7429
rect 26068 7392 26096 7432
rect 37734 7420 37740 7432
rect 37792 7420 37798 7472
rect 38102 7420 38108 7472
rect 38160 7460 38166 7472
rect 40678 7460 40684 7472
rect 38160 7432 40684 7460
rect 38160 7420 38166 7432
rect 40678 7420 40684 7432
rect 40736 7420 40742 7472
rect 25424 7364 26096 7392
rect 25225 7355 25283 7361
rect 28810 7352 28816 7404
rect 28868 7392 28874 7404
rect 28905 7395 28963 7401
rect 28905 7392 28917 7395
rect 28868 7364 28917 7392
rect 28868 7352 28874 7364
rect 28905 7361 28917 7364
rect 28951 7392 28963 7395
rect 28951 7364 29684 7392
rect 28951 7361 28963 7364
rect 28905 7355 28963 7361
rect 13814 7284 13820 7336
rect 13872 7284 13878 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 15102 7324 15108 7336
rect 13964 7296 15108 7324
rect 13964 7284 13970 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 16592 7324 16620 7352
rect 15304 7296 16620 7324
rect 15304 7256 15332 7296
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18288 7296 18889 7324
rect 18288 7284 18294 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 19024 7296 19257 7324
rect 19024 7284 19030 7296
rect 19245 7293 19257 7296
rect 19291 7293 19303 7327
rect 19245 7287 19303 7293
rect 24305 7327 24363 7333
rect 24305 7293 24317 7327
rect 24351 7293 24363 7327
rect 24305 7287 24363 7293
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7293 27583 7327
rect 27525 7287 27583 7293
rect 28353 7327 28411 7333
rect 28353 7293 28365 7327
rect 28399 7324 28411 7327
rect 28997 7327 29055 7333
rect 28997 7324 29009 7327
rect 28399 7296 29009 7324
rect 28399 7293 28411 7296
rect 28353 7287 28411 7293
rect 28997 7293 29009 7296
rect 29043 7324 29055 7327
rect 29656 7324 29684 7364
rect 29730 7352 29736 7404
rect 29788 7392 29794 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29788 7364 29837 7392
rect 29788 7352 29794 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 29825 7355 29883 7361
rect 30929 7395 30987 7401
rect 30929 7361 30941 7395
rect 30975 7361 30987 7395
rect 32677 7395 32735 7401
rect 32677 7392 32689 7395
rect 30929 7355 30987 7361
rect 31128 7364 32689 7392
rect 30944 7324 30972 7355
rect 31128 7336 31156 7364
rect 32677 7361 32689 7364
rect 32723 7392 32735 7395
rect 33965 7395 34023 7401
rect 33965 7392 33977 7395
rect 32723 7364 33977 7392
rect 32723 7361 32735 7364
rect 32677 7355 32735 7361
rect 33965 7361 33977 7364
rect 34011 7361 34023 7395
rect 33965 7355 34023 7361
rect 34333 7395 34391 7401
rect 34333 7361 34345 7395
rect 34379 7361 34391 7395
rect 34333 7355 34391 7361
rect 29043 7296 29097 7324
rect 29656 7296 30972 7324
rect 29043 7293 29055 7296
rect 28997 7287 29055 7293
rect 23569 7259 23627 7265
rect 13464 7228 15332 7256
rect 16868 7228 22048 7256
rect 13357 7219 13415 7225
rect 3752 7160 4568 7188
rect 7009 7191 7067 7197
rect 3752 7148 3758 7160
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7374 7188 7380 7200
rect 7055 7160 7380 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7374 7148 7380 7160
rect 7432 7188 7438 7200
rect 7650 7188 7656 7200
rect 7432 7160 7656 7188
rect 7432 7148 7438 7160
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8478 7188 8484 7200
rect 8343 7160 8484 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 8662 7188 8668 7200
rect 8536 7160 8668 7188
rect 8536 7148 8542 7160
rect 8662 7148 8668 7160
rect 8720 7188 8726 7200
rect 8987 7191 9045 7197
rect 8987 7188 8999 7191
rect 8720 7160 8999 7188
rect 8720 7148 8726 7160
rect 8987 7157 8999 7160
rect 9033 7157 9045 7191
rect 8987 7151 9045 7157
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 12434 7188 12440 7200
rect 11379 7160 12440 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14148 7160 14933 7188
rect 14148 7148 14154 7160
rect 14921 7157 14933 7160
rect 14967 7188 14979 7191
rect 15194 7188 15200 7200
rect 14967 7160 15200 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15194 7148 15200 7160
rect 15252 7188 15258 7200
rect 16022 7188 16028 7200
rect 15252 7160 16028 7188
rect 15252 7148 15258 7160
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16868 7197 16896 7228
rect 22020 7200 22048 7228
rect 23569 7225 23581 7259
rect 23615 7256 23627 7259
rect 24320 7256 24348 7287
rect 24854 7256 24860 7268
rect 23615 7228 24860 7256
rect 23615 7225 23627 7228
rect 23569 7219 23627 7225
rect 24854 7216 24860 7228
rect 24912 7216 24918 7268
rect 26602 7216 26608 7268
rect 26660 7256 26666 7268
rect 27540 7256 27568 7287
rect 26660 7228 27568 7256
rect 29012 7256 29040 7287
rect 30190 7256 30196 7268
rect 29012 7228 30196 7256
rect 26660 7216 26666 7228
rect 30190 7216 30196 7228
rect 30248 7216 30254 7268
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16724 7160 16865 7188
rect 16724 7148 16730 7160
rect 16853 7157 16865 7160
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18141 7191 18199 7197
rect 18141 7188 18153 7191
rect 18012 7160 18153 7188
rect 18012 7148 18018 7160
rect 18141 7157 18153 7160
rect 18187 7157 18199 7191
rect 18141 7151 18199 7157
rect 18322 7148 18328 7200
rect 18380 7148 18386 7200
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 21266 7188 21272 7200
rect 19935 7160 21272 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21542 7148 21548 7200
rect 21600 7148 21606 7200
rect 22002 7148 22008 7200
rect 22060 7148 22066 7200
rect 23750 7148 23756 7200
rect 23808 7148 23814 7200
rect 26786 7148 26792 7200
rect 26844 7188 26850 7200
rect 26973 7191 27031 7197
rect 26973 7188 26985 7191
rect 26844 7160 26985 7188
rect 26844 7148 26850 7160
rect 26973 7157 26985 7160
rect 27019 7157 27031 7191
rect 26973 7151 27031 7157
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 27893 7191 27951 7197
rect 27893 7188 27905 7191
rect 27672 7160 27905 7188
rect 27672 7148 27678 7160
rect 27893 7157 27905 7160
rect 27939 7188 27951 7191
rect 29454 7188 29460 7200
rect 27939 7160 29460 7188
rect 27939 7157 27951 7160
rect 27893 7151 27951 7157
rect 29454 7148 29460 7160
rect 29512 7188 29518 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29512 7160 29561 7188
rect 29512 7148 29518 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 30374 7148 30380 7200
rect 30432 7148 30438 7200
rect 30558 7148 30564 7200
rect 30616 7148 30622 7200
rect 30944 7188 30972 7296
rect 31021 7327 31079 7333
rect 31021 7293 31033 7327
rect 31067 7293 31079 7327
rect 31021 7287 31079 7293
rect 31036 7256 31064 7287
rect 31110 7284 31116 7336
rect 31168 7284 31174 7336
rect 33410 7284 33416 7336
rect 33468 7284 33474 7336
rect 34348 7324 34376 7355
rect 34882 7352 34888 7404
rect 34940 7392 34946 7404
rect 35253 7395 35311 7401
rect 35253 7392 35265 7395
rect 34940 7364 35265 7392
rect 34940 7352 34946 7364
rect 35253 7361 35265 7364
rect 35299 7361 35311 7395
rect 35253 7355 35311 7361
rect 35618 7352 35624 7404
rect 35676 7392 35682 7404
rect 35676 7364 36492 7392
rect 35676 7352 35682 7364
rect 35894 7324 35900 7336
rect 34348 7296 35900 7324
rect 35894 7284 35900 7296
rect 35952 7284 35958 7336
rect 36078 7284 36084 7336
rect 36136 7284 36142 7336
rect 36464 7324 36492 7364
rect 36538 7352 36544 7404
rect 36596 7392 36602 7404
rect 37182 7392 37188 7404
rect 36596 7364 37188 7392
rect 36596 7352 36602 7364
rect 37182 7352 37188 7364
rect 37240 7352 37246 7404
rect 37829 7395 37887 7401
rect 37829 7361 37841 7395
rect 37875 7392 37887 7395
rect 37918 7392 37924 7404
rect 37875 7364 37924 7392
rect 37875 7361 37887 7364
rect 37829 7355 37887 7361
rect 37918 7352 37924 7364
rect 37976 7352 37982 7404
rect 38470 7352 38476 7404
rect 38528 7392 38534 7404
rect 39669 7395 39727 7401
rect 39669 7392 39681 7395
rect 38528 7364 39681 7392
rect 38528 7352 38534 7364
rect 39669 7361 39681 7364
rect 39715 7392 39727 7395
rect 40402 7392 40408 7404
rect 39715 7364 40408 7392
rect 39715 7361 39727 7364
rect 39669 7355 39727 7361
rect 40402 7352 40408 7364
rect 40460 7352 40466 7404
rect 36722 7324 36728 7336
rect 36464 7296 36728 7324
rect 36722 7284 36728 7296
rect 36780 7324 36786 7336
rect 37553 7327 37611 7333
rect 37553 7324 37565 7327
rect 36780 7296 37565 7324
rect 36780 7284 36786 7296
rect 37553 7293 37565 7296
rect 37599 7324 37611 7327
rect 38010 7324 38016 7336
rect 37599 7296 38016 7324
rect 37599 7293 37611 7296
rect 37553 7287 37611 7293
rect 38010 7284 38016 7296
rect 38068 7284 38074 7336
rect 38194 7284 38200 7336
rect 38252 7324 38258 7336
rect 38378 7324 38384 7336
rect 38252 7296 38384 7324
rect 38252 7284 38258 7296
rect 38378 7284 38384 7296
rect 38436 7324 38442 7336
rect 40126 7324 40132 7336
rect 38436 7296 40132 7324
rect 38436 7284 38442 7296
rect 40126 7284 40132 7296
rect 40184 7284 40190 7336
rect 40494 7284 40500 7336
rect 40552 7284 40558 7336
rect 40880 7324 40908 7491
rect 41414 7488 41420 7500
rect 41472 7488 41478 7540
rect 41506 7488 41512 7540
rect 41564 7488 41570 7540
rect 42242 7488 42248 7540
rect 42300 7528 42306 7540
rect 42429 7531 42487 7537
rect 42429 7528 42441 7531
rect 42300 7500 42441 7528
rect 42300 7488 42306 7500
rect 42429 7497 42441 7500
rect 42475 7497 42487 7531
rect 42429 7491 42487 7497
rect 43530 7488 43536 7540
rect 43588 7528 43594 7540
rect 44913 7531 44971 7537
rect 44913 7528 44925 7531
rect 43588 7500 44925 7528
rect 43588 7488 43594 7500
rect 44913 7497 44925 7500
rect 44959 7497 44971 7531
rect 44913 7491 44971 7497
rect 46750 7488 46756 7540
rect 46808 7488 46814 7540
rect 47578 7488 47584 7540
rect 47636 7488 47642 7540
rect 48590 7488 48596 7540
rect 48648 7488 48654 7540
rect 49142 7488 49148 7540
rect 49200 7528 49206 7540
rect 49329 7531 49387 7537
rect 49329 7528 49341 7531
rect 49200 7500 49341 7528
rect 49200 7488 49206 7500
rect 49329 7497 49341 7500
rect 49375 7497 49387 7531
rect 49329 7491 49387 7497
rect 51994 7488 52000 7540
rect 52052 7528 52058 7540
rect 53466 7528 53472 7540
rect 52052 7500 53472 7528
rect 52052 7488 52058 7500
rect 53466 7488 53472 7500
rect 53524 7488 53530 7540
rect 54018 7488 54024 7540
rect 54076 7488 54082 7540
rect 54110 7488 54116 7540
rect 54168 7488 54174 7540
rect 56778 7488 56784 7540
rect 56836 7528 56842 7540
rect 57241 7531 57299 7537
rect 57241 7528 57253 7531
rect 56836 7500 57253 7528
rect 56836 7488 56842 7500
rect 57241 7497 57253 7500
rect 57287 7497 57299 7531
rect 57241 7491 57299 7497
rect 57606 7488 57612 7540
rect 57664 7488 57670 7540
rect 57882 7488 57888 7540
rect 57940 7488 57946 7540
rect 41966 7420 41972 7472
rect 42024 7460 42030 7472
rect 42153 7463 42211 7469
rect 42153 7460 42165 7463
rect 42024 7432 42165 7460
rect 42024 7420 42030 7432
rect 42153 7429 42165 7432
rect 42199 7460 42211 7463
rect 43990 7460 43996 7472
rect 42199 7432 43996 7460
rect 42199 7429 42211 7432
rect 42153 7423 42211 7429
rect 43990 7420 43996 7432
rect 44048 7420 44054 7472
rect 44082 7420 44088 7472
rect 44140 7460 44146 7472
rect 52546 7460 52552 7472
rect 44140 7432 52552 7460
rect 44140 7420 44146 7432
rect 52546 7420 52552 7432
rect 52604 7420 52610 7472
rect 53837 7463 53895 7469
rect 53837 7429 53849 7463
rect 53883 7460 53895 7463
rect 54036 7460 54064 7488
rect 55582 7460 55588 7472
rect 53883 7432 55588 7460
rect 53883 7429 53895 7432
rect 53837 7423 53895 7429
rect 55582 7420 55588 7432
rect 55640 7460 55646 7472
rect 55861 7463 55919 7469
rect 55861 7460 55873 7463
rect 55640 7432 55873 7460
rect 55640 7420 55646 7432
rect 55861 7429 55873 7432
rect 55907 7429 55919 7463
rect 58066 7460 58072 7472
rect 55861 7423 55919 7429
rect 56336 7432 58072 7460
rect 41414 7352 41420 7404
rect 41472 7352 41478 7404
rect 42702 7352 42708 7404
rect 42760 7392 42766 7404
rect 42797 7395 42855 7401
rect 42797 7392 42809 7395
rect 42760 7364 42809 7392
rect 42760 7352 42766 7364
rect 42797 7361 42809 7364
rect 42843 7361 42855 7395
rect 42797 7355 42855 7361
rect 42889 7395 42947 7401
rect 42889 7361 42901 7395
rect 42935 7392 42947 7395
rect 43257 7395 43315 7401
rect 43257 7392 43269 7395
rect 42935 7364 43269 7392
rect 42935 7361 42947 7364
rect 42889 7355 42947 7361
rect 43257 7361 43269 7364
rect 43303 7361 43315 7395
rect 44177 7395 44235 7401
rect 44177 7392 44189 7395
rect 43257 7355 43315 7361
rect 43364 7364 44189 7392
rect 41601 7327 41659 7333
rect 41601 7324 41613 7327
rect 40880 7296 41613 7324
rect 41601 7293 41613 7296
rect 41647 7293 41659 7327
rect 41601 7287 41659 7293
rect 41690 7284 41696 7336
rect 41748 7324 41754 7336
rect 42981 7327 43039 7333
rect 42981 7324 42993 7327
rect 41748 7296 42993 7324
rect 41748 7284 41754 7296
rect 42981 7293 42993 7296
rect 43027 7324 43039 7327
rect 43364 7324 43392 7364
rect 44177 7361 44189 7364
rect 44223 7361 44235 7395
rect 44177 7355 44235 7361
rect 43027 7296 43392 7324
rect 43027 7293 43039 7296
rect 42981 7287 43039 7293
rect 43438 7284 43444 7336
rect 43496 7324 43502 7336
rect 43809 7327 43867 7333
rect 43809 7324 43821 7327
rect 43496 7296 43821 7324
rect 43496 7284 43502 7296
rect 43809 7293 43821 7296
rect 43855 7293 43867 7327
rect 44192 7324 44220 7355
rect 45370 7352 45376 7404
rect 45428 7392 45434 7404
rect 46017 7395 46075 7401
rect 46017 7392 46029 7395
rect 45428 7364 46029 7392
rect 45428 7352 45434 7364
rect 46017 7361 46029 7364
rect 46063 7361 46075 7395
rect 46017 7355 46075 7361
rect 48225 7395 48283 7401
rect 48225 7361 48237 7395
rect 48271 7392 48283 7395
rect 48314 7392 48320 7404
rect 48271 7364 48320 7392
rect 48271 7361 48283 7364
rect 48225 7355 48283 7361
rect 48314 7352 48320 7364
rect 48372 7352 48378 7404
rect 48682 7352 48688 7404
rect 48740 7392 48746 7404
rect 49145 7395 49203 7401
rect 49145 7392 49157 7395
rect 48740 7364 49157 7392
rect 48740 7352 48746 7364
rect 49145 7361 49157 7364
rect 49191 7361 49203 7395
rect 49145 7355 49203 7361
rect 49878 7352 49884 7404
rect 49936 7352 49942 7404
rect 49973 7395 50031 7401
rect 49973 7361 49985 7395
rect 50019 7392 50031 7395
rect 50246 7392 50252 7404
rect 50019 7364 50252 7392
rect 50019 7361 50031 7364
rect 49973 7355 50031 7361
rect 50246 7352 50252 7364
rect 50304 7352 50310 7404
rect 51721 7395 51779 7401
rect 51721 7392 51733 7395
rect 51046 7364 51733 7392
rect 48774 7324 48780 7336
rect 44192 7296 48780 7324
rect 43809 7287 43867 7293
rect 48774 7284 48780 7296
rect 48832 7284 48838 7336
rect 49896 7324 49924 7352
rect 51046 7324 51074 7364
rect 51721 7361 51733 7364
rect 51767 7392 51779 7395
rect 52178 7392 52184 7404
rect 51767 7364 52184 7392
rect 51767 7361 51779 7364
rect 51721 7355 51779 7361
rect 52178 7352 52184 7364
rect 52236 7352 52242 7404
rect 54757 7395 54815 7401
rect 54757 7361 54769 7395
rect 54803 7392 54815 7395
rect 55122 7392 55128 7404
rect 54803 7364 55128 7392
rect 54803 7361 54815 7364
rect 54757 7355 54815 7361
rect 55122 7352 55128 7364
rect 55180 7352 55186 7404
rect 56336 7401 56364 7432
rect 58066 7420 58072 7432
rect 58124 7420 58130 7472
rect 56321 7395 56379 7401
rect 56321 7361 56333 7395
rect 56367 7361 56379 7395
rect 56321 7355 56379 7361
rect 57517 7395 57575 7401
rect 57517 7361 57529 7395
rect 57563 7392 57575 7395
rect 57606 7392 57612 7404
rect 57563 7364 57612 7392
rect 57563 7361 57575 7364
rect 57517 7355 57575 7361
rect 57606 7352 57612 7364
rect 57664 7352 57670 7404
rect 49896 7296 51074 7324
rect 52196 7324 52224 7352
rect 55217 7327 55275 7333
rect 55217 7324 55229 7327
rect 52196 7296 55229 7324
rect 55217 7293 55229 7296
rect 55263 7324 55275 7327
rect 55858 7324 55864 7336
rect 55263 7296 55864 7324
rect 55263 7293 55275 7296
rect 55217 7287 55275 7293
rect 55858 7284 55864 7296
rect 55916 7284 55922 7336
rect 56502 7284 56508 7336
rect 56560 7324 56566 7336
rect 58437 7327 58495 7333
rect 58437 7324 58449 7327
rect 56560 7296 58449 7324
rect 56560 7284 56566 7296
rect 58437 7293 58449 7296
rect 58483 7293 58495 7327
rect 58437 7287 58495 7293
rect 32306 7256 32312 7268
rect 31036 7228 32312 7256
rect 32306 7216 32312 7228
rect 32364 7216 32370 7268
rect 32674 7216 32680 7268
rect 32732 7256 32738 7268
rect 39850 7256 39856 7268
rect 32732 7228 39856 7256
rect 32732 7216 32738 7228
rect 39850 7216 39856 7228
rect 39908 7216 39914 7268
rect 44910 7216 44916 7268
rect 44968 7256 44974 7268
rect 56965 7259 57023 7265
rect 44968 7228 51074 7256
rect 44968 7216 44974 7228
rect 32490 7188 32496 7200
rect 30944 7160 32496 7188
rect 32490 7148 32496 7160
rect 32548 7148 32554 7200
rect 33410 7148 33416 7200
rect 33468 7188 33474 7200
rect 35618 7188 35624 7200
rect 33468 7160 35624 7188
rect 33468 7148 33474 7160
rect 35618 7148 35624 7160
rect 35676 7148 35682 7200
rect 36446 7148 36452 7200
rect 36504 7148 36510 7200
rect 38470 7148 38476 7200
rect 38528 7188 38534 7200
rect 38657 7191 38715 7197
rect 38657 7188 38669 7191
rect 38528 7160 38669 7188
rect 38528 7148 38534 7160
rect 38657 7157 38669 7160
rect 38703 7157 38715 7191
rect 38657 7151 38715 7157
rect 38746 7148 38752 7200
rect 38804 7188 38810 7200
rect 39022 7188 39028 7200
rect 38804 7160 39028 7188
rect 38804 7148 38810 7160
rect 39022 7148 39028 7160
rect 39080 7148 39086 7200
rect 44637 7191 44695 7197
rect 44637 7157 44649 7191
rect 44683 7188 44695 7191
rect 44818 7188 44824 7200
rect 44683 7160 44824 7188
rect 44683 7157 44695 7160
rect 44637 7151 44695 7157
rect 44818 7148 44824 7160
rect 44876 7148 44882 7200
rect 45186 7148 45192 7200
rect 45244 7188 45250 7200
rect 45281 7191 45339 7197
rect 45281 7188 45293 7191
rect 45244 7160 45293 7188
rect 45244 7148 45250 7160
rect 45281 7157 45293 7160
rect 45327 7188 45339 7191
rect 45649 7191 45707 7197
rect 45649 7188 45661 7191
rect 45327 7160 45661 7188
rect 45327 7157 45339 7160
rect 45281 7151 45339 7157
rect 45649 7157 45661 7160
rect 45695 7157 45707 7191
rect 45649 7151 45707 7157
rect 46474 7148 46480 7200
rect 46532 7188 46538 7200
rect 47118 7188 47124 7200
rect 46532 7160 47124 7188
rect 46532 7148 46538 7160
rect 47118 7148 47124 7160
rect 47176 7148 47182 7200
rect 51046 7188 51074 7228
rect 51552 7228 54800 7256
rect 51552 7188 51580 7228
rect 54772 7200 54800 7228
rect 56965 7225 56977 7259
rect 57011 7256 57023 7259
rect 58250 7256 58256 7268
rect 57011 7228 58256 7256
rect 57011 7225 57023 7228
rect 56965 7219 57023 7225
rect 58250 7216 58256 7228
rect 58308 7216 58314 7268
rect 51046 7160 51580 7188
rect 51994 7148 52000 7200
rect 52052 7148 52058 7200
rect 52549 7191 52607 7197
rect 52549 7157 52561 7191
rect 52595 7188 52607 7191
rect 52638 7188 52644 7200
rect 52595 7160 52644 7188
rect 52595 7157 52607 7160
rect 52549 7151 52607 7157
rect 52638 7148 52644 7160
rect 52696 7148 52702 7200
rect 52914 7148 52920 7200
rect 52972 7148 52978 7200
rect 54754 7148 54760 7200
rect 54812 7148 54818 7200
rect 55490 7148 55496 7200
rect 55548 7148 55554 7200
rect 1104 7098 58880 7120
rect 1104 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 22616 7098
rect 22668 7046 22680 7098
rect 22732 7046 22744 7098
rect 22796 7046 22808 7098
rect 22860 7046 22872 7098
rect 22924 7046 37060 7098
rect 37112 7046 37124 7098
rect 37176 7046 37188 7098
rect 37240 7046 37252 7098
rect 37304 7046 37316 7098
rect 37368 7046 51504 7098
rect 51556 7046 51568 7098
rect 51620 7046 51632 7098
rect 51684 7046 51696 7098
rect 51748 7046 51760 7098
rect 51812 7046 58880 7098
rect 1104 7024 58880 7046
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 4525 6987 4583 6993
rect 4525 6984 4537 6987
rect 3476 6956 4537 6984
rect 3476 6944 3482 6956
rect 4525 6953 4537 6956
rect 4571 6953 4583 6987
rect 4525 6947 4583 6953
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12308 6956 13768 6984
rect 12308 6944 12314 6956
rect 5074 6916 5080 6928
rect 5000 6888 5080 6916
rect 3326 6808 3332 6860
rect 3384 6808 3390 6860
rect 4338 6808 4344 6860
rect 4396 6808 4402 6860
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 5000 6789 5028 6888
rect 5074 6876 5080 6888
rect 5132 6916 5138 6928
rect 5445 6919 5503 6925
rect 5445 6916 5457 6919
rect 5132 6888 5457 6916
rect 5132 6876 5138 6888
rect 5445 6885 5457 6888
rect 5491 6885 5503 6919
rect 5445 6879 5503 6885
rect 12342 6876 12348 6928
rect 12400 6876 12406 6928
rect 13740 6916 13768 6956
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13872 6956 14105 6984
rect 13872 6944 13878 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 23477 6987 23535 6993
rect 20496 6956 23336 6984
rect 20496 6944 20502 6956
rect 13906 6916 13912 6928
rect 13740 6888 13912 6916
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 21358 6916 21364 6928
rect 19812 6888 20024 6916
rect 21319 6888 21364 6916
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6454 6848 6460 6860
rect 5675 6820 6460 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6454 6808 6460 6820
rect 6512 6848 6518 6860
rect 7098 6848 7104 6860
rect 6512 6820 7104 6848
rect 6512 6808 6518 6820
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7558 6848 7564 6860
rect 7423 6820 7564 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7800 6820 7941 6848
rect 7800 6808 7806 6820
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 6871 6752 7512 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 3084 6715 3142 6721
rect 3084 6681 3096 6715
rect 3130 6712 3142 6715
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3130 6684 3801 6712
rect 3130 6681 3142 6684
rect 3084 6675 3142 6681
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 5000 6712 5028 6743
rect 4120 6684 5028 6712
rect 5169 6715 5227 6721
rect 4120 6672 4126 6684
rect 5169 6681 5181 6715
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 3694 6644 3700 6656
rect 1995 6616 3700 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4890 6644 4896 6656
rect 4028 6616 4896 6644
rect 4028 6604 4034 6616
rect 4890 6604 4896 6616
rect 4948 6644 4954 6656
rect 5184 6644 5212 6675
rect 4948 6616 5212 6644
rect 5997 6647 6055 6653
rect 4948 6604 4954 6616
rect 5997 6613 6009 6647
rect 6043 6644 6055 6647
rect 6362 6644 6368 6656
rect 6043 6616 6368 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 6822 6644 6828 6656
rect 6687 6616 6828 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 6822 6604 6828 6616
rect 6880 6644 6886 6656
rect 7098 6644 7104 6656
rect 6880 6616 7104 6644
rect 6880 6604 6886 6616
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7484 6653 7512 6752
rect 8128 6712 8156 6811
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 12360 6848 12388 6876
rect 8628 6820 10364 6848
rect 8628 6808 8634 6820
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 9122 6780 9128 6792
rect 8260 6752 9128 6780
rect 8260 6740 8266 6752
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9180 6752 9413 6780
rect 9180 6740 9186 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 10336 6789 10364 6820
rect 11348 6820 12388 6848
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 11348 6780 11376 6820
rect 12360 6789 12388 6820
rect 13372 6820 16988 6848
rect 10367 6752 11376 6780
rect 12345 6783 12403 6789
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 12345 6749 12357 6783
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12601 6783 12659 6789
rect 12601 6780 12613 6783
rect 12492 6752 12613 6780
rect 12492 6740 12498 6752
rect 12601 6749 12613 6752
rect 12647 6749 12659 6783
rect 12601 6743 12659 6749
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 8128 6684 8585 6712
rect 8573 6681 8585 6684
rect 8619 6712 8631 6715
rect 9030 6712 9036 6724
rect 8619 6684 9036 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 9030 6672 9036 6684
rect 9088 6712 9094 6724
rect 10588 6715 10646 6721
rect 9088 6684 10548 6712
rect 9088 6672 9094 6684
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 7837 6647 7895 6653
rect 7837 6613 7849 6647
rect 7883 6644 7895 6647
rect 9122 6644 9128 6656
rect 7883 6616 9128 6644
rect 7883 6613 7895 6616
rect 7837 6607 7895 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 10226 6604 10232 6656
rect 10284 6604 10290 6656
rect 10520 6644 10548 6684
rect 10588 6681 10600 6715
rect 10634 6712 10646 6715
rect 11054 6712 11060 6724
rect 10634 6684 11060 6712
rect 10634 6681 10646 6684
rect 10588 6675 10646 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 12250 6712 12256 6724
rect 11624 6684 12256 6712
rect 11624 6644 11652 6684
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 13372 6712 13400 6820
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 12406 6684 13400 6712
rect 10520 6616 11652 6644
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12158 6644 12164 6656
rect 11848 6616 12164 6644
rect 11848 6604 11854 6616
rect 12158 6604 12164 6616
rect 12216 6644 12222 6656
rect 12406 6644 12434 6684
rect 12216 6616 12434 6644
rect 13725 6647 13783 6653
rect 12216 6604 12222 6616
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 14274 6644 14280 6656
rect 13771 6616 14280 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14274 6604 14280 6616
rect 14332 6644 14338 6656
rect 14660 6644 14688 6743
rect 14734 6740 14740 6792
rect 14792 6780 14798 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 14792 6752 15393 6780
rect 14792 6740 14798 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16224 6712 16252 6743
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16724 6752 16865 6780
rect 16724 6740 16730 6752
rect 16853 6749 16865 6752
rect 16899 6749 16911 6783
rect 16960 6780 16988 6820
rect 17954 6808 17960 6860
rect 18012 6848 18018 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18012 6820 18889 6848
rect 18012 6808 18018 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 19242 6808 19248 6860
rect 19300 6808 19306 6860
rect 19610 6848 19616 6860
rect 19352 6820 19616 6848
rect 17972 6780 18000 6808
rect 19352 6780 19380 6820
rect 19610 6808 19616 6820
rect 19668 6848 19674 6860
rect 19812 6848 19840 6888
rect 19668 6820 19840 6848
rect 19668 6808 19674 6820
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 19996 6848 20024 6888
rect 21358 6876 21364 6888
rect 21416 6876 21422 6928
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 19996 6820 20177 6848
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20254 6808 20260 6860
rect 20312 6857 20318 6860
rect 20312 6851 20340 6857
rect 20328 6817 20340 6851
rect 21376 6848 21404 6876
rect 22005 6851 22063 6857
rect 22005 6848 22017 6851
rect 21376 6820 22017 6848
rect 20312 6811 20340 6817
rect 22005 6817 22017 6820
rect 22051 6817 22063 6851
rect 23308 6848 23336 6956
rect 23477 6953 23489 6987
rect 23523 6984 23535 6987
rect 23566 6984 23572 6996
rect 23523 6956 23572 6984
rect 23523 6953 23535 6956
rect 23477 6947 23535 6953
rect 23566 6944 23572 6956
rect 23624 6944 23630 6996
rect 24670 6944 24676 6996
rect 24728 6984 24734 6996
rect 24728 6956 25636 6984
rect 24728 6944 24734 6956
rect 23658 6848 23664 6860
rect 23308 6820 23664 6848
rect 22005 6811 22063 6817
rect 20312 6808 20318 6811
rect 23658 6808 23664 6820
rect 23716 6808 23722 6860
rect 23750 6808 23756 6860
rect 23808 6848 23814 6860
rect 23937 6851 23995 6857
rect 23937 6848 23949 6851
rect 23808 6820 23949 6848
rect 23808 6808 23814 6820
rect 23937 6817 23949 6820
rect 23983 6817 23995 6851
rect 23937 6811 23995 6817
rect 24121 6851 24179 6857
rect 24121 6817 24133 6851
rect 24167 6848 24179 6851
rect 24302 6848 24308 6860
rect 24167 6820 24308 6848
rect 24167 6817 24179 6820
rect 24121 6811 24179 6817
rect 16960 6752 18000 6780
rect 18248 6752 19380 6780
rect 19429 6783 19487 6789
rect 16853 6743 16911 6749
rect 17120 6715 17178 6721
rect 16224 6684 17080 6712
rect 14332 6616 14688 6644
rect 14332 6604 14338 6616
rect 14826 6604 14832 6656
rect 14884 6604 14890 6656
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 15930 6644 15936 6656
rect 15887 6616 15936 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16758 6604 16764 6656
rect 16816 6604 16822 6656
rect 17052 6644 17080 6684
rect 17120 6681 17132 6715
rect 17166 6712 17178 6715
rect 17770 6712 17776 6724
rect 17166 6684 17776 6712
rect 17166 6681 17178 6684
rect 17120 6675 17178 6681
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 17310 6644 17316 6656
rect 17052 6616 17316 6644
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 18248 6653 18276 6752
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 18693 6715 18751 6721
rect 18693 6681 18705 6715
rect 18739 6712 18751 6715
rect 19334 6712 19340 6724
rect 18739 6684 19340 6712
rect 18739 6681 18751 6684
rect 18693 6675 18751 6681
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 18322 6604 18328 6656
rect 18380 6604 18386 6656
rect 18782 6604 18788 6656
rect 18840 6604 18846 6656
rect 19444 6644 19472 6743
rect 20438 6740 20444 6792
rect 20496 6740 20502 6792
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 24136 6780 24164 6811
rect 24302 6808 24308 6820
rect 24360 6808 24366 6860
rect 24854 6808 24860 6860
rect 24912 6848 24918 6860
rect 25608 6857 25636 6956
rect 25774 6944 25780 6996
rect 25832 6944 25838 6996
rect 26329 6987 26387 6993
rect 26329 6953 26341 6987
rect 26375 6984 26387 6987
rect 26510 6984 26516 6996
rect 26375 6956 26516 6984
rect 26375 6953 26387 6956
rect 26329 6947 26387 6953
rect 26510 6944 26516 6956
rect 26568 6944 26574 6996
rect 30374 6944 30380 6996
rect 30432 6984 30438 6996
rect 31110 6984 31116 6996
rect 30432 6956 31116 6984
rect 30432 6944 30438 6956
rect 31110 6944 31116 6956
rect 31168 6944 31174 6996
rect 41414 6984 41420 6996
rect 36832 6956 38654 6984
rect 25792 6916 25820 6944
rect 36832 6928 36860 6956
rect 25792 6888 26924 6916
rect 25317 6851 25375 6857
rect 25317 6848 25329 6851
rect 24912 6820 25329 6848
rect 24912 6808 24918 6820
rect 25317 6817 25329 6820
rect 25363 6817 25375 6851
rect 25317 6811 25375 6817
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6848 25651 6851
rect 25682 6848 25688 6860
rect 25639 6820 25688 6848
rect 25639 6817 25651 6820
rect 25593 6811 25651 6817
rect 25682 6808 25688 6820
rect 25740 6808 25746 6860
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26602 6848 26608 6860
rect 26283 6820 26608 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 26786 6808 26792 6860
rect 26844 6808 26850 6860
rect 26896 6857 26924 6888
rect 30190 6876 30196 6928
rect 30248 6876 30254 6928
rect 34974 6876 34980 6928
rect 35032 6916 35038 6928
rect 35710 6916 35716 6928
rect 35032 6888 35716 6916
rect 35032 6876 35038 6888
rect 35710 6876 35716 6888
rect 35768 6876 35774 6928
rect 35894 6876 35900 6928
rect 35952 6916 35958 6928
rect 36354 6916 36360 6928
rect 35952 6888 36360 6916
rect 35952 6876 35958 6888
rect 36354 6876 36360 6888
rect 36412 6876 36418 6928
rect 36814 6876 36820 6928
rect 36872 6876 36878 6928
rect 36909 6919 36967 6925
rect 36909 6885 36921 6919
rect 36955 6916 36967 6919
rect 37182 6916 37188 6928
rect 36955 6888 37188 6916
rect 36955 6885 36967 6888
rect 36909 6879 36967 6885
rect 37182 6876 37188 6888
rect 37240 6876 37246 6928
rect 26881 6851 26939 6857
rect 26881 6817 26893 6851
rect 26927 6817 26939 6851
rect 26881 6811 26939 6817
rect 27798 6808 27804 6860
rect 27856 6808 27862 6860
rect 28994 6808 29000 6860
rect 29052 6848 29058 6860
rect 30009 6851 30067 6857
rect 30009 6848 30021 6851
rect 29052 6820 30021 6848
rect 29052 6808 29058 6820
rect 30009 6817 30021 6820
rect 30055 6817 30067 6851
rect 30009 6811 30067 6817
rect 30101 6851 30159 6857
rect 30101 6817 30113 6851
rect 30147 6848 30159 6851
rect 30208 6848 30236 6876
rect 30147 6820 30236 6848
rect 30147 6817 30159 6820
rect 30101 6811 30159 6817
rect 30466 6808 30472 6860
rect 30524 6808 30530 6860
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 31021 6851 31079 6857
rect 31021 6848 31033 6851
rect 30616 6820 31033 6848
rect 30616 6808 30622 6820
rect 31021 6817 31033 6820
rect 31067 6817 31079 6851
rect 33873 6851 33931 6857
rect 33873 6848 33885 6851
rect 31021 6811 31079 6817
rect 33428 6820 33885 6848
rect 21968 6752 24164 6780
rect 21968 6740 21974 6752
rect 25038 6740 25044 6792
rect 25096 6740 25102 6792
rect 25130 6740 25136 6792
rect 25188 6789 25194 6792
rect 25188 6783 25237 6789
rect 25188 6749 25191 6783
rect 25225 6749 25237 6783
rect 25188 6743 25237 6749
rect 25188 6740 25194 6743
rect 26050 6740 26056 6792
rect 26108 6780 26114 6792
rect 28537 6783 28595 6789
rect 28537 6780 28549 6783
rect 26108 6752 28549 6780
rect 26108 6740 26114 6752
rect 28537 6749 28549 6752
rect 28583 6749 28595 6783
rect 28537 6743 28595 6749
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6780 29423 6783
rect 31757 6783 31815 6789
rect 29411 6752 29592 6780
rect 29411 6749 29423 6752
rect 29365 6743 29423 6749
rect 22272 6715 22330 6721
rect 22272 6681 22284 6715
rect 22318 6712 22330 6715
rect 22462 6712 22468 6724
rect 22318 6684 22468 6712
rect 22318 6681 22330 6684
rect 22272 6675 22330 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 23400 6684 24532 6712
rect 19702 6644 19708 6656
rect 19444 6616 19708 6644
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 23400 6653 23428 6684
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20956 6616 21097 6644
rect 20956 6604 20962 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 23385 6647 23443 6653
rect 23385 6613 23397 6647
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 23845 6647 23903 6653
rect 23845 6613 23857 6647
rect 23891 6644 23903 6647
rect 23934 6644 23940 6656
rect 23891 6616 23940 6644
rect 23891 6613 23903 6616
rect 23845 6607 23903 6613
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 24394 6604 24400 6656
rect 24452 6604 24458 6656
rect 24504 6644 24532 6684
rect 26694 6672 26700 6724
rect 26752 6712 26758 6724
rect 27525 6715 27583 6721
rect 26752 6684 27292 6712
rect 26752 6672 26758 6684
rect 25130 6644 25136 6656
rect 24504 6616 25136 6644
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 27154 6604 27160 6656
rect 27212 6604 27218 6656
rect 27264 6644 27292 6684
rect 27525 6681 27537 6715
rect 27571 6712 27583 6715
rect 27985 6715 28043 6721
rect 27985 6712 27997 6715
rect 27571 6684 27997 6712
rect 27571 6681 27583 6684
rect 27525 6675 27583 6681
rect 27985 6681 27997 6684
rect 28031 6681 28043 6715
rect 27985 6675 28043 6681
rect 27617 6647 27675 6653
rect 27617 6644 27629 6647
rect 27264 6616 27629 6644
rect 27617 6613 27629 6616
rect 27663 6613 27675 6647
rect 27617 6607 27675 6613
rect 28721 6647 28779 6653
rect 28721 6613 28733 6647
rect 28767 6644 28779 6647
rect 28810 6644 28816 6656
rect 28767 6616 28816 6644
rect 28767 6613 28779 6616
rect 28721 6607 28779 6613
rect 28810 6604 28816 6616
rect 28868 6604 28874 6656
rect 29564 6653 29592 6752
rect 31757 6749 31769 6783
rect 31803 6749 31815 6783
rect 31757 6743 31815 6749
rect 29917 6715 29975 6721
rect 29917 6681 29929 6715
rect 29963 6712 29975 6715
rect 31205 6715 31263 6721
rect 31205 6712 31217 6715
rect 29963 6684 31217 6712
rect 29963 6681 29975 6684
rect 29917 6675 29975 6681
rect 31205 6681 31217 6684
rect 31251 6681 31263 6715
rect 31205 6675 31263 6681
rect 31772 6656 31800 6743
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 33428 6780 33456 6820
rect 33873 6817 33885 6820
rect 33919 6817 33931 6851
rect 33873 6811 33931 6817
rect 35618 6808 35624 6860
rect 35676 6848 35682 6860
rect 35676 6820 36124 6848
rect 35676 6808 35682 6820
rect 32548 6752 33456 6780
rect 33505 6783 33563 6789
rect 32548 6740 32554 6752
rect 33505 6749 33517 6783
rect 33551 6780 33563 6783
rect 33594 6780 33600 6792
rect 33551 6752 33600 6780
rect 33551 6749 33563 6752
rect 33505 6743 33563 6749
rect 33594 6740 33600 6752
rect 33652 6780 33658 6792
rect 33652 6752 34284 6780
rect 33652 6740 33658 6752
rect 33260 6715 33318 6721
rect 33260 6681 33272 6715
rect 33306 6712 33318 6715
rect 33410 6712 33416 6724
rect 33306 6684 33416 6712
rect 33306 6681 33318 6684
rect 33260 6675 33318 6681
rect 33410 6672 33416 6684
rect 33468 6672 33474 6724
rect 33686 6672 33692 6724
rect 33744 6672 33750 6724
rect 34256 6721 34284 6752
rect 35986 6740 35992 6792
rect 36044 6740 36050 6792
rect 36096 6780 36124 6820
rect 36262 6808 36268 6860
rect 36320 6808 36326 6860
rect 37553 6851 37611 6857
rect 37553 6848 37565 6851
rect 36372 6820 37565 6848
rect 36372 6780 36400 6820
rect 37553 6817 37565 6820
rect 37599 6817 37611 6851
rect 37553 6811 37611 6817
rect 36096 6752 36400 6780
rect 36449 6783 36507 6789
rect 36449 6749 36461 6783
rect 36495 6780 36507 6783
rect 37001 6783 37059 6789
rect 37001 6780 37013 6783
rect 36495 6752 37013 6780
rect 36495 6749 36507 6752
rect 36449 6743 36507 6749
rect 37001 6749 37013 6752
rect 37047 6749 37059 6783
rect 38626 6780 38654 6956
rect 41386 6944 41420 6984
rect 41472 6984 41478 6996
rect 42702 6984 42708 6996
rect 41472 6956 42708 6984
rect 41472 6944 41478 6956
rect 42702 6944 42708 6956
rect 42760 6944 42766 6996
rect 45462 6944 45468 6996
rect 45520 6944 45526 6996
rect 54386 6984 54392 6996
rect 52472 6956 54392 6984
rect 41386 6916 41414 6944
rect 41248 6888 41414 6916
rect 40402 6808 40408 6860
rect 40460 6808 40466 6860
rect 41248 6848 41276 6888
rect 43990 6876 43996 6928
rect 44048 6916 44054 6928
rect 44361 6919 44419 6925
rect 44361 6916 44373 6919
rect 44048 6888 44373 6916
rect 44048 6876 44054 6888
rect 44361 6885 44373 6888
rect 44407 6916 44419 6919
rect 45186 6916 45192 6928
rect 44407 6888 45192 6916
rect 44407 6885 44419 6888
rect 44361 6879 44419 6885
rect 45186 6876 45192 6888
rect 45244 6916 45250 6928
rect 45281 6919 45339 6925
rect 45281 6916 45293 6919
rect 45244 6888 45293 6916
rect 45244 6876 45250 6888
rect 45281 6885 45293 6888
rect 45327 6916 45339 6919
rect 45327 6888 48544 6916
rect 45327 6885 45339 6888
rect 45281 6879 45339 6885
rect 48516 6860 48544 6888
rect 52472 6860 52500 6956
rect 54386 6944 54392 6956
rect 54444 6944 54450 6996
rect 55582 6944 55588 6996
rect 55640 6944 55646 6996
rect 53190 6876 53196 6928
rect 53248 6916 53254 6928
rect 53469 6919 53527 6925
rect 53469 6916 53481 6919
rect 53248 6888 53481 6916
rect 53248 6876 53254 6888
rect 53469 6885 53481 6888
rect 53515 6885 53527 6919
rect 56594 6916 56600 6928
rect 53469 6879 53527 6885
rect 56244 6888 56600 6916
rect 42199 6851 42257 6857
rect 42199 6848 42211 6851
rect 40604 6820 41276 6848
rect 41386 6820 42211 6848
rect 39669 6783 39727 6789
rect 38626 6752 38792 6780
rect 37001 6743 37059 6749
rect 34241 6715 34299 6721
rect 34241 6681 34253 6715
rect 34287 6712 34299 6715
rect 35250 6712 35256 6724
rect 34287 6684 35256 6712
rect 34287 6681 34299 6684
rect 34241 6675 34299 6681
rect 35250 6672 35256 6684
rect 35308 6712 35314 6724
rect 35345 6715 35403 6721
rect 35345 6712 35357 6715
rect 35308 6684 35357 6712
rect 35308 6672 35314 6684
rect 35345 6681 35357 6684
rect 35391 6712 35403 6715
rect 37550 6712 37556 6724
rect 35391 6684 37556 6712
rect 35391 6681 35403 6684
rect 35345 6675 35403 6681
rect 37550 6672 37556 6684
rect 37608 6712 37614 6724
rect 37921 6715 37979 6721
rect 37921 6712 37933 6715
rect 37608 6684 37933 6712
rect 37608 6672 37614 6684
rect 37921 6681 37933 6684
rect 37967 6712 37979 6715
rect 38654 6712 38660 6724
rect 37967 6684 38660 6712
rect 37967 6681 37979 6684
rect 37921 6675 37979 6681
rect 38654 6672 38660 6684
rect 38712 6672 38718 6724
rect 29549 6647 29607 6653
rect 29549 6613 29561 6647
rect 29595 6613 29607 6647
rect 29549 6607 29607 6613
rect 31018 6604 31024 6656
rect 31076 6644 31082 6656
rect 31754 6644 31760 6656
rect 31076 6616 31760 6644
rect 31076 6604 31082 6616
rect 31754 6604 31760 6616
rect 31812 6604 31818 6656
rect 32125 6647 32183 6653
rect 32125 6613 32137 6647
rect 32171 6644 32183 6647
rect 33502 6644 33508 6656
rect 32171 6616 33508 6644
rect 32171 6613 32183 6616
rect 32125 6607 32183 6613
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 35434 6604 35440 6656
rect 35492 6604 35498 6656
rect 36078 6604 36084 6656
rect 36136 6644 36142 6656
rect 36541 6647 36599 6653
rect 36541 6644 36553 6647
rect 36136 6616 36553 6644
rect 36136 6604 36142 6616
rect 36541 6613 36553 6616
rect 36587 6644 36599 6647
rect 38286 6644 38292 6656
rect 36587 6616 38292 6644
rect 36587 6613 36599 6616
rect 36541 6607 36599 6613
rect 38286 6604 38292 6616
rect 38344 6604 38350 6656
rect 38381 6647 38439 6653
rect 38381 6613 38393 6647
rect 38427 6644 38439 6647
rect 38562 6644 38568 6656
rect 38427 6616 38568 6644
rect 38427 6613 38439 6616
rect 38381 6607 38439 6613
rect 38562 6604 38568 6616
rect 38620 6644 38626 6656
rect 38764 6644 38792 6752
rect 39669 6749 39681 6783
rect 39715 6780 39727 6783
rect 39715 6752 39896 6780
rect 39715 6749 39727 6752
rect 39669 6743 39727 6749
rect 38620 6616 38792 6644
rect 39025 6647 39083 6653
rect 38620 6604 38626 6616
rect 39025 6613 39037 6647
rect 39071 6644 39083 6647
rect 39114 6644 39120 6656
rect 39071 6616 39120 6644
rect 39071 6613 39083 6616
rect 39025 6607 39083 6613
rect 39114 6604 39120 6616
rect 39172 6604 39178 6656
rect 39868 6653 39896 6752
rect 40126 6740 40132 6792
rect 40184 6780 40190 6792
rect 40313 6783 40371 6789
rect 40313 6780 40325 6783
rect 40184 6752 40325 6780
rect 40184 6740 40190 6752
rect 40313 6749 40325 6752
rect 40359 6780 40371 6783
rect 40604 6780 40632 6820
rect 40359 6752 40632 6780
rect 41233 6783 41291 6789
rect 40359 6749 40371 6752
rect 40313 6743 40371 6749
rect 41233 6749 41245 6783
rect 41279 6780 41291 6783
rect 41386 6780 41414 6820
rect 42199 6817 42211 6820
rect 42245 6817 42257 6851
rect 42199 6811 42257 6817
rect 42337 6851 42395 6857
rect 42337 6817 42349 6851
rect 42383 6848 42395 6851
rect 42518 6848 42524 6860
rect 42383 6820 42524 6848
rect 42383 6817 42395 6820
rect 42337 6811 42395 6817
rect 42518 6808 42524 6820
rect 42576 6808 42582 6860
rect 42610 6808 42616 6860
rect 42668 6808 42674 6860
rect 43254 6808 43260 6860
rect 43312 6808 43318 6860
rect 46658 6808 46664 6860
rect 46716 6848 46722 6860
rect 47397 6851 47455 6857
rect 47397 6848 47409 6851
rect 46716 6820 47409 6848
rect 46716 6808 46722 6820
rect 47397 6817 47409 6820
rect 47443 6848 47455 6851
rect 47854 6848 47860 6860
rect 47443 6820 47860 6848
rect 47443 6817 47455 6820
rect 47397 6811 47455 6817
rect 47854 6808 47860 6820
rect 47912 6808 47918 6860
rect 48498 6808 48504 6860
rect 48556 6808 48562 6860
rect 51813 6851 51871 6857
rect 51813 6848 51825 6851
rect 51276 6820 51825 6848
rect 41279 6752 41414 6780
rect 41279 6749 41291 6752
rect 41233 6743 41291 6749
rect 40221 6715 40279 6721
rect 40221 6681 40233 6715
rect 40267 6712 40279 6715
rect 40681 6715 40739 6721
rect 40681 6712 40693 6715
rect 40267 6684 40693 6712
rect 40267 6681 40279 6684
rect 40221 6675 40279 6681
rect 40681 6681 40693 6684
rect 40727 6681 40739 6715
rect 40681 6675 40739 6681
rect 41248 6656 41276 6743
rect 42058 6740 42064 6792
rect 42116 6740 42122 6792
rect 43070 6740 43076 6792
rect 43128 6740 43134 6792
rect 45646 6740 45652 6792
rect 45704 6780 45710 6792
rect 46293 6783 46351 6789
rect 46293 6780 46305 6783
rect 45704 6752 46305 6780
rect 45704 6740 45710 6752
rect 46293 6749 46305 6752
rect 46339 6749 46351 6783
rect 46293 6743 46351 6749
rect 46750 6740 46756 6792
rect 46808 6780 46814 6792
rect 47029 6783 47087 6789
rect 47029 6780 47041 6783
rect 46808 6752 47041 6780
rect 46808 6740 46814 6752
rect 47029 6749 47041 6752
rect 47075 6780 47087 6783
rect 47302 6780 47308 6792
rect 47075 6752 47308 6780
rect 47075 6749 47087 6752
rect 47029 6743 47087 6749
rect 47302 6740 47308 6752
rect 47360 6740 47366 6792
rect 51276 6780 51304 6820
rect 51813 6817 51825 6820
rect 51859 6848 51871 6851
rect 52454 6848 52460 6860
rect 51859 6820 52460 6848
rect 51859 6817 51871 6820
rect 51813 6811 51871 6817
rect 52454 6808 52460 6820
rect 52512 6808 52518 6860
rect 52638 6808 52644 6860
rect 52696 6848 52702 6860
rect 52733 6851 52791 6857
rect 52733 6848 52745 6851
rect 52696 6820 52745 6848
rect 52696 6808 52702 6820
rect 52733 6817 52745 6820
rect 52779 6817 52791 6851
rect 54205 6851 54263 6857
rect 54205 6848 54217 6851
rect 52733 6811 52791 6817
rect 53024 6820 54217 6848
rect 47412 6752 51304 6780
rect 45557 6715 45615 6721
rect 45557 6681 45569 6715
rect 45603 6712 45615 6715
rect 45830 6712 45836 6724
rect 45603 6684 45836 6712
rect 45603 6681 45615 6684
rect 45557 6675 45615 6681
rect 45830 6672 45836 6684
rect 45888 6672 45894 6724
rect 46474 6672 46480 6724
rect 46532 6712 46538 6724
rect 46658 6712 46664 6724
rect 46532 6684 46664 6712
rect 46532 6672 46538 6684
rect 46658 6672 46664 6684
rect 46716 6712 46722 6724
rect 47412 6712 47440 6752
rect 51902 6740 51908 6792
rect 51960 6740 51966 6792
rect 53024 6789 53052 6820
rect 54205 6817 54217 6820
rect 54251 6817 54263 6851
rect 54205 6811 54263 6817
rect 55490 6808 55496 6860
rect 55548 6848 55554 6860
rect 56244 6857 56272 6888
rect 56594 6876 56600 6888
rect 56652 6876 56658 6928
rect 56229 6851 56287 6857
rect 56229 6848 56241 6851
rect 55548 6820 56241 6848
rect 55548 6808 55554 6820
rect 56229 6817 56241 6820
rect 56275 6817 56287 6851
rect 56229 6811 56287 6817
rect 56778 6808 56784 6860
rect 56836 6808 56842 6860
rect 57882 6848 57888 6860
rect 57072 6820 57888 6848
rect 57072 6789 57100 6820
rect 57882 6808 57888 6820
rect 57940 6808 57946 6860
rect 53009 6783 53067 6789
rect 53009 6749 53021 6783
rect 53055 6749 53067 6783
rect 54021 6783 54079 6789
rect 54021 6780 54033 6783
rect 53009 6743 53067 6749
rect 53484 6752 54033 6780
rect 49878 6712 49884 6724
rect 46716 6684 47440 6712
rect 47780 6684 49884 6712
rect 46716 6672 46722 6684
rect 39853 6647 39911 6653
rect 39853 6613 39865 6647
rect 39899 6613 39911 6647
rect 39853 6607 39911 6613
rect 41230 6604 41236 6656
rect 41288 6604 41294 6656
rect 41417 6647 41475 6653
rect 41417 6613 41429 6647
rect 41463 6644 41475 6647
rect 42794 6644 42800 6656
rect 41463 6616 42800 6644
rect 41463 6613 41475 6616
rect 41417 6607 41475 6613
rect 42794 6604 42800 6616
rect 42852 6604 42858 6656
rect 43622 6604 43628 6656
rect 43680 6604 43686 6656
rect 44729 6647 44787 6653
rect 44729 6613 44741 6647
rect 44775 6644 44787 6647
rect 44818 6644 44824 6656
rect 44775 6616 44824 6644
rect 44775 6613 44787 6616
rect 44729 6607 44787 6613
rect 44818 6604 44824 6616
rect 44876 6604 44882 6656
rect 45738 6604 45744 6656
rect 45796 6604 45802 6656
rect 47486 6604 47492 6656
rect 47544 6644 47550 6656
rect 47780 6653 47808 6684
rect 49878 6672 49884 6684
rect 49936 6672 49942 6724
rect 51166 6712 51172 6724
rect 50356 6684 51172 6712
rect 47765 6647 47823 6653
rect 47765 6644 47777 6647
rect 47544 6616 47777 6644
rect 47544 6604 47550 6616
rect 47765 6613 47777 6616
rect 47811 6613 47823 6647
rect 47765 6607 47823 6613
rect 48038 6604 48044 6656
rect 48096 6644 48102 6656
rect 48133 6647 48191 6653
rect 48133 6644 48145 6647
rect 48096 6616 48145 6644
rect 48096 6604 48102 6616
rect 48133 6613 48145 6616
rect 48179 6613 48191 6647
rect 48133 6607 48191 6613
rect 48314 6604 48320 6656
rect 48372 6644 48378 6656
rect 48961 6647 49019 6653
rect 48961 6644 48973 6647
rect 48372 6616 48973 6644
rect 48372 6604 48378 6616
rect 48961 6613 48973 6616
rect 49007 6644 49019 6647
rect 49050 6644 49056 6656
rect 49007 6616 49056 6644
rect 49007 6613 49019 6616
rect 48961 6607 49019 6613
rect 49050 6604 49056 6616
rect 49108 6644 49114 6656
rect 49786 6644 49792 6656
rect 49108 6616 49792 6644
rect 49108 6604 49114 6616
rect 49786 6604 49792 6616
rect 49844 6604 49850 6656
rect 50246 6604 50252 6656
rect 50304 6644 50310 6656
rect 50356 6653 50384 6684
rect 51166 6672 51172 6684
rect 51224 6672 51230 6724
rect 50341 6647 50399 6653
rect 50341 6644 50353 6647
rect 50304 6616 50353 6644
rect 50304 6604 50310 6616
rect 50341 6613 50353 6616
rect 50387 6613 50399 6647
rect 50341 6607 50399 6613
rect 50798 6604 50804 6656
rect 50856 6644 50862 6656
rect 50893 6647 50951 6653
rect 50893 6644 50905 6647
rect 50856 6616 50905 6644
rect 50856 6604 50862 6616
rect 50893 6613 50905 6616
rect 50939 6644 50951 6647
rect 51261 6647 51319 6653
rect 51261 6644 51273 6647
rect 50939 6616 51273 6644
rect 50939 6613 50951 6616
rect 50893 6607 50951 6613
rect 51261 6613 51273 6616
rect 51307 6644 51319 6647
rect 51994 6644 52000 6656
rect 51307 6616 52000 6644
rect 51307 6613 51319 6616
rect 51261 6607 51319 6613
rect 51994 6604 52000 6616
rect 52052 6604 52058 6656
rect 52270 6604 52276 6656
rect 52328 6644 52334 6656
rect 52549 6647 52607 6653
rect 52549 6644 52561 6647
rect 52328 6616 52561 6644
rect 52328 6604 52334 6616
rect 52549 6613 52561 6616
rect 52595 6613 52607 6647
rect 52549 6607 52607 6613
rect 52917 6647 52975 6653
rect 52917 6613 52929 6647
rect 52963 6644 52975 6647
rect 53098 6644 53104 6656
rect 52963 6616 53104 6644
rect 52963 6613 52975 6616
rect 52917 6607 52975 6613
rect 53098 6604 53104 6616
rect 53156 6604 53162 6656
rect 53377 6647 53435 6653
rect 53377 6613 53389 6647
rect 53423 6644 53435 6647
rect 53484 6644 53512 6752
rect 54021 6749 54033 6752
rect 54067 6749 54079 6783
rect 54021 6743 54079 6749
rect 54757 6783 54815 6789
rect 54757 6749 54769 6783
rect 54803 6749 54815 6783
rect 54757 6743 54815 6749
rect 57057 6783 57115 6789
rect 57057 6749 57069 6783
rect 57103 6749 57115 6783
rect 58069 6783 58127 6789
rect 58069 6780 58081 6783
rect 57057 6743 57115 6749
rect 57440 6752 58081 6780
rect 53423 6616 53512 6644
rect 53423 6613 53435 6616
rect 53377 6607 53435 6613
rect 54110 6604 54116 6656
rect 54168 6644 54174 6656
rect 54772 6644 54800 6743
rect 56045 6715 56103 6721
rect 56045 6681 56057 6715
rect 56091 6712 56103 6715
rect 56091 6684 57008 6712
rect 56091 6681 56103 6684
rect 56045 6675 56103 6681
rect 56980 6656 57008 6684
rect 54168 6616 54800 6644
rect 55677 6647 55735 6653
rect 54168 6604 54174 6616
rect 55677 6613 55689 6647
rect 55723 6644 55735 6647
rect 55950 6644 55956 6656
rect 55723 6616 55956 6644
rect 55723 6613 55735 6616
rect 55677 6607 55735 6613
rect 55950 6604 55956 6616
rect 56008 6604 56014 6656
rect 56137 6647 56195 6653
rect 56137 6613 56149 6647
rect 56183 6644 56195 6647
rect 56778 6644 56784 6656
rect 56183 6616 56784 6644
rect 56183 6613 56195 6616
rect 56137 6607 56195 6613
rect 56778 6604 56784 6616
rect 56836 6604 56842 6656
rect 56962 6604 56968 6656
rect 57020 6604 57026 6656
rect 57440 6653 57468 6752
rect 58069 6749 58081 6752
rect 58115 6749 58127 6783
rect 58069 6743 58127 6749
rect 58529 6783 58587 6789
rect 58529 6749 58541 6783
rect 58575 6749 58587 6783
rect 58529 6743 58587 6749
rect 57974 6672 57980 6724
rect 58032 6712 58038 6724
rect 58544 6712 58572 6743
rect 58032 6684 58572 6712
rect 58032 6672 58038 6684
rect 57425 6647 57483 6653
rect 57425 6613 57437 6647
rect 57471 6613 57483 6647
rect 57425 6607 57483 6613
rect 57514 6604 57520 6656
rect 57572 6604 57578 6656
rect 58342 6604 58348 6656
rect 58400 6604 58406 6656
rect 1104 6554 59040 6576
rect 1104 6502 15394 6554
rect 15446 6502 15458 6554
rect 15510 6502 15522 6554
rect 15574 6502 15586 6554
rect 15638 6502 15650 6554
rect 15702 6502 29838 6554
rect 29890 6502 29902 6554
rect 29954 6502 29966 6554
rect 30018 6502 30030 6554
rect 30082 6502 30094 6554
rect 30146 6502 44282 6554
rect 44334 6502 44346 6554
rect 44398 6502 44410 6554
rect 44462 6502 44474 6554
rect 44526 6502 44538 6554
rect 44590 6502 58726 6554
rect 58778 6502 58790 6554
rect 58842 6502 58854 6554
rect 58906 6502 58918 6554
rect 58970 6502 58982 6554
rect 59034 6502 59040 6554
rect 1104 6480 59040 6502
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6440 6975 6443
rect 7742 6440 7748 6452
rect 6963 6412 7748 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7742 6400 7748 6412
rect 7800 6440 7806 6452
rect 8202 6440 8208 6452
rect 7800 6412 8208 6440
rect 7800 6400 7806 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8570 6400 8576 6452
rect 8628 6400 8634 6452
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10042 6440 10048 6452
rect 9907 6412 10048 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11606 6440 11612 6452
rect 11563 6412 11612 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 13906 6440 13912 6452
rect 12483 6412 13912 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 14369 6443 14427 6449
rect 14369 6409 14381 6443
rect 14415 6440 14427 6443
rect 14734 6440 14740 6452
rect 14415 6412 14740 6440
rect 14415 6409 14427 6412
rect 14369 6403 14427 6409
rect 5994 6332 6000 6384
rect 6052 6332 6058 6384
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 8122 6375 8180 6381
rect 8122 6372 8134 6375
rect 7616 6344 8134 6372
rect 7616 6332 7622 6344
rect 8122 6341 8134 6344
rect 8168 6341 8180 6375
rect 8122 6335 8180 6341
rect 8588 6372 8616 6400
rect 10226 6381 10232 6384
rect 10220 6372 10232 6381
rect 8588 6344 9996 6372
rect 10187 6344 10232 6372
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5442 6304 5448 6316
rect 5399 6276 5448 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 7374 6304 7380 6316
rect 5736 6276 7380 6304
rect 5736 6248 5764 6276
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 8588 6304 8616 6344
rect 8435 6276 8616 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9493 6307 9551 6313
rect 9088 6276 9168 6304
rect 9088 6264 9094 6276
rect 3326 6196 3332 6248
rect 3384 6196 3390 6248
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 2363 6140 3280 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 3252 6112 3280 6140
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 4080 6168 4108 6199
rect 4982 6196 4988 6248
rect 5040 6196 5046 6248
rect 5718 6196 5724 6248
rect 5776 6196 5782 6248
rect 7006 6196 7012 6248
rect 7064 6196 7070 6248
rect 9140 6245 9168 6276
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9582 6304 9588 6316
rect 9539 6276 9588 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9968 6313 9996 6344
rect 10220 6335 10232 6344
rect 10226 6332 10232 6335
rect 10284 6332 10290 6384
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 14292 6313 14320 6400
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 11974 6196 11980 6248
rect 12032 6196 12038 6248
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 13219 6239 13277 6245
rect 13219 6236 13231 6239
rect 12406 6208 13231 6236
rect 7024 6168 7052 6196
rect 4028 6140 7052 6168
rect 4028 6128 4034 6140
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 12406 6168 12434 6208
rect 13219 6205 13231 6208
rect 13265 6205 13277 6239
rect 13219 6199 13277 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 14093 6239 14151 6245
rect 13403 6208 13584 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 11388 6140 12434 6168
rect 11388 6128 11394 6140
rect 2682 6060 2688 6112
rect 2740 6060 2746 6112
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 3234 6060 3240 6112
rect 3292 6060 3298 6112
rect 3510 6060 3516 6112
rect 3568 6060 3574 6112
rect 4430 6060 4436 6112
rect 4488 6060 4494 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7190 6100 7196 6112
rect 7055 6072 7196 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7190 6060 7196 6072
rect 7248 6100 7254 6112
rect 8018 6100 8024 6112
rect 7248 6072 8024 6100
rect 7248 6060 7254 6072
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 13556 6100 13584 6208
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14384 6236 14412 6403
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 16758 6400 16764 6452
rect 16816 6400 16822 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 18141 6443 18199 6449
rect 18141 6440 18153 6443
rect 17368 6412 18153 6440
rect 17368 6400 17374 6412
rect 18141 6409 18153 6412
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 18506 6400 18512 6452
rect 18564 6400 18570 6452
rect 18782 6400 18788 6452
rect 18840 6440 18846 6452
rect 18969 6443 19027 6449
rect 18969 6440 18981 6443
rect 18840 6412 18981 6440
rect 18840 6400 18846 6412
rect 18969 6409 18981 6412
rect 19015 6409 19027 6443
rect 18969 6403 19027 6409
rect 19610 6400 19616 6452
rect 19668 6400 19674 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 19760 6412 22416 6440
rect 19760 6400 19766 6412
rect 15504 6375 15562 6381
rect 15504 6341 15516 6375
rect 15550 6372 15562 6375
rect 15841 6375 15899 6381
rect 15841 6372 15853 6375
rect 15550 6344 15853 6372
rect 15550 6341 15562 6344
rect 15504 6335 15562 6341
rect 15841 6341 15853 6344
rect 15887 6341 15899 6375
rect 16776 6372 16804 6400
rect 16914 6375 16972 6381
rect 16914 6372 16926 6375
rect 16776 6344 16926 6372
rect 15841 6335 15899 6341
rect 16914 6341 16926 6344
rect 16960 6341 16972 6375
rect 16914 6335 16972 6341
rect 18601 6375 18659 6381
rect 18601 6341 18613 6375
rect 18647 6372 18659 6375
rect 18647 6344 19564 6372
rect 18647 6341 18659 6344
rect 18601 6335 18659 6341
rect 19536 6316 19564 6344
rect 16666 6304 16672 6316
rect 15764 6276 16672 6304
rect 15764 6248 15792 6276
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 18472 6276 18828 6304
rect 18472 6264 18478 6276
rect 14139 6208 14412 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 15746 6196 15752 6248
rect 15804 6196 15810 6248
rect 16390 6196 16396 6248
rect 16448 6196 16454 6248
rect 13630 6128 13636 6180
rect 13688 6128 13694 6180
rect 18049 6171 18107 6177
rect 18049 6137 18061 6171
rect 18095 6168 18107 6171
rect 18432 6168 18460 6264
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 18800 6236 18828 6276
rect 19518 6264 19524 6316
rect 19576 6264 19582 6316
rect 19628 6313 19656 6400
rect 19886 6332 19892 6384
rect 19944 6372 19950 6384
rect 22278 6372 22284 6384
rect 19944 6344 22284 6372
rect 19944 6332 19950 6344
rect 22278 6332 22284 6344
rect 22336 6332 22342 6384
rect 19613 6307 19671 6313
rect 19613 6273 19625 6307
rect 19659 6273 19671 6307
rect 20254 6304 20260 6316
rect 19613 6267 19671 6273
rect 19720 6276 20260 6304
rect 19720 6236 19748 6276
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20806 6264 20812 6316
rect 20864 6313 20870 6316
rect 20864 6267 20876 6313
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21358 6304 21364 6316
rect 21131 6276 21364 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 20864 6264 20870 6267
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 22388 6313 22416 6412
rect 25130 6400 25136 6452
rect 25188 6400 25194 6452
rect 25225 6443 25283 6449
rect 25225 6409 25237 6443
rect 25271 6440 25283 6443
rect 26050 6440 26056 6452
rect 25271 6412 26056 6440
rect 25271 6409 25283 6412
rect 25225 6403 25283 6409
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 29917 6443 29975 6449
rect 26160 6412 27108 6440
rect 23109 6375 23167 6381
rect 23109 6341 23121 6375
rect 23155 6372 23167 6375
rect 23934 6372 23940 6384
rect 23155 6344 23940 6372
rect 23155 6341 23167 6344
rect 23109 6335 23167 6341
rect 23934 6332 23940 6344
rect 23992 6332 23998 6384
rect 25148 6372 25176 6400
rect 24136 6344 25176 6372
rect 24136 6313 24164 6344
rect 25314 6332 25320 6384
rect 25372 6372 25378 6384
rect 26160 6372 26188 6412
rect 25372 6344 26188 6372
rect 26360 6375 26418 6381
rect 25372 6332 25378 6344
rect 26360 6341 26372 6375
rect 26406 6372 26418 6375
rect 26973 6375 27031 6381
rect 26973 6372 26985 6375
rect 26406 6344 26985 6372
rect 26406 6341 26418 6344
rect 26360 6335 26418 6341
rect 26973 6341 26985 6344
rect 27019 6341 27031 6375
rect 27080 6372 27108 6412
rect 29917 6409 29929 6443
rect 29963 6409 29975 6443
rect 29917 6403 29975 6409
rect 29932 6372 29960 6403
rect 37182 6400 37188 6452
rect 37240 6440 37246 6452
rect 40221 6443 40279 6449
rect 37240 6412 37872 6440
rect 37240 6400 37246 6412
rect 31018 6372 31024 6384
rect 27080 6344 28948 6372
rect 29932 6344 31024 6372
rect 26973 6335 27031 6341
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6304 23075 6307
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 23063 6276 23489 6304
rect 23063 6273 23075 6276
rect 23017 6267 23075 6273
rect 23477 6273 23489 6276
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 24762 6264 24768 6316
rect 24820 6264 24826 6316
rect 24949 6307 25007 6313
rect 24949 6273 24961 6307
rect 24995 6304 25007 6307
rect 26510 6304 26516 6316
rect 24995 6276 26516 6304
rect 24995 6273 25007 6276
rect 24949 6267 25007 6273
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 27154 6264 27160 6316
rect 27212 6304 27218 6316
rect 28810 6313 28816 6316
rect 27525 6307 27583 6313
rect 27525 6304 27537 6307
rect 27212 6276 27537 6304
rect 27212 6264 27218 6276
rect 27525 6273 27537 6276
rect 27571 6273 27583 6307
rect 27525 6267 27583 6273
rect 28793 6307 28816 6313
rect 28793 6273 28805 6307
rect 28793 6267 28816 6273
rect 28810 6264 28816 6267
rect 28868 6264 28874 6316
rect 28920 6304 28948 6344
rect 31018 6332 31024 6344
rect 31076 6332 31082 6384
rect 32214 6372 32220 6384
rect 31864 6344 32220 6372
rect 28920 6276 30420 6304
rect 18800 6208 19748 6236
rect 23201 6239 23259 6245
rect 23201 6205 23213 6239
rect 23247 6205 23259 6239
rect 23201 6199 23259 6205
rect 26605 6239 26663 6245
rect 26605 6205 26617 6239
rect 26651 6236 26663 6239
rect 28537 6239 28595 6245
rect 28537 6236 28549 6239
rect 26651 6208 27752 6236
rect 26651 6205 26663 6208
rect 26605 6199 26663 6205
rect 18095 6140 18460 6168
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 11756 6072 13584 6100
rect 18708 6100 18736 6196
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 23216 6168 23244 6199
rect 21692 6140 23244 6168
rect 21692 6128 21698 6140
rect 23658 6128 23664 6180
rect 23716 6168 23722 6180
rect 24489 6171 24547 6177
rect 24489 6168 24501 6171
rect 23716 6140 24501 6168
rect 23716 6128 23722 6140
rect 24489 6137 24501 6140
rect 24535 6168 24547 6171
rect 24535 6140 25084 6168
rect 24535 6137 24547 6140
rect 24489 6131 24547 6137
rect 25056 6112 25084 6140
rect 21082 6100 21088 6112
rect 18708 6072 21088 6100
rect 11756 6060 11762 6072
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21232 6072 21833 6100
rect 21232 6060 21238 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 22649 6103 22707 6109
rect 22649 6069 22661 6103
rect 22695 6100 22707 6103
rect 23014 6100 23020 6112
rect 22695 6072 23020 6100
rect 22695 6069 22707 6072
rect 22649 6063 22707 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 25038 6060 25044 6112
rect 25096 6060 25102 6112
rect 27614 6060 27620 6112
rect 27672 6100 27678 6112
rect 27724 6100 27752 6208
rect 28368 6208 28549 6236
rect 28368 6109 28396 6208
rect 28537 6205 28549 6208
rect 28583 6205 28595 6239
rect 28537 6199 28595 6205
rect 27893 6103 27951 6109
rect 27893 6100 27905 6103
rect 27672 6072 27905 6100
rect 27672 6060 27678 6072
rect 27893 6069 27905 6072
rect 27939 6100 27951 6103
rect 28353 6103 28411 6109
rect 28353 6100 28365 6103
rect 27939 6072 28365 6100
rect 27939 6069 27951 6072
rect 27893 6063 27951 6069
rect 28353 6069 28365 6072
rect 28399 6069 28411 6103
rect 28353 6063 28411 6069
rect 30009 6103 30067 6109
rect 30009 6069 30021 6103
rect 30055 6100 30067 6103
rect 30190 6100 30196 6112
rect 30055 6072 30196 6100
rect 30055 6069 30067 6072
rect 30009 6063 30067 6069
rect 30190 6060 30196 6072
rect 30248 6060 30254 6112
rect 30392 6100 30420 6276
rect 31110 6264 31116 6316
rect 31168 6313 31174 6316
rect 31168 6267 31180 6313
rect 31168 6264 31174 6267
rect 31386 6196 31392 6248
rect 31444 6196 31450 6248
rect 31864 6109 31892 6344
rect 32214 6332 32220 6344
rect 32272 6372 32278 6384
rect 34885 6375 34943 6381
rect 34885 6372 34897 6375
rect 32272 6344 34897 6372
rect 32272 6332 32278 6344
rect 33226 6264 33232 6316
rect 33284 6313 33290 6316
rect 33612 6313 33640 6344
rect 34885 6341 34897 6344
rect 34931 6341 34943 6375
rect 35250 6372 35256 6384
rect 34885 6335 34943 6341
rect 35176 6344 35256 6372
rect 35176 6313 35204 6344
rect 35250 6332 35256 6344
rect 35308 6332 35314 6384
rect 35434 6381 35440 6384
rect 35428 6372 35440 6381
rect 35395 6344 35440 6372
rect 35428 6335 35440 6344
rect 35434 6332 35440 6335
rect 35492 6332 35498 6384
rect 35526 6332 35532 6384
rect 35584 6332 35590 6384
rect 36262 6332 36268 6384
rect 36320 6372 36326 6384
rect 36320 6344 36952 6372
rect 36320 6332 36326 6344
rect 33284 6267 33296 6313
rect 33597 6307 33655 6313
rect 33597 6273 33609 6307
rect 33643 6273 33655 6307
rect 33597 6267 33655 6273
rect 35161 6307 35219 6313
rect 35161 6273 35173 6307
rect 35207 6273 35219 6307
rect 35544 6304 35572 6332
rect 35161 6267 35219 6273
rect 35268 6276 35572 6304
rect 33284 6264 33290 6267
rect 33505 6239 33563 6245
rect 33505 6205 33517 6239
rect 33551 6205 33563 6239
rect 33505 6199 33563 6205
rect 33520 6168 33548 6199
rect 34422 6196 34428 6248
rect 34480 6236 34486 6248
rect 35268 6236 35296 6276
rect 36446 6264 36452 6316
rect 36504 6264 36510 6316
rect 36924 6313 36952 6344
rect 36909 6307 36967 6313
rect 36909 6273 36921 6307
rect 36955 6304 36967 6307
rect 37458 6304 37464 6316
rect 36955 6276 37464 6304
rect 36955 6273 36967 6276
rect 36909 6267 36967 6273
rect 37458 6264 37464 6276
rect 37516 6264 37522 6316
rect 37844 6313 37872 6412
rect 40221 6409 40233 6443
rect 40267 6440 40279 6443
rect 41230 6440 41236 6452
rect 40267 6412 41236 6440
rect 40267 6409 40279 6412
rect 40221 6403 40279 6409
rect 41230 6400 41236 6412
rect 41288 6400 41294 6452
rect 42058 6400 42064 6452
rect 42116 6440 42122 6452
rect 42116 6412 42840 6440
rect 42116 6400 42122 6412
rect 38657 6375 38715 6381
rect 38657 6372 38669 6375
rect 37936 6344 38669 6372
rect 37829 6307 37887 6313
rect 37829 6273 37841 6307
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 34480 6208 35296 6236
rect 34480 6196 34486 6208
rect 36170 6196 36176 6248
rect 36228 6196 36234 6248
rect 36464 6236 36492 6264
rect 37936 6236 37964 6344
rect 38657 6341 38669 6344
rect 38703 6372 38715 6375
rect 40494 6372 40500 6384
rect 38703 6344 40500 6372
rect 38703 6341 38715 6344
rect 38657 6335 38715 6341
rect 40494 6332 40500 6344
rect 40552 6332 40558 6384
rect 42245 6375 42303 6381
rect 42245 6341 42257 6375
rect 42291 6372 42303 6375
rect 42674 6375 42732 6381
rect 42674 6372 42686 6375
rect 42291 6344 42686 6372
rect 42291 6341 42303 6344
rect 42245 6335 42303 6341
rect 42674 6341 42686 6344
rect 42720 6341 42732 6375
rect 42812 6372 42840 6412
rect 43070 6400 43076 6452
rect 43128 6440 43134 6452
rect 43809 6443 43867 6449
rect 43809 6440 43821 6443
rect 43128 6412 43821 6440
rect 43128 6400 43134 6412
rect 43809 6409 43821 6412
rect 43855 6409 43867 6443
rect 43809 6403 43867 6409
rect 43622 6372 43628 6384
rect 42812 6344 43628 6372
rect 42674 6335 42732 6341
rect 43622 6332 43628 6344
rect 43680 6332 43686 6384
rect 39114 6313 39120 6316
rect 39097 6307 39120 6313
rect 39097 6273 39109 6307
rect 39097 6267 39120 6273
rect 39114 6264 39120 6267
rect 39172 6264 39178 6316
rect 40402 6264 40408 6316
rect 40460 6304 40466 6316
rect 43824 6304 43852 6403
rect 45738 6400 45744 6452
rect 45796 6400 45802 6452
rect 48774 6400 48780 6452
rect 48832 6400 48838 6452
rect 51629 6443 51687 6449
rect 51629 6440 51641 6443
rect 49160 6412 51641 6440
rect 44082 6332 44088 6384
rect 44140 6372 44146 6384
rect 44818 6372 44824 6384
rect 44140 6344 44824 6372
rect 44140 6332 44146 6344
rect 44818 6332 44824 6344
rect 44876 6372 44882 6384
rect 45364 6375 45422 6381
rect 44876 6344 45324 6372
rect 44876 6332 44882 6344
rect 44453 6307 44511 6313
rect 44453 6304 44465 6307
rect 40460 6276 43760 6304
rect 43824 6276 44465 6304
rect 40460 6264 40466 6276
rect 36464 6208 37964 6236
rect 38654 6196 38660 6248
rect 38712 6236 38718 6248
rect 38841 6239 38899 6245
rect 38841 6236 38853 6239
rect 38712 6208 38853 6236
rect 38712 6196 38718 6208
rect 38841 6205 38853 6208
rect 38887 6205 38899 6239
rect 38841 6199 38899 6205
rect 40862 6196 40868 6248
rect 40920 6196 40926 6248
rect 41690 6196 41696 6248
rect 41748 6196 41754 6248
rect 42429 6239 42487 6245
rect 42429 6205 42441 6239
rect 42475 6205 42487 6239
rect 42429 6199 42487 6205
rect 33594 6168 33600 6180
rect 33520 6140 33600 6168
rect 33594 6128 33600 6140
rect 33652 6128 33658 6180
rect 36188 6168 36216 6196
rect 38197 6171 38255 6177
rect 38197 6168 38209 6171
rect 36188 6140 38209 6168
rect 38197 6137 38209 6140
rect 38243 6168 38255 6171
rect 38746 6168 38752 6180
rect 38243 6140 38752 6168
rect 38243 6137 38255 6140
rect 38197 6131 38255 6137
rect 38746 6128 38752 6140
rect 38804 6128 38810 6180
rect 42444 6168 42472 6199
rect 41386 6140 42472 6168
rect 43732 6168 43760 6276
rect 44453 6273 44465 6276
rect 44499 6273 44511 6307
rect 44453 6267 44511 6273
rect 45097 6307 45155 6313
rect 45097 6273 45109 6307
rect 45143 6304 45155 6307
rect 45186 6304 45192 6316
rect 45143 6276 45192 6304
rect 45143 6273 45155 6276
rect 45097 6267 45155 6273
rect 45186 6264 45192 6276
rect 45244 6264 45250 6316
rect 45296 6304 45324 6344
rect 45364 6341 45376 6375
rect 45410 6372 45422 6375
rect 45756 6372 45784 6400
rect 45410 6344 45784 6372
rect 45410 6341 45422 6344
rect 45364 6335 45422 6341
rect 48314 6304 48320 6316
rect 45296 6276 48320 6304
rect 48314 6264 48320 6276
rect 48372 6264 48378 6316
rect 47118 6236 47124 6248
rect 46492 6208 47124 6236
rect 46492 6177 46520 6208
rect 47118 6196 47124 6208
rect 47176 6196 47182 6248
rect 48792 6236 48820 6400
rect 49053 6239 49111 6245
rect 49053 6236 49065 6239
rect 48792 6208 49065 6236
rect 49053 6205 49065 6208
rect 49099 6205 49111 6239
rect 49053 6199 49111 6205
rect 46477 6171 46535 6177
rect 43732 6140 45140 6168
rect 31849 6103 31907 6109
rect 31849 6100 31861 6103
rect 30392 6072 31861 6100
rect 31849 6069 31861 6072
rect 31895 6069 31907 6103
rect 31849 6063 31907 6069
rect 32125 6103 32183 6109
rect 32125 6069 32137 6103
rect 32171 6100 32183 6103
rect 32766 6100 32772 6112
rect 32171 6072 32772 6100
rect 32171 6069 32183 6072
rect 32125 6063 32183 6069
rect 32766 6060 32772 6072
rect 32824 6060 32830 6112
rect 36538 6060 36544 6112
rect 36596 6060 36602 6112
rect 36906 6060 36912 6112
rect 36964 6100 36970 6112
rect 37277 6103 37335 6109
rect 37277 6100 37289 6103
rect 36964 6072 37289 6100
rect 36964 6060 36970 6072
rect 37277 6069 37289 6072
rect 37323 6069 37335 6103
rect 37277 6063 37335 6069
rect 39758 6060 39764 6112
rect 39816 6100 39822 6112
rect 40313 6103 40371 6109
rect 40313 6100 40325 6103
rect 39816 6072 40325 6100
rect 39816 6060 39822 6072
rect 40313 6069 40325 6072
rect 40359 6069 40371 6103
rect 40313 6063 40371 6069
rect 41138 6060 41144 6112
rect 41196 6100 41202 6112
rect 41233 6103 41291 6109
rect 41233 6100 41245 6103
rect 41196 6072 41245 6100
rect 41196 6060 41202 6072
rect 41233 6069 41245 6072
rect 41279 6100 41291 6103
rect 41386 6100 41414 6140
rect 41279 6072 41414 6100
rect 41279 6069 41291 6072
rect 41233 6063 41291 6069
rect 43346 6060 43352 6112
rect 43404 6100 43410 6112
rect 43901 6103 43959 6109
rect 43901 6100 43913 6103
rect 43404 6072 43913 6100
rect 43404 6060 43410 6072
rect 43901 6069 43913 6072
rect 43947 6069 43959 6103
rect 43901 6063 43959 6069
rect 44818 6060 44824 6112
rect 44876 6060 44882 6112
rect 45112 6100 45140 6140
rect 46477 6137 46489 6171
rect 46523 6137 46535 6171
rect 48130 6168 48136 6180
rect 46477 6131 46535 6137
rect 47780 6140 48136 6168
rect 46198 6100 46204 6112
rect 45112 6072 46204 6100
rect 46198 6060 46204 6072
rect 46256 6060 46262 6112
rect 46566 6060 46572 6112
rect 46624 6060 46630 6112
rect 47670 6060 47676 6112
rect 47728 6100 47734 6112
rect 47780 6109 47808 6140
rect 48130 6128 48136 6140
rect 48188 6168 48194 6180
rect 49160 6168 49188 6412
rect 51629 6409 51641 6412
rect 51675 6409 51687 6443
rect 51629 6403 51687 6409
rect 51813 6443 51871 6449
rect 51813 6409 51825 6443
rect 51859 6440 51871 6443
rect 51902 6440 51908 6452
rect 51859 6412 51908 6440
rect 51859 6409 51871 6412
rect 51813 6403 51871 6409
rect 49237 6375 49295 6381
rect 49237 6341 49249 6375
rect 49283 6372 49295 6375
rect 50525 6375 50583 6381
rect 50525 6372 50537 6375
rect 49283 6344 50537 6372
rect 49283 6341 49295 6344
rect 49237 6335 49295 6341
rect 50525 6341 50537 6344
rect 50571 6341 50583 6375
rect 50525 6335 50583 6341
rect 49329 6307 49387 6313
rect 49329 6273 49341 6307
rect 49375 6304 49387 6307
rect 49602 6304 49608 6316
rect 49375 6276 49608 6304
rect 49375 6273 49387 6276
rect 49329 6267 49387 6273
rect 49602 6264 49608 6276
rect 49660 6264 49666 6316
rect 50341 6239 50399 6245
rect 50341 6236 50353 6239
rect 49712 6208 50353 6236
rect 49712 6177 49740 6208
rect 50341 6205 50353 6208
rect 50387 6205 50399 6239
rect 50341 6199 50399 6205
rect 51074 6196 51080 6248
rect 51132 6196 51138 6248
rect 51644 6236 51672 6403
rect 51902 6400 51908 6412
rect 51960 6400 51966 6452
rect 52181 6443 52239 6449
rect 52181 6409 52193 6443
rect 52227 6440 52239 6443
rect 53098 6440 53104 6452
rect 52227 6412 53104 6440
rect 52227 6409 52239 6412
rect 52181 6403 52239 6409
rect 53098 6400 53104 6412
rect 53156 6400 53162 6452
rect 53190 6400 53196 6452
rect 53248 6400 53254 6452
rect 54110 6400 54116 6452
rect 54168 6400 54174 6452
rect 57514 6440 57520 6452
rect 57440 6412 57520 6440
rect 53000 6375 53058 6381
rect 53000 6341 53012 6375
rect 53046 6372 53058 6375
rect 53208 6372 53236 6400
rect 53046 6344 53236 6372
rect 53046 6341 53058 6344
rect 53000 6335 53058 6341
rect 52273 6307 52331 6313
rect 52273 6273 52285 6307
rect 52319 6304 52331 6307
rect 52546 6304 52552 6316
rect 52319 6276 52552 6304
rect 52319 6273 52331 6276
rect 52273 6267 52331 6273
rect 52546 6264 52552 6276
rect 52604 6264 52610 6316
rect 52733 6307 52791 6313
rect 52733 6273 52745 6307
rect 52779 6304 52791 6307
rect 52822 6304 52828 6316
rect 52779 6276 52828 6304
rect 52779 6273 52791 6276
rect 52733 6267 52791 6273
rect 52822 6264 52828 6276
rect 52880 6264 52886 6316
rect 52365 6239 52423 6245
rect 52365 6236 52377 6239
rect 51644 6208 52377 6236
rect 52365 6205 52377 6208
rect 52411 6205 52423 6239
rect 54128 6236 54156 6400
rect 54938 6264 54944 6316
rect 54996 6264 55002 6316
rect 57440 6313 57468 6412
rect 57514 6400 57520 6412
rect 57572 6400 57578 6452
rect 57882 6400 57888 6452
rect 57940 6400 57946 6452
rect 57440 6307 57503 6313
rect 57440 6276 57457 6307
rect 57445 6273 57457 6276
rect 57491 6273 57503 6307
rect 57445 6267 57503 6273
rect 57698 6264 57704 6316
rect 57756 6264 57762 6316
rect 55079 6239 55137 6245
rect 55079 6236 55091 6239
rect 54128 6208 55091 6236
rect 52365 6199 52423 6205
rect 55079 6205 55091 6208
rect 55125 6205 55137 6239
rect 55079 6199 55137 6205
rect 55214 6196 55220 6248
rect 55272 6196 55278 6248
rect 55493 6239 55551 6245
rect 55493 6205 55505 6239
rect 55539 6236 55551 6239
rect 55582 6236 55588 6248
rect 55539 6208 55588 6236
rect 55539 6205 55551 6208
rect 55493 6199 55551 6205
rect 55582 6196 55588 6208
rect 55640 6196 55646 6248
rect 55953 6239 56011 6245
rect 55953 6205 55965 6239
rect 55999 6205 56011 6239
rect 55953 6199 56011 6205
rect 56137 6239 56195 6245
rect 56137 6205 56149 6239
rect 56183 6236 56195 6239
rect 56686 6236 56692 6248
rect 56183 6208 56692 6236
rect 56183 6205 56195 6208
rect 56137 6199 56195 6205
rect 48188 6140 49188 6168
rect 49697 6171 49755 6177
rect 48188 6128 48194 6140
rect 49697 6137 49709 6171
rect 49743 6137 49755 6171
rect 49697 6131 49755 6137
rect 47765 6103 47823 6109
rect 47765 6100 47777 6103
rect 47728 6072 47777 6100
rect 47728 6060 47734 6072
rect 47765 6069 47777 6072
rect 47811 6069 47823 6103
rect 47765 6063 47823 6069
rect 48498 6060 48504 6112
rect 48556 6060 48562 6112
rect 49786 6060 49792 6112
rect 49844 6060 49850 6112
rect 54297 6103 54355 6109
rect 54297 6069 54309 6103
rect 54343 6100 54355 6103
rect 55858 6100 55864 6112
rect 54343 6072 55864 6100
rect 54343 6069 54355 6072
rect 54297 6063 54355 6069
rect 55858 6060 55864 6072
rect 55916 6060 55922 6112
rect 55968 6100 55996 6199
rect 56686 6196 56692 6208
rect 56744 6196 56750 6248
rect 57900 6245 57928 6400
rect 57885 6239 57943 6245
rect 57885 6205 57897 6239
rect 57931 6205 57943 6239
rect 57885 6199 57943 6205
rect 58437 6239 58495 6245
rect 58437 6205 58449 6239
rect 58483 6205 58495 6239
rect 58437 6199 58495 6205
rect 58452 6168 58480 6199
rect 57716 6140 58480 6168
rect 56321 6103 56379 6109
rect 56321 6100 56333 6103
rect 55968 6072 56333 6100
rect 56321 6069 56333 6072
rect 56367 6100 56379 6103
rect 57716 6100 57744 6140
rect 56367 6072 57744 6100
rect 56367 6069 56379 6072
rect 56321 6063 56379 6069
rect 1104 6010 58880 6032
rect 1104 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 22616 6010
rect 22668 5958 22680 6010
rect 22732 5958 22744 6010
rect 22796 5958 22808 6010
rect 22860 5958 22872 6010
rect 22924 5958 37060 6010
rect 37112 5958 37124 6010
rect 37176 5958 37188 6010
rect 37240 5958 37252 6010
rect 37304 5958 37316 6010
rect 37368 5958 51504 6010
rect 51556 5958 51568 6010
rect 51620 5958 51632 6010
rect 51684 5958 51696 6010
rect 51748 5958 51760 6010
rect 51812 5958 58880 6010
rect 1104 5936 58880 5958
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 5442 5896 5448 5908
rect 4295 5868 5448 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6178 5896 6184 5908
rect 6135 5868 6184 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6178 5856 6184 5868
rect 6236 5896 6242 5908
rect 6822 5896 6828 5908
rect 6236 5868 6828 5896
rect 6236 5856 6242 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 9732 5868 10701 5896
rect 9732 5856 9738 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 10689 5859 10747 5865
rect 11517 5899 11575 5905
rect 11517 5865 11529 5899
rect 11563 5896 11575 5899
rect 11974 5896 11980 5908
rect 11563 5868 11980 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12820 5868 14596 5896
rect 5721 5831 5779 5837
rect 5721 5797 5733 5831
rect 5767 5797 5779 5831
rect 7392 5828 7420 5856
rect 12820 5840 12848 5868
rect 10597 5831 10655 5837
rect 10597 5828 10609 5831
rect 7392 5800 10609 5828
rect 5721 5791 5779 5797
rect 10597 5797 10609 5800
rect 10643 5828 10655 5831
rect 10643 5800 12388 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 5736 5760 5764 5791
rect 7098 5760 7104 5772
rect 5736 5732 7104 5760
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 7742 5760 7748 5772
rect 7423 5732 7748 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 8018 5720 8024 5772
rect 8076 5720 8082 5772
rect 8754 5720 8760 5772
rect 8812 5760 8818 5772
rect 9306 5760 9312 5772
rect 8812 5732 9312 5760
rect 8812 5720 8818 5732
rect 9306 5720 9312 5732
rect 9364 5760 9370 5772
rect 9364 5732 9674 5760
rect 9364 5720 9370 5732
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 1762 5692 1768 5704
rect 1719 5664 1768 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 1762 5652 1768 5664
rect 1820 5692 1826 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1820 5664 2053 5692
rect 1820 5652 1826 5664
rect 2041 5661 2053 5664
rect 2087 5692 2099 5695
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 2087 5664 2145 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2133 5661 2145 5664
rect 2179 5692 2191 5695
rect 2682 5692 2688 5704
rect 2179 5664 2688 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2774 5652 2780 5704
rect 2832 5652 2838 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 2400 5627 2458 5633
rect 2400 5593 2412 5627
rect 2446 5624 2458 5627
rect 2792 5624 2820 5652
rect 2446 5596 2820 5624
rect 2446 5593 2458 5596
rect 2400 5587 2458 5593
rect 4356 5568 4384 5655
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4597 5695 4655 5701
rect 4597 5692 4609 5695
rect 4488 5664 4609 5692
rect 4488 5652 4494 5664
rect 4597 5661 4609 5664
rect 4643 5661 4655 5695
rect 4597 5655 4655 5661
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 7006 5701 7012 5704
rect 6984 5695 7012 5701
rect 6984 5661 6996 5695
rect 6984 5655 7012 5661
rect 7006 5652 7012 5655
rect 7064 5652 7070 5704
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 8128 5624 8156 5655
rect 8076 5596 8156 5624
rect 9646 5624 9674 5732
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 11238 5760 11244 5772
rect 10284 5732 11244 5760
rect 10284 5720 10290 5732
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11756 5732 12081 5760
rect 11756 5720 11762 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12360 5760 12388 5800
rect 12802 5788 12808 5840
rect 12860 5788 12866 5840
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 13630 5828 13636 5840
rect 12952 5800 13636 5828
rect 12952 5788 12958 5800
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5828 13783 5831
rect 14458 5828 14464 5840
rect 13771 5800 14464 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 14458 5788 14464 5800
rect 14516 5788 14522 5840
rect 13173 5763 13231 5769
rect 13173 5760 13185 5763
rect 12360 5732 13185 5760
rect 12069 5723 12127 5729
rect 13173 5729 13185 5732
rect 13219 5760 13231 5763
rect 14090 5760 14096 5772
rect 13219 5732 14096 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 14568 5760 14596 5868
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 16390 5896 16396 5908
rect 15243 5868 16396 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 17770 5856 17776 5908
rect 17828 5856 17834 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 20438 5896 20444 5908
rect 19484 5868 20444 5896
rect 19484 5856 19490 5868
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20864 5868 20913 5896
rect 20864 5856 20870 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 22278 5856 22284 5908
rect 22336 5856 22342 5908
rect 22462 5856 22468 5908
rect 22520 5856 22526 5908
rect 23014 5856 23020 5908
rect 23072 5856 23078 5908
rect 28445 5899 28503 5905
rect 28445 5865 28457 5899
rect 28491 5896 28503 5899
rect 28534 5896 28540 5908
rect 28491 5868 28540 5896
rect 28491 5865 28503 5868
rect 28445 5859 28503 5865
rect 28534 5856 28540 5868
rect 28592 5856 28598 5908
rect 30374 5896 30380 5908
rect 28736 5868 30380 5896
rect 14936 5828 14964 5856
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 14936 5800 17233 5828
rect 17221 5797 17233 5800
rect 17267 5828 17279 5831
rect 18690 5828 18696 5840
rect 17267 5800 18696 5828
rect 17267 5797 17279 5800
rect 17221 5791 17279 5797
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 18969 5831 19027 5837
rect 18969 5797 18981 5831
rect 19015 5828 19027 5831
rect 19886 5828 19892 5840
rect 19015 5800 19892 5828
rect 19015 5797 19027 5800
rect 18969 5791 19027 5797
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 20180 5800 21312 5828
rect 14642 5760 14648 5772
rect 14568 5732 14648 5760
rect 14642 5720 14648 5732
rect 14700 5760 14706 5772
rect 14700 5732 15240 5760
rect 14700 5720 14706 5732
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5692 10011 5695
rect 10134 5692 10140 5704
rect 9999 5664 10140 5692
rect 9999 5661 10011 5664
rect 9953 5655 10011 5661
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 14550 5692 14556 5704
rect 14200 5664 14556 5692
rect 12802 5624 12808 5636
rect 9646 5596 12808 5624
rect 8076 5584 8082 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13722 5624 13728 5636
rect 13412 5596 13728 5624
rect 13412 5584 13418 5596
rect 13722 5584 13728 5596
rect 13780 5624 13786 5636
rect 14200 5624 14228 5664
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 15212 5692 15240 5732
rect 15930 5720 15936 5772
rect 15988 5760 15994 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 15988 5732 17601 5760
rect 15988 5720 15994 5732
rect 17589 5729 17601 5732
rect 17635 5760 17647 5763
rect 17954 5760 17960 5772
rect 17635 5732 17960 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18322 5720 18328 5772
rect 18380 5720 18386 5772
rect 20180 5769 20208 5800
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19904 5732 20177 5760
rect 16298 5692 16304 5704
rect 15212 5664 16304 5692
rect 16298 5652 16304 5664
rect 16356 5692 16362 5704
rect 19904 5701 19932 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 21174 5760 21180 5772
rect 20165 5723 20223 5729
rect 20456 5732 21180 5760
rect 20456 5701 20484 5732
rect 21174 5720 21180 5732
rect 21232 5720 21238 5772
rect 21284 5760 21312 5800
rect 22922 5760 22928 5772
rect 21284 5732 22928 5760
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 23032 5769 23060 5856
rect 24578 5788 24584 5840
rect 24636 5828 24642 5840
rect 24673 5831 24731 5837
rect 24673 5828 24685 5831
rect 24636 5800 24685 5828
rect 24636 5788 24642 5800
rect 24673 5797 24685 5800
rect 24719 5797 24731 5831
rect 24673 5791 24731 5797
rect 25593 5831 25651 5837
rect 25593 5797 25605 5831
rect 25639 5797 25651 5831
rect 25593 5791 25651 5797
rect 23017 5763 23075 5769
rect 23017 5729 23029 5763
rect 23063 5729 23075 5763
rect 23017 5723 23075 5729
rect 19889 5695 19947 5701
rect 19889 5692 19901 5695
rect 16356 5664 19901 5692
rect 16356 5652 16362 5664
rect 19889 5661 19901 5664
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 20441 5655 20499 5661
rect 20824 5664 21465 5692
rect 15565 5627 15623 5633
rect 15565 5624 15577 5627
rect 13780 5596 14228 5624
rect 14292 5596 15577 5624
rect 13780 5584 13786 5596
rect 4338 5516 4344 5568
rect 4396 5516 4402 5568
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 7558 5556 7564 5568
rect 6227 5528 7564 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8720 5528 8769 5556
rect 8720 5516 8726 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 11054 5516 11060 5568
rect 11112 5516 11118 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11882 5556 11888 5568
rect 11195 5528 11888 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 12943 5528 13277 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13265 5519 13323 5525
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14292 5565 14320 5596
rect 15565 5593 15577 5596
rect 15611 5624 15623 5627
rect 15746 5624 15752 5636
rect 15611 5596 15752 5624
rect 15611 5593 15623 5596
rect 15565 5587 15623 5593
rect 15746 5584 15752 5596
rect 15804 5624 15810 5636
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 15804 5596 15945 5624
rect 15804 5584 15810 5596
rect 15933 5593 15945 5596
rect 15979 5624 15991 5627
rect 16206 5624 16212 5636
rect 15979 5596 16212 5624
rect 15979 5593 15991 5596
rect 15933 5587 15991 5593
rect 16206 5584 16212 5596
rect 16264 5624 16270 5636
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 16264 5596 16497 5624
rect 16264 5584 16270 5596
rect 16485 5593 16497 5596
rect 16531 5624 16543 5627
rect 16853 5627 16911 5633
rect 16853 5624 16865 5627
rect 16531 5596 16865 5624
rect 16531 5593 16543 5596
rect 16485 5587 16543 5593
rect 16853 5593 16865 5596
rect 16899 5593 16911 5627
rect 16853 5587 16911 5593
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 13872 5528 14289 5556
rect 13872 5516 13878 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14277 5519 14335 5525
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14608 5528 14749 5556
rect 14608 5516 14614 5528
rect 14737 5525 14749 5528
rect 14783 5525 14795 5559
rect 14737 5519 14795 5525
rect 19426 5516 19432 5568
rect 19484 5516 19490 5568
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 20254 5556 20260 5568
rect 19576 5528 20260 5556
rect 19576 5516 19582 5528
rect 20254 5516 20260 5528
rect 20312 5556 20318 5568
rect 20824 5565 20852 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 24026 5692 24032 5704
rect 21453 5655 21511 5661
rect 22756 5664 24032 5692
rect 21082 5584 21088 5636
rect 21140 5624 21146 5636
rect 22005 5627 22063 5633
rect 22005 5624 22017 5627
rect 21140 5596 22017 5624
rect 21140 5584 21146 5596
rect 22005 5593 22017 5596
rect 22051 5624 22063 5627
rect 22756 5624 22784 5664
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 24688 5692 24716 5791
rect 24949 5763 25007 5769
rect 24949 5729 24961 5763
rect 24995 5760 25007 5763
rect 25608 5760 25636 5791
rect 25866 5788 25872 5840
rect 25924 5828 25930 5840
rect 25924 5800 27476 5828
rect 25924 5788 25930 5800
rect 26145 5763 26203 5769
rect 26145 5760 26157 5763
rect 24995 5732 25636 5760
rect 25884 5732 26157 5760
rect 24995 5729 25007 5732
rect 24949 5723 25007 5729
rect 25501 5695 25559 5701
rect 24688 5664 25452 5692
rect 23477 5627 23535 5633
rect 23477 5624 23489 5627
rect 22051 5596 22784 5624
rect 22848 5596 23489 5624
rect 22051 5593 22063 5596
rect 22005 5587 22063 5593
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 20312 5528 20361 5556
rect 20312 5516 20318 5528
rect 20349 5525 20361 5528
rect 20395 5525 20407 5559
rect 20349 5519 20407 5525
rect 20809 5559 20867 5565
rect 20809 5525 20821 5559
rect 20855 5525 20867 5559
rect 20809 5519 20867 5525
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 22848 5556 22876 5596
rect 23477 5593 23489 5596
rect 23523 5624 23535 5627
rect 24762 5624 24768 5636
rect 23523 5596 24768 5624
rect 23523 5593 23535 5596
rect 23477 5587 23535 5593
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 25314 5584 25320 5636
rect 25372 5584 25378 5636
rect 25424 5624 25452 5664
rect 25501 5661 25513 5695
rect 25547 5692 25559 5695
rect 25590 5692 25596 5704
rect 25547 5664 25596 5692
rect 25547 5661 25559 5664
rect 25501 5655 25559 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 25884 5624 25912 5732
rect 26145 5729 26157 5732
rect 26191 5729 26203 5763
rect 26145 5723 26203 5729
rect 25961 5695 26019 5701
rect 25961 5661 25973 5695
rect 26007 5692 26019 5695
rect 26694 5692 26700 5704
rect 26007 5664 26700 5692
rect 26007 5661 26019 5664
rect 25961 5655 26019 5661
rect 26694 5652 26700 5664
rect 26752 5652 26758 5704
rect 26970 5652 26976 5704
rect 27028 5652 27034 5704
rect 27448 5701 27476 5800
rect 27433 5695 27491 5701
rect 27433 5661 27445 5695
rect 27479 5692 27491 5695
rect 27798 5692 27804 5704
rect 27479 5664 27804 5692
rect 27479 5661 27491 5664
rect 27433 5655 27491 5661
rect 27798 5652 27804 5664
rect 27856 5652 27862 5704
rect 28736 5624 28764 5868
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 33410 5856 33416 5908
rect 33468 5896 33474 5908
rect 33689 5899 33747 5905
rect 33689 5896 33701 5899
rect 33468 5868 33701 5896
rect 33468 5856 33474 5868
rect 33689 5865 33701 5868
rect 33735 5865 33747 5899
rect 33689 5859 33747 5865
rect 38013 5899 38071 5905
rect 38013 5865 38025 5899
rect 38059 5896 38071 5899
rect 38102 5896 38108 5908
rect 38059 5868 38108 5896
rect 38059 5865 38071 5868
rect 38013 5859 38071 5865
rect 38102 5856 38108 5868
rect 38160 5896 38166 5908
rect 38286 5896 38292 5908
rect 38160 5868 38292 5896
rect 38160 5856 38166 5868
rect 38286 5856 38292 5868
rect 38344 5856 38350 5908
rect 38470 5856 38476 5908
rect 38528 5856 38534 5908
rect 38654 5856 38660 5908
rect 38712 5896 38718 5908
rect 38749 5899 38807 5905
rect 38749 5896 38761 5899
rect 38712 5868 38761 5896
rect 38712 5856 38718 5868
rect 38749 5865 38761 5868
rect 38795 5896 38807 5899
rect 41138 5896 41144 5908
rect 38795 5868 41144 5896
rect 38795 5865 38807 5868
rect 38749 5859 38807 5865
rect 41138 5856 41144 5868
rect 41196 5856 41202 5908
rect 41690 5856 41696 5908
rect 41748 5896 41754 5908
rect 42337 5899 42395 5905
rect 42337 5896 42349 5899
rect 41748 5868 42349 5896
rect 41748 5856 41754 5868
rect 42337 5865 42349 5868
rect 42383 5865 42395 5899
rect 42337 5859 42395 5865
rect 43622 5856 43628 5908
rect 43680 5896 43686 5908
rect 43717 5899 43775 5905
rect 43717 5896 43729 5899
rect 43680 5868 43729 5896
rect 43680 5856 43686 5868
rect 43717 5865 43729 5868
rect 43763 5865 43775 5899
rect 43717 5859 43775 5865
rect 46569 5899 46627 5905
rect 46569 5865 46581 5899
rect 46615 5896 46627 5899
rect 48593 5899 48651 5905
rect 46615 5868 47808 5896
rect 46615 5865 46627 5868
rect 46569 5859 46627 5865
rect 28828 5800 29684 5828
rect 28828 5769 28856 5800
rect 28813 5763 28871 5769
rect 28813 5729 28825 5763
rect 28859 5729 28871 5763
rect 28813 5723 28871 5729
rect 29656 5704 29684 5800
rect 32122 5788 32128 5840
rect 32180 5788 32186 5840
rect 33502 5828 33508 5840
rect 32600 5800 33508 5828
rect 30190 5720 30196 5772
rect 30248 5760 30254 5772
rect 32600 5769 32628 5800
rect 33502 5788 33508 5800
rect 33560 5828 33566 5840
rect 33870 5828 33876 5840
rect 33560 5800 33876 5828
rect 33560 5788 33566 5800
rect 33870 5788 33876 5800
rect 33928 5788 33934 5840
rect 35618 5788 35624 5840
rect 35676 5788 35682 5840
rect 38562 5788 38568 5840
rect 38620 5828 38626 5840
rect 41874 5828 41880 5840
rect 38620 5800 41880 5828
rect 38620 5788 38626 5800
rect 41874 5788 41880 5800
rect 41932 5828 41938 5840
rect 42058 5828 42064 5840
rect 41932 5800 42064 5828
rect 41932 5788 41938 5800
rect 42058 5788 42064 5800
rect 42116 5788 42122 5840
rect 47780 5772 47808 5868
rect 48593 5865 48605 5899
rect 48639 5896 48651 5899
rect 51074 5896 51080 5908
rect 48639 5868 51080 5896
rect 48639 5865 48651 5868
rect 48593 5859 48651 5865
rect 47854 5788 47860 5840
rect 47912 5788 47918 5840
rect 31849 5763 31907 5769
rect 31849 5760 31861 5763
rect 30248 5732 31861 5760
rect 30248 5720 30254 5732
rect 31849 5729 31861 5732
rect 31895 5729 31907 5763
rect 31849 5723 31907 5729
rect 32585 5763 32643 5769
rect 32585 5729 32597 5763
rect 32631 5729 32643 5763
rect 32585 5723 32643 5729
rect 33045 5763 33103 5769
rect 33045 5729 33057 5763
rect 33091 5760 33103 5763
rect 33318 5760 33324 5772
rect 33091 5732 33324 5760
rect 33091 5729 33103 5732
rect 33045 5723 33103 5729
rect 33318 5720 33324 5732
rect 33376 5720 33382 5772
rect 35253 5763 35311 5769
rect 35253 5760 35265 5763
rect 33428 5732 35265 5760
rect 29549 5695 29607 5701
rect 29549 5692 29561 5695
rect 25424 5596 28764 5624
rect 28808 5664 29561 5692
rect 21416 5528 22876 5556
rect 21416 5516 21422 5528
rect 22922 5516 22928 5568
rect 22980 5556 22986 5568
rect 24213 5559 24271 5565
rect 24213 5556 24225 5559
rect 22980 5528 24225 5556
rect 22980 5516 22986 5528
rect 24213 5525 24225 5528
rect 24259 5556 24271 5559
rect 25332 5556 25360 5584
rect 25774 5556 25780 5568
rect 24259 5528 25780 5556
rect 24259 5525 24271 5528
rect 24213 5519 24271 5525
rect 25774 5516 25780 5528
rect 25832 5516 25838 5568
rect 26053 5559 26111 5565
rect 26053 5525 26065 5559
rect 26099 5556 26111 5559
rect 26421 5559 26479 5565
rect 26421 5556 26433 5559
rect 26099 5528 26433 5556
rect 26099 5525 26111 5528
rect 26053 5519 26111 5525
rect 26421 5525 26433 5528
rect 26467 5525 26479 5559
rect 26421 5519 26479 5525
rect 27614 5516 27620 5568
rect 27672 5556 27678 5568
rect 27709 5559 27767 5565
rect 27709 5556 27721 5559
rect 27672 5528 27721 5556
rect 27672 5516 27678 5528
rect 27709 5525 27721 5528
rect 27755 5525 27767 5559
rect 27709 5519 27767 5525
rect 28169 5559 28227 5565
rect 28169 5525 28181 5559
rect 28215 5556 28227 5559
rect 28258 5556 28264 5568
rect 28215 5528 28264 5556
rect 28215 5525 28227 5528
rect 28169 5519 28227 5525
rect 28258 5516 28264 5528
rect 28316 5516 28322 5568
rect 28534 5516 28540 5568
rect 28592 5556 28598 5568
rect 28808 5556 28836 5664
rect 29549 5661 29561 5664
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 30377 5695 30435 5701
rect 30377 5692 30389 5695
rect 29696 5664 30389 5692
rect 29696 5652 29702 5664
rect 30377 5661 30389 5664
rect 30423 5692 30435 5695
rect 30926 5692 30932 5704
rect 30423 5664 30932 5692
rect 30423 5661 30435 5664
rect 30377 5655 30435 5661
rect 30926 5652 30932 5664
rect 30984 5652 30990 5704
rect 31570 5652 31576 5704
rect 31628 5652 31634 5704
rect 31754 5701 31760 5704
rect 31732 5695 31760 5701
rect 31732 5661 31744 5695
rect 31732 5655 31760 5661
rect 31754 5652 31760 5655
rect 31812 5652 31818 5704
rect 32766 5652 32772 5704
rect 32824 5692 32830 5704
rect 33428 5692 33456 5732
rect 35253 5729 35265 5732
rect 35299 5729 35311 5763
rect 35253 5723 35311 5729
rect 38746 5720 38752 5772
rect 38804 5760 38810 5772
rect 39485 5763 39543 5769
rect 39485 5760 39497 5763
rect 38804 5732 39497 5760
rect 38804 5720 38810 5732
rect 39485 5729 39497 5732
rect 39531 5729 39543 5763
rect 40126 5760 40132 5772
rect 39485 5723 39543 5729
rect 39776 5732 40132 5760
rect 32824 5664 33456 5692
rect 32824 5652 32830 5664
rect 33502 5652 33508 5704
rect 33560 5692 33566 5704
rect 34241 5695 34299 5701
rect 34241 5692 34253 5695
rect 33560 5664 34253 5692
rect 33560 5652 33566 5664
rect 34241 5661 34253 5664
rect 34287 5661 34299 5695
rect 34241 5655 34299 5661
rect 36745 5695 36803 5701
rect 36745 5661 36757 5695
rect 36791 5692 36803 5695
rect 36906 5692 36912 5704
rect 36791 5664 36912 5692
rect 36791 5661 36803 5664
rect 36745 5655 36803 5661
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 37001 5695 37059 5701
rect 37001 5661 37013 5695
rect 37047 5692 37059 5695
rect 37550 5692 37556 5704
rect 37047 5664 37556 5692
rect 37047 5661 37059 5664
rect 37001 5655 37059 5661
rect 37550 5652 37556 5664
rect 37608 5652 37614 5704
rect 37645 5695 37703 5701
rect 37645 5661 37657 5695
rect 37691 5661 37703 5695
rect 37645 5655 37703 5661
rect 39301 5695 39359 5701
rect 39301 5661 39313 5695
rect 39347 5692 39359 5695
rect 39776 5692 39804 5732
rect 40126 5720 40132 5732
rect 40184 5720 40190 5772
rect 40218 5720 40224 5772
rect 40276 5760 40282 5772
rect 42981 5763 43039 5769
rect 42981 5760 42993 5763
rect 40276 5732 42993 5760
rect 40276 5720 40282 5732
rect 42981 5729 42993 5732
rect 43027 5760 43039 5763
rect 44453 5763 44511 5769
rect 44453 5760 44465 5763
rect 43027 5732 44465 5760
rect 43027 5729 43039 5732
rect 42981 5723 43039 5729
rect 44453 5729 44465 5732
rect 44499 5729 44511 5763
rect 44453 5723 44511 5729
rect 45186 5720 45192 5772
rect 45244 5720 45250 5772
rect 47118 5720 47124 5772
rect 47176 5760 47182 5772
rect 47443 5763 47501 5769
rect 47443 5760 47455 5763
rect 47176 5732 47455 5760
rect 47176 5720 47182 5732
rect 47443 5729 47455 5732
rect 47489 5729 47501 5763
rect 47443 5723 47501 5729
rect 47581 5763 47639 5769
rect 47581 5729 47593 5763
rect 47627 5760 47639 5763
rect 47762 5760 47768 5772
rect 47627 5732 47768 5760
rect 47627 5729 47639 5732
rect 47581 5723 47639 5729
rect 47762 5720 47768 5732
rect 47820 5720 47826 5772
rect 48501 5763 48559 5769
rect 48501 5729 48513 5763
rect 48547 5760 48559 5763
rect 48608 5760 48636 5859
rect 51074 5856 51080 5868
rect 51132 5856 51138 5908
rect 53101 5899 53159 5905
rect 53101 5865 53113 5899
rect 53147 5896 53159 5899
rect 53374 5896 53380 5908
rect 53147 5868 53380 5896
rect 53147 5865 53159 5868
rect 53101 5859 53159 5865
rect 53374 5856 53380 5868
rect 53432 5896 53438 5908
rect 55214 5896 55220 5908
rect 53432 5868 55220 5896
rect 53432 5856 53438 5868
rect 55214 5856 55220 5868
rect 55272 5856 55278 5908
rect 56686 5856 56692 5908
rect 56744 5856 56750 5908
rect 56778 5856 56784 5908
rect 56836 5856 56842 5908
rect 58434 5856 58440 5908
rect 58492 5856 58498 5908
rect 50893 5831 50951 5837
rect 50893 5797 50905 5831
rect 50939 5828 50951 5831
rect 50939 5800 51074 5828
rect 50939 5797 50951 5800
rect 50893 5791 50951 5797
rect 48547 5732 48636 5760
rect 48547 5729 48559 5732
rect 48501 5723 48559 5729
rect 50246 5720 50252 5772
rect 50304 5720 50310 5772
rect 51046 5760 51074 5800
rect 51537 5763 51595 5769
rect 51537 5760 51549 5763
rect 51046 5732 51549 5760
rect 51537 5729 51549 5732
rect 51583 5729 51595 5763
rect 57698 5760 57704 5772
rect 51537 5723 51595 5729
rect 56336 5732 57704 5760
rect 39347 5664 39804 5692
rect 39853 5695 39911 5701
rect 39347 5661 39359 5664
rect 39301 5655 39359 5661
rect 39853 5661 39865 5695
rect 39899 5692 39911 5695
rect 40770 5692 40776 5704
rect 39899 5664 40776 5692
rect 39899 5661 39911 5664
rect 39853 5655 39911 5661
rect 28905 5627 28963 5633
rect 28905 5593 28917 5627
rect 28951 5624 28963 5627
rect 29270 5624 29276 5636
rect 28951 5596 29276 5624
rect 28951 5593 28963 5596
rect 28905 5587 28963 5593
rect 29270 5584 29276 5596
rect 29328 5584 29334 5636
rect 33137 5627 33195 5633
rect 33137 5593 33149 5627
rect 33183 5624 33195 5627
rect 34701 5627 34759 5633
rect 34701 5624 34713 5627
rect 33183 5596 34713 5624
rect 33183 5593 33195 5596
rect 33137 5587 33195 5593
rect 34701 5593 34713 5596
rect 34747 5593 34759 5627
rect 34701 5587 34759 5593
rect 36538 5584 36544 5636
rect 36596 5624 36602 5636
rect 37660 5624 37688 5655
rect 40770 5652 40776 5664
rect 40828 5692 40834 5704
rect 42705 5695 42763 5701
rect 40828 5664 41414 5692
rect 40828 5652 40834 5664
rect 36596 5596 37688 5624
rect 36596 5584 36602 5596
rect 37918 5584 37924 5636
rect 37976 5584 37982 5636
rect 39393 5627 39451 5633
rect 39393 5593 39405 5627
rect 39439 5624 39451 5627
rect 39758 5624 39764 5636
rect 39439 5596 39764 5624
rect 39439 5593 39451 5596
rect 39393 5587 39451 5593
rect 39758 5584 39764 5596
rect 39816 5584 39822 5636
rect 41386 5624 41414 5664
rect 42705 5661 42717 5695
rect 42751 5692 42763 5695
rect 43346 5692 43352 5704
rect 42751 5664 43352 5692
rect 42751 5661 42763 5664
rect 42705 5655 42763 5661
rect 43346 5652 43352 5664
rect 43404 5652 43410 5704
rect 47302 5652 47308 5704
rect 47360 5652 47366 5704
rect 48317 5695 48375 5701
rect 48317 5661 48329 5695
rect 48363 5692 48375 5695
rect 48866 5692 48872 5704
rect 48363 5664 48872 5692
rect 48363 5661 48375 5664
rect 48317 5655 48375 5661
rect 48866 5652 48872 5664
rect 48924 5652 48930 5704
rect 49694 5652 49700 5704
rect 49752 5701 49758 5704
rect 49752 5692 49764 5701
rect 49973 5695 50031 5701
rect 49752 5664 49797 5692
rect 49752 5655 49764 5664
rect 49973 5661 49985 5695
rect 50019 5692 50031 5695
rect 50154 5692 50160 5704
rect 50019 5664 50160 5692
rect 50019 5661 50031 5664
rect 49973 5655 50031 5661
rect 49752 5652 49758 5655
rect 50154 5652 50160 5664
rect 50212 5652 50218 5704
rect 50430 5652 50436 5704
rect 50488 5692 50494 5704
rect 50985 5695 51043 5701
rect 50985 5692 50997 5695
rect 50488 5664 50997 5692
rect 50488 5652 50494 5664
rect 50985 5661 50997 5664
rect 51031 5661 51043 5695
rect 50985 5655 51043 5661
rect 51721 5695 51779 5701
rect 51721 5661 51733 5695
rect 51767 5692 51779 5695
rect 52822 5692 52828 5704
rect 51767 5664 52828 5692
rect 51767 5661 51779 5664
rect 51721 5655 51779 5661
rect 52822 5652 52828 5664
rect 52880 5692 52886 5704
rect 54941 5695 54999 5701
rect 54941 5692 54953 5695
rect 52880 5664 54953 5692
rect 52880 5652 52886 5664
rect 54941 5661 54953 5664
rect 54987 5692 54999 5695
rect 55309 5695 55367 5701
rect 55309 5692 55321 5695
rect 54987 5664 55321 5692
rect 54987 5661 54999 5664
rect 54941 5655 54999 5661
rect 55309 5661 55321 5664
rect 55355 5692 55367 5695
rect 56336 5692 56364 5732
rect 57698 5720 57704 5732
rect 57756 5720 57762 5772
rect 55355 5664 56364 5692
rect 55355 5661 55367 5664
rect 55309 5655 55367 5661
rect 56686 5652 56692 5704
rect 56744 5692 56750 5704
rect 57333 5695 57391 5701
rect 57333 5692 57345 5695
rect 56744 5664 57345 5692
rect 56744 5652 56750 5664
rect 57333 5661 57345 5664
rect 57379 5661 57391 5695
rect 57333 5655 57391 5661
rect 58069 5695 58127 5701
rect 58069 5661 58081 5695
rect 58115 5661 58127 5695
rect 58069 5655 58127 5661
rect 44174 5624 44180 5636
rect 41386 5596 44180 5624
rect 44174 5584 44180 5596
rect 44232 5584 44238 5636
rect 45456 5627 45514 5633
rect 45456 5593 45468 5627
rect 45502 5624 45514 5627
rect 46014 5624 46020 5636
rect 45502 5596 46020 5624
rect 45502 5593 45514 5596
rect 45456 5587 45514 5593
rect 46014 5584 46020 5596
rect 46072 5584 46078 5636
rect 51988 5627 52046 5633
rect 51988 5593 52000 5627
rect 52034 5624 52046 5627
rect 52270 5624 52276 5636
rect 52034 5596 52276 5624
rect 52034 5593 52046 5596
rect 51988 5587 52046 5593
rect 52270 5584 52276 5596
rect 52328 5584 52334 5636
rect 52730 5584 52736 5636
rect 52788 5624 52794 5636
rect 53193 5627 53251 5633
rect 53193 5624 53205 5627
rect 52788 5596 53205 5624
rect 52788 5584 52794 5596
rect 53193 5593 53205 5596
rect 53239 5624 53251 5627
rect 54018 5624 54024 5636
rect 53239 5596 54024 5624
rect 53239 5593 53251 5596
rect 53193 5587 53251 5593
rect 54018 5584 54024 5596
rect 54076 5584 54082 5636
rect 55576 5627 55634 5633
rect 55576 5593 55588 5627
rect 55622 5624 55634 5627
rect 55674 5624 55680 5636
rect 55622 5596 55680 5624
rect 55622 5593 55634 5596
rect 55576 5587 55634 5593
rect 55674 5584 55680 5596
rect 55732 5584 55738 5636
rect 56502 5584 56508 5636
rect 56560 5624 56566 5636
rect 58084 5624 58112 5655
rect 58250 5652 58256 5704
rect 58308 5652 58314 5704
rect 56560 5596 58112 5624
rect 56560 5584 56566 5596
rect 28592 5528 28836 5556
rect 28592 5516 28598 5528
rect 28994 5516 29000 5568
rect 29052 5516 29058 5568
rect 29362 5516 29368 5568
rect 29420 5516 29426 5568
rect 30929 5559 30987 5565
rect 30929 5525 30941 5559
rect 30975 5556 30987 5559
rect 32674 5556 32680 5568
rect 30975 5528 32680 5556
rect 30975 5525 30987 5528
rect 30929 5519 30987 5525
rect 32674 5516 32680 5528
rect 32732 5516 32738 5568
rect 32858 5516 32864 5568
rect 32916 5556 32922 5568
rect 33229 5559 33287 5565
rect 33229 5556 33241 5559
rect 32916 5528 33241 5556
rect 32916 5516 32922 5528
rect 33229 5525 33241 5528
rect 33275 5525 33287 5559
rect 33229 5519 33287 5525
rect 33594 5516 33600 5568
rect 33652 5516 33658 5568
rect 37090 5516 37096 5568
rect 37148 5516 37154 5568
rect 38746 5516 38752 5568
rect 38804 5556 38810 5568
rect 38933 5559 38991 5565
rect 38933 5556 38945 5559
rect 38804 5528 38945 5556
rect 38804 5516 38810 5528
rect 38933 5525 38945 5528
rect 38979 5525 38991 5559
rect 38933 5519 38991 5525
rect 41138 5516 41144 5568
rect 41196 5556 41202 5568
rect 41782 5556 41788 5568
rect 41196 5528 41788 5556
rect 41196 5516 41202 5528
rect 41782 5516 41788 5528
rect 41840 5516 41846 5568
rect 41969 5559 42027 5565
rect 41969 5525 41981 5559
rect 42015 5556 42027 5559
rect 42150 5556 42156 5568
rect 42015 5528 42156 5556
rect 42015 5525 42027 5528
rect 41969 5519 42027 5525
rect 42150 5516 42156 5528
rect 42208 5516 42214 5568
rect 42702 5516 42708 5568
rect 42760 5556 42766 5568
rect 42797 5559 42855 5565
rect 42797 5556 42809 5559
rect 42760 5528 42809 5556
rect 42760 5516 42766 5528
rect 42797 5525 42809 5528
rect 42843 5525 42855 5559
rect 42797 5519 42855 5525
rect 43441 5559 43499 5565
rect 43441 5525 43453 5559
rect 43487 5556 43499 5559
rect 44818 5556 44824 5568
rect 43487 5528 44824 5556
rect 43487 5525 43499 5528
rect 43441 5519 43499 5525
rect 44818 5516 44824 5528
rect 44876 5516 44882 5568
rect 46661 5559 46719 5565
rect 46661 5525 46673 5559
rect 46707 5556 46719 5559
rect 47946 5556 47952 5568
rect 46707 5528 47952 5556
rect 46707 5525 46719 5528
rect 46661 5519 46719 5525
rect 47946 5516 47952 5528
rect 48004 5516 48010 5568
rect 49602 5516 49608 5568
rect 49660 5556 49666 5568
rect 50433 5559 50491 5565
rect 50433 5556 50445 5559
rect 49660 5528 50445 5556
rect 49660 5516 49666 5528
rect 50433 5525 50445 5528
rect 50479 5525 50491 5559
rect 50433 5519 50491 5525
rect 50525 5559 50583 5565
rect 50525 5525 50537 5559
rect 50571 5556 50583 5559
rect 51074 5556 51080 5568
rect 50571 5528 51080 5556
rect 50571 5525 50583 5528
rect 50525 5519 50583 5525
rect 51074 5516 51080 5528
rect 51132 5516 51138 5568
rect 57514 5516 57520 5568
rect 57572 5516 57578 5568
rect 1104 5466 59040 5488
rect 1104 5414 15394 5466
rect 15446 5414 15458 5466
rect 15510 5414 15522 5466
rect 15574 5414 15586 5466
rect 15638 5414 15650 5466
rect 15702 5414 29838 5466
rect 29890 5414 29902 5466
rect 29954 5414 29966 5466
rect 30018 5414 30030 5466
rect 30082 5414 30094 5466
rect 30146 5414 44282 5466
rect 44334 5414 44346 5466
rect 44398 5414 44410 5466
rect 44462 5414 44474 5466
rect 44526 5414 44538 5466
rect 44590 5414 58726 5466
rect 58778 5414 58790 5466
rect 58842 5414 58854 5466
rect 58906 5414 58918 5466
rect 58970 5414 58982 5466
rect 59034 5414 59040 5466
rect 1104 5392 59040 5414
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 4338 5352 4344 5364
rect 2740 5324 4344 5352
rect 2740 5312 2746 5324
rect 4338 5312 4344 5324
rect 4396 5352 4402 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 4396 5324 6101 5352
rect 4396 5312 4402 5324
rect 6089 5321 6101 5324
rect 6135 5352 6147 5355
rect 6362 5352 6368 5364
rect 6135 5324 6368 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7432 5324 7481 5352
rect 7432 5312 7438 5324
rect 7469 5321 7481 5324
rect 7515 5352 7527 5355
rect 7742 5352 7748 5364
rect 7515 5324 7748 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 10134 5352 10140 5364
rect 8588 5324 10140 5352
rect 3421 5287 3479 5293
rect 3421 5253 3433 5287
rect 3467 5284 3479 5287
rect 3510 5284 3516 5296
rect 3467 5256 3516 5284
rect 3467 5253 3479 5256
rect 3421 5247 3479 5253
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 4801 5287 4859 5293
rect 4801 5253 4813 5287
rect 4847 5284 4859 5287
rect 5166 5284 5172 5296
rect 4847 5256 5172 5284
rect 4847 5253 4859 5256
rect 4801 5247 4859 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 5626 5284 5632 5296
rect 5307 5256 5632 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 8588 5284 8616 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 11054 5352 11060 5364
rect 10735 5324 11060 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11204 5324 14044 5352
rect 11204 5312 11210 5324
rect 6656 5256 8616 5284
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 5353 5219 5411 5225
rect 2271 5188 3648 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 3510 5108 3516 5160
rect 3568 5108 3574 5160
rect 3620 5157 3648 5188
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5399 5188 6377 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5994 5148 6000 5160
rect 5491 5120 6000 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2958 5080 2964 5092
rect 1903 5052 2964 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3326 5080 3332 5092
rect 3099 5052 3332 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3620 5080 3648 5111
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6656 5080 6684 5256
rect 8662 5244 8668 5296
rect 8720 5293 8726 5296
rect 8720 5287 8743 5293
rect 8731 5253 8743 5287
rect 8720 5247 8743 5253
rect 8720 5244 8726 5247
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 8904 5256 9996 5284
rect 8904 5244 8910 5256
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7098 5216 7104 5228
rect 7055 5188 7104 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9048 5188 9689 5216
rect 9048 5080 9076 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 3620 5052 6684 5080
rect 8956 5052 9076 5080
rect 9968 5080 9996 5256
rect 11882 5244 11888 5296
rect 11940 5284 11946 5296
rect 13354 5284 13360 5296
rect 11940 5256 13360 5284
rect 11940 5244 11946 5256
rect 13354 5244 13360 5256
rect 13412 5244 13418 5296
rect 13572 5287 13630 5293
rect 13572 5253 13584 5287
rect 13618 5284 13630 5287
rect 13909 5287 13967 5293
rect 13909 5284 13921 5287
rect 13618 5256 13921 5284
rect 13618 5253 13630 5256
rect 13572 5247 13630 5253
rect 13909 5253 13921 5256
rect 13955 5253 13967 5287
rect 14016 5284 14044 5324
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14700 5324 14841 5352
rect 14700 5312 14706 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 19886 5352 19892 5364
rect 16172 5324 19892 5352
rect 16172 5312 16178 5324
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20625 5355 20683 5361
rect 20625 5321 20637 5355
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 20349 5287 20407 5293
rect 14016 5256 20300 5284
rect 13909 5247 13967 5253
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10597 5219 10655 5225
rect 10091 5188 10548 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10520 5148 10548 5188
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 10643 5188 11805 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16540 5176 16574 5216
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18012 5188 18429 5216
rect 18012 5176 18018 5188
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 19521 5219 19579 5225
rect 18463 5188 19472 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 11054 5148 11060 5160
rect 10520 5120 11060 5148
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 11698 5108 11704 5160
rect 11756 5108 11762 5160
rect 13814 5108 13820 5160
rect 13872 5108 13878 5160
rect 12066 5080 12072 5092
rect 9968 5052 12072 5080
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 4614 5012 4620 5024
rect 2915 4984 4620 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4893 5015 4951 5021
rect 4893 4981 4905 5015
rect 4939 5012 4951 5015
rect 4982 5012 4988 5024
rect 4939 4984 4988 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 7374 5012 7380 5024
rect 5224 4984 7380 5012
rect 5224 4972 5230 4984
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7561 5015 7619 5021
rect 7561 4981 7573 5015
rect 7607 5012 7619 5015
rect 7834 5012 7840 5024
rect 7607 4984 7840 5012
rect 7607 4981 7619 4984
rect 7561 4975 7619 4981
rect 7834 4972 7840 4984
rect 7892 5012 7898 5024
rect 8956 5012 8984 5052
rect 12066 5040 12072 5052
rect 12124 5080 12130 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 12124 5052 12572 5080
rect 12124 5040 12130 5052
rect 7892 4984 8984 5012
rect 7892 4972 7898 4984
rect 9030 4972 9036 5024
rect 9088 4972 9094 5024
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 12216 4984 12265 5012
rect 12216 4972 12222 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 12400 4984 12449 5012
rect 12400 4972 12406 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12544 5012 12572 5052
rect 13832 5052 15761 5080
rect 13832 5012 13860 5052
rect 15749 5049 15761 5052
rect 15795 5080 15807 5083
rect 16546 5080 16574 5176
rect 17218 5108 17224 5160
rect 17276 5108 17282 5160
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 19242 5108 19248 5160
rect 19300 5108 19306 5160
rect 19444 5148 19472 5188
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 19794 5216 19800 5228
rect 19567 5188 19800 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 20272 5216 20300 5256
rect 20349 5253 20361 5287
rect 20395 5284 20407 5287
rect 20640 5284 20668 5315
rect 21358 5312 21364 5364
rect 21416 5352 21422 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21416 5324 21557 5352
rect 21416 5312 21422 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 26697 5355 26755 5361
rect 21545 5315 21603 5321
rect 21652 5324 26648 5352
rect 21652 5284 21680 5324
rect 20395 5256 20668 5284
rect 20732 5256 21680 5284
rect 20395 5253 20407 5256
rect 20349 5247 20407 5253
rect 20732 5216 20760 5256
rect 22186 5244 22192 5296
rect 22244 5244 22250 5296
rect 23017 5287 23075 5293
rect 23017 5253 23029 5287
rect 23063 5284 23075 5287
rect 23934 5284 23940 5296
rect 23063 5256 23940 5284
rect 23063 5253 23075 5256
rect 23017 5247 23075 5253
rect 23934 5244 23940 5256
rect 23992 5244 23998 5296
rect 25332 5256 26556 5284
rect 20272 5188 20760 5216
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 22204 5216 22232 5244
rect 23109 5219 23167 5225
rect 21315 5188 22692 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 19705 5151 19763 5157
rect 19705 5148 19717 5151
rect 19444 5120 19717 5148
rect 19705 5117 19717 5120
rect 19751 5148 19763 5151
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19751 5120 19993 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 18966 5080 18972 5092
rect 15795 5052 16160 5080
rect 16546 5052 18972 5080
rect 15795 5049 15807 5052
rect 15749 5043 15807 5049
rect 16132 5024 16160 5052
rect 18966 5040 18972 5052
rect 19024 5080 19030 5092
rect 19426 5080 19432 5092
rect 19024 5052 19432 5080
rect 19024 5040 19030 5052
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 19996 5080 20024 5111
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 20824 5148 20852 5179
rect 20772 5120 20852 5148
rect 22557 5151 22615 5157
rect 20772 5108 20778 5120
rect 22557 5117 22569 5151
rect 22603 5117 22615 5151
rect 22664 5148 22692 5188
rect 23109 5185 23121 5219
rect 23155 5216 23167 5219
rect 23477 5219 23535 5225
rect 23477 5216 23489 5219
rect 23155 5188 23489 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 23477 5185 23489 5188
rect 23523 5185 23535 5219
rect 23477 5179 23535 5185
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24176 5188 24256 5216
rect 24176 5176 24182 5188
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 22664 5120 23213 5148
rect 22557 5111 22615 5117
rect 23201 5117 23213 5120
rect 23247 5117 23259 5151
rect 23201 5111 23259 5117
rect 21542 5080 21548 5092
rect 19996 5052 21548 5080
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 22572 5080 22600 5111
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 22572 5052 22661 5080
rect 22649 5049 22661 5052
rect 22695 5049 22707 5083
rect 24228 5080 24256 5188
rect 24854 5176 24860 5228
rect 24912 5216 24918 5228
rect 25332 5225 25360 5256
rect 25590 5225 25596 5228
rect 25317 5219 25375 5225
rect 25317 5216 25329 5219
rect 24912 5188 25329 5216
rect 24912 5176 24918 5188
rect 25317 5185 25329 5188
rect 25363 5185 25375 5219
rect 25584 5216 25596 5225
rect 25551 5188 25596 5216
rect 25317 5179 25375 5185
rect 25584 5179 25596 5188
rect 25590 5176 25596 5179
rect 25648 5176 25654 5228
rect 24670 5108 24676 5160
rect 24728 5148 24734 5160
rect 24765 5151 24823 5157
rect 24765 5148 24777 5151
rect 24728 5120 24777 5148
rect 24728 5108 24734 5120
rect 24765 5117 24777 5120
rect 24811 5117 24823 5151
rect 26528 5148 26556 5256
rect 26620 5216 26648 5324
rect 26697 5321 26709 5355
rect 26743 5352 26755 5355
rect 26970 5352 26976 5364
rect 26743 5324 26976 5352
rect 26743 5321 26755 5324
rect 26697 5315 26755 5321
rect 26970 5312 26976 5324
rect 27028 5312 27034 5364
rect 27982 5312 27988 5364
rect 28040 5312 28046 5364
rect 29270 5312 29276 5364
rect 29328 5352 29334 5364
rect 29549 5355 29607 5361
rect 29549 5352 29561 5355
rect 29328 5324 29561 5352
rect 29328 5312 29334 5324
rect 29549 5321 29561 5324
rect 29595 5321 29607 5355
rect 29549 5315 29607 5321
rect 29638 5312 29644 5364
rect 29696 5312 29702 5364
rect 30282 5312 30288 5364
rect 30340 5312 30346 5364
rect 30929 5355 30987 5361
rect 30929 5321 30941 5355
rect 30975 5352 30987 5355
rect 31110 5352 31116 5364
rect 30975 5324 31116 5352
rect 30975 5321 30987 5324
rect 30929 5315 30987 5321
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 31294 5312 31300 5364
rect 31352 5312 31358 5364
rect 32122 5312 32128 5364
rect 32180 5352 32186 5364
rect 35253 5355 35311 5361
rect 35253 5352 35265 5355
rect 32180 5324 35265 5352
rect 32180 5312 32186 5324
rect 35253 5321 35265 5324
rect 35299 5321 35311 5355
rect 35253 5315 35311 5321
rect 35713 5355 35771 5361
rect 35713 5321 35725 5355
rect 35759 5352 35771 5355
rect 35986 5352 35992 5364
rect 35759 5324 35992 5352
rect 35759 5321 35771 5324
rect 35713 5315 35771 5321
rect 27338 5244 27344 5296
rect 27396 5284 27402 5296
rect 29457 5287 29515 5293
rect 27396 5256 29040 5284
rect 27396 5244 27402 5256
rect 26620 5188 27752 5216
rect 27157 5151 27215 5157
rect 27157 5148 27169 5151
rect 26528 5120 27169 5148
rect 24765 5111 24823 5117
rect 27157 5117 27169 5120
rect 27203 5148 27215 5151
rect 27525 5151 27583 5157
rect 27525 5148 27537 5151
rect 27203 5120 27537 5148
rect 27203 5117 27215 5120
rect 27157 5111 27215 5117
rect 27525 5117 27537 5120
rect 27571 5148 27583 5151
rect 27614 5148 27620 5160
rect 27571 5120 27620 5148
rect 27571 5117 27583 5120
rect 27525 5111 27583 5117
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 24228 5052 25360 5080
rect 22649 5043 22707 5049
rect 25332 5024 25360 5052
rect 27724 5024 27752 5188
rect 28629 5083 28687 5089
rect 28629 5049 28641 5083
rect 28675 5080 28687 5083
rect 28675 5052 28856 5080
rect 28675 5049 28687 5052
rect 28629 5043 28687 5049
rect 28828 5024 28856 5052
rect 12544 4984 13860 5012
rect 15381 5015 15439 5021
rect 12437 4975 12495 4981
rect 15381 4981 15393 5015
rect 15427 5012 15439 5015
rect 15930 5012 15936 5024
rect 15427 4984 15936 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 16114 4972 16120 5024
rect 16172 4972 16178 5024
rect 16666 4972 16672 5024
rect 16724 4972 16730 5024
rect 17494 4972 17500 5024
rect 17552 4972 17558 5024
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18564 4984 18613 5012
rect 18564 4972 18570 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 19334 4972 19340 5024
rect 19392 4972 19398 5024
rect 20254 4972 20260 5024
rect 20312 4972 20318 5024
rect 21910 4972 21916 5024
rect 21968 4972 21974 5024
rect 24210 4972 24216 5024
rect 24268 4972 24274 5024
rect 25222 4972 25228 5024
rect 25280 4972 25286 5024
rect 25314 4972 25320 5024
rect 25372 4972 25378 5024
rect 27706 4972 27712 5024
rect 27764 4972 27770 5024
rect 27798 4972 27804 5024
rect 27856 5012 27862 5024
rect 28353 5015 28411 5021
rect 28353 5012 28365 5015
rect 27856 4984 28365 5012
rect 27856 4972 27862 4984
rect 28353 4981 28365 4984
rect 28399 5012 28411 5015
rect 28718 5012 28724 5024
rect 28399 4984 28724 5012
rect 28399 4981 28411 4984
rect 28353 4975 28411 4981
rect 28718 4972 28724 4984
rect 28776 4972 28782 5024
rect 28810 4972 28816 5024
rect 28868 4972 28874 5024
rect 29012 5012 29040 5256
rect 29457 5253 29469 5287
rect 29503 5284 29515 5287
rect 29656 5284 29684 5312
rect 29503 5256 29684 5284
rect 30300 5284 30328 5312
rect 32582 5284 32588 5296
rect 30300 5256 32588 5284
rect 29503 5253 29515 5256
rect 29457 5247 29515 5253
rect 32582 5244 32588 5256
rect 32640 5244 32646 5296
rect 32769 5287 32827 5293
rect 32769 5253 32781 5287
rect 32815 5284 32827 5287
rect 33965 5287 34023 5293
rect 33965 5284 33977 5287
rect 32815 5256 33977 5284
rect 32815 5253 32827 5256
rect 32769 5247 32827 5253
rect 33965 5253 33977 5256
rect 34011 5253 34023 5287
rect 33965 5247 34023 5253
rect 34882 5244 34888 5296
rect 34940 5244 34946 5296
rect 35268 5284 35296 5315
rect 35986 5312 35992 5324
rect 36044 5312 36050 5364
rect 36078 5312 36084 5364
rect 36136 5312 36142 5364
rect 36173 5355 36231 5361
rect 36173 5321 36185 5355
rect 36219 5352 36231 5355
rect 37090 5352 37096 5364
rect 36219 5324 37096 5352
rect 36219 5321 36231 5324
rect 36173 5315 36231 5321
rect 37090 5312 37096 5324
rect 37148 5312 37154 5364
rect 37642 5312 37648 5364
rect 37700 5312 37706 5364
rect 40494 5312 40500 5364
rect 40552 5312 40558 5364
rect 41782 5312 41788 5364
rect 41840 5352 41846 5364
rect 42153 5355 42211 5361
rect 42153 5352 42165 5355
rect 41840 5324 42165 5352
rect 41840 5312 41846 5324
rect 42153 5321 42165 5324
rect 42199 5352 42211 5355
rect 43533 5355 43591 5361
rect 43533 5352 43545 5355
rect 42199 5324 43545 5352
rect 42199 5321 42211 5324
rect 42153 5315 42211 5321
rect 43533 5321 43545 5324
rect 43579 5352 43591 5355
rect 43901 5355 43959 5361
rect 43901 5352 43913 5355
rect 43579 5324 43913 5352
rect 43579 5321 43591 5324
rect 43533 5315 43591 5321
rect 43901 5321 43913 5324
rect 43947 5352 43959 5355
rect 44174 5352 44180 5364
rect 43947 5324 44180 5352
rect 43947 5321 43959 5324
rect 43901 5315 43959 5321
rect 44174 5312 44180 5324
rect 44232 5352 44238 5364
rect 44637 5355 44695 5361
rect 44637 5352 44649 5355
rect 44232 5324 44649 5352
rect 44232 5312 44238 5324
rect 44637 5321 44649 5324
rect 44683 5352 44695 5355
rect 45186 5352 45192 5364
rect 44683 5324 45192 5352
rect 44683 5321 44695 5324
rect 44637 5315 44695 5321
rect 45186 5312 45192 5324
rect 45244 5312 45250 5364
rect 45646 5312 45652 5364
rect 45704 5312 45710 5364
rect 46017 5355 46075 5361
rect 46017 5321 46029 5355
rect 46063 5352 46075 5355
rect 46566 5352 46572 5364
rect 46063 5324 46572 5352
rect 46063 5321 46075 5324
rect 46017 5315 46075 5321
rect 46566 5312 46572 5324
rect 46624 5312 46630 5364
rect 48516 5324 50752 5352
rect 36446 5284 36452 5296
rect 35268 5256 36452 5284
rect 36446 5244 36452 5256
rect 36504 5244 36510 5296
rect 36722 5244 36728 5296
rect 36780 5244 36786 5296
rect 38841 5287 38899 5293
rect 38841 5253 38853 5287
rect 38887 5284 38899 5287
rect 39178 5287 39236 5293
rect 39178 5284 39190 5287
rect 38887 5256 39190 5284
rect 38887 5253 38899 5256
rect 38841 5247 38899 5253
rect 39178 5253 39190 5256
rect 39224 5253 39236 5287
rect 39178 5247 39236 5253
rect 29362 5176 29368 5228
rect 29420 5216 29426 5228
rect 30285 5219 30343 5225
rect 30285 5216 30297 5219
rect 29420 5188 30297 5216
rect 29420 5176 29426 5188
rect 30285 5185 30297 5188
rect 30331 5185 30343 5219
rect 30285 5179 30343 5185
rect 31294 5176 31300 5228
rect 31352 5216 31358 5228
rect 32122 5216 32128 5228
rect 31352 5188 32128 5216
rect 31352 5176 31358 5188
rect 32122 5176 32128 5188
rect 32180 5176 32186 5228
rect 32677 5219 32735 5225
rect 32677 5216 32689 5219
rect 32416 5188 32689 5216
rect 32416 5160 32444 5188
rect 32677 5185 32689 5188
rect 32723 5216 32735 5219
rect 32858 5216 32864 5228
rect 32723 5188 32864 5216
rect 32723 5185 32735 5188
rect 32677 5179 32735 5185
rect 32858 5176 32864 5188
rect 32916 5176 32922 5228
rect 33226 5176 33232 5228
rect 33284 5176 33290 5228
rect 33594 5176 33600 5228
rect 33652 5216 33658 5228
rect 33781 5219 33839 5225
rect 33781 5216 33793 5219
rect 33652 5188 33793 5216
rect 33652 5176 33658 5188
rect 33781 5185 33793 5188
rect 33827 5185 33839 5219
rect 33781 5179 33839 5185
rect 33870 5176 33876 5228
rect 33928 5216 33934 5228
rect 34517 5219 34575 5225
rect 34517 5216 34529 5219
rect 33928 5188 34529 5216
rect 33928 5176 33934 5188
rect 34517 5185 34529 5188
rect 34563 5185 34575 5219
rect 34900 5216 34928 5244
rect 35802 5216 35808 5228
rect 34900 5188 35808 5216
rect 34517 5179 34575 5185
rect 35802 5176 35808 5188
rect 35860 5176 35866 5228
rect 36170 5176 36176 5228
rect 36228 5216 36234 5228
rect 36228 5188 36308 5216
rect 36228 5176 36234 5188
rect 30190 5108 30196 5160
rect 30248 5108 30254 5160
rect 31386 5108 31392 5160
rect 31444 5148 31450 5160
rect 31665 5151 31723 5157
rect 31665 5148 31677 5151
rect 31444 5120 31677 5148
rect 31444 5108 31450 5120
rect 31665 5117 31677 5120
rect 31711 5148 31723 5151
rect 32306 5148 32312 5160
rect 31711 5120 32312 5148
rect 31711 5117 31723 5120
rect 31665 5111 31723 5117
rect 32306 5108 32312 5120
rect 32364 5108 32370 5160
rect 32398 5108 32404 5160
rect 32456 5108 32462 5160
rect 32585 5151 32643 5157
rect 32585 5117 32597 5151
rect 32631 5148 32643 5151
rect 34422 5148 34428 5160
rect 32631 5120 34428 5148
rect 32631 5117 32643 5120
rect 32585 5111 32643 5117
rect 29089 5083 29147 5089
rect 29089 5049 29101 5083
rect 29135 5080 29147 5083
rect 32600 5080 32628 5111
rect 34422 5108 34428 5120
rect 34480 5108 34486 5160
rect 36280 5157 36308 5188
rect 38654 5176 38660 5228
rect 38712 5216 38718 5228
rect 38933 5219 38991 5225
rect 38933 5216 38945 5219
rect 38712 5188 38945 5216
rect 38712 5176 38718 5188
rect 38933 5185 38945 5188
rect 38979 5185 38991 5219
rect 40512 5216 40540 5312
rect 42794 5244 42800 5296
rect 42852 5244 42858 5296
rect 47486 5284 47492 5296
rect 45296 5256 47492 5284
rect 41230 5216 41236 5228
rect 40512 5188 41236 5216
rect 38933 5179 38991 5185
rect 41230 5176 41236 5188
rect 41288 5216 41294 5228
rect 42610 5216 42616 5228
rect 41288 5188 42616 5216
rect 41288 5176 41294 5188
rect 42610 5176 42616 5188
rect 42668 5216 42674 5228
rect 44177 5219 44235 5225
rect 44177 5216 44189 5219
rect 42668 5188 44189 5216
rect 42668 5176 42674 5188
rect 44177 5185 44189 5188
rect 44223 5185 44235 5219
rect 44177 5179 44235 5185
rect 36265 5151 36323 5157
rect 36265 5117 36277 5151
rect 36311 5117 36323 5151
rect 36265 5111 36323 5117
rect 37734 5108 37740 5160
rect 37792 5108 37798 5160
rect 37921 5151 37979 5157
rect 37921 5117 37933 5151
rect 37967 5148 37979 5151
rect 38289 5151 38347 5157
rect 37967 5120 38056 5148
rect 37967 5117 37979 5120
rect 37921 5111 37979 5117
rect 29135 5052 32628 5080
rect 33137 5083 33195 5089
rect 29135 5049 29147 5052
rect 29089 5043 29147 5049
rect 33137 5049 33149 5083
rect 33183 5080 33195 5083
rect 33502 5080 33508 5092
rect 33183 5052 33508 5080
rect 33183 5049 33195 5052
rect 33137 5043 33195 5049
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 33594 5040 33600 5092
rect 33652 5080 33658 5092
rect 33778 5080 33784 5092
rect 33652 5052 33784 5080
rect 33652 5040 33658 5052
rect 33778 5040 33784 5052
rect 33836 5080 33842 5092
rect 38028 5080 38056 5120
rect 38289 5117 38301 5151
rect 38335 5148 38347 5151
rect 38746 5148 38752 5160
rect 38335 5120 38752 5148
rect 38335 5117 38347 5120
rect 38289 5111 38347 5117
rect 38746 5108 38752 5120
rect 38804 5108 38810 5160
rect 39960 5120 41000 5148
rect 33836 5052 38056 5080
rect 33836 5040 33842 5052
rect 38028 5024 38056 5052
rect 34606 5012 34612 5024
rect 29012 4984 34612 5012
rect 34606 4972 34612 4984
rect 34664 4972 34670 5024
rect 35802 4972 35808 5024
rect 35860 5012 35866 5024
rect 36906 5012 36912 5024
rect 35860 4984 36912 5012
rect 35860 4972 35866 4984
rect 36906 4972 36912 4984
rect 36964 4972 36970 5024
rect 37277 5015 37335 5021
rect 37277 4981 37289 5015
rect 37323 5012 37335 5015
rect 37550 5012 37556 5024
rect 37323 4984 37556 5012
rect 37323 4981 37335 4984
rect 37277 4975 37335 4981
rect 37550 4972 37556 4984
rect 37608 4972 37614 5024
rect 38010 4972 38016 5024
rect 38068 5012 38074 5024
rect 39960 5012 39988 5120
rect 40313 5083 40371 5089
rect 40313 5049 40325 5083
rect 40359 5080 40371 5083
rect 40862 5080 40868 5092
rect 40359 5052 40868 5080
rect 40359 5049 40371 5052
rect 40313 5043 40371 5049
rect 40862 5040 40868 5052
rect 40920 5040 40926 5092
rect 40972 5080 41000 5120
rect 41046 5108 41052 5160
rect 41104 5108 41110 5160
rect 42521 5151 42579 5157
rect 42521 5117 42533 5151
rect 42567 5117 42579 5151
rect 42521 5111 42579 5117
rect 41417 5083 41475 5089
rect 41417 5080 41429 5083
rect 40972 5052 41429 5080
rect 41417 5049 41429 5052
rect 41463 5080 41475 5083
rect 42536 5080 42564 5111
rect 42702 5108 42708 5160
rect 42760 5108 42766 5160
rect 45002 5080 45008 5092
rect 41463 5052 45008 5080
rect 41463 5049 41475 5052
rect 41417 5043 41475 5049
rect 45002 5040 45008 5052
rect 45060 5080 45066 5092
rect 45296 5089 45324 5256
rect 47486 5244 47492 5256
rect 47544 5244 47550 5296
rect 46845 5219 46903 5225
rect 46845 5216 46857 5219
rect 46124 5188 46857 5216
rect 46124 5157 46152 5188
rect 46845 5185 46857 5188
rect 46891 5185 46903 5219
rect 46845 5179 46903 5185
rect 46937 5219 46995 5225
rect 46937 5185 46949 5219
rect 46983 5216 46995 5219
rect 47581 5219 47639 5225
rect 47581 5216 47593 5219
rect 46983 5188 47593 5216
rect 46983 5185 46995 5188
rect 46937 5179 46995 5185
rect 47581 5185 47593 5188
rect 47627 5185 47639 5219
rect 47581 5179 47639 5185
rect 47762 5176 47768 5228
rect 47820 5216 47826 5228
rect 48133 5219 48191 5225
rect 48133 5216 48145 5219
rect 47820 5188 48145 5216
rect 47820 5176 47826 5188
rect 48133 5185 48145 5188
rect 48179 5185 48191 5219
rect 48133 5179 48191 5185
rect 46109 5151 46167 5157
rect 46109 5117 46121 5151
rect 46155 5117 46167 5151
rect 46109 5111 46167 5117
rect 45281 5083 45339 5089
rect 45281 5080 45293 5083
rect 45060 5052 45293 5080
rect 45060 5040 45066 5052
rect 45281 5049 45293 5052
rect 45327 5049 45339 5083
rect 45281 5043 45339 5049
rect 38068 4984 39988 5012
rect 40405 5015 40463 5021
rect 38068 4972 38074 4984
rect 40405 4981 40417 5015
rect 40451 5012 40463 5015
rect 40494 5012 40500 5024
rect 40451 4984 40500 5012
rect 40451 4981 40463 4984
rect 40405 4975 40463 4981
rect 40494 4972 40500 4984
rect 40552 4972 40558 5024
rect 40880 5012 40908 5040
rect 41322 5012 41328 5024
rect 40880 4984 41328 5012
rect 41322 4972 41328 4984
rect 41380 4972 41386 5024
rect 41785 5015 41843 5021
rect 41785 4981 41797 5015
rect 41831 5012 41843 5015
rect 42150 5012 42156 5024
rect 41831 4984 42156 5012
rect 41831 4981 41843 4984
rect 41785 4975 41843 4981
rect 42150 4972 42156 4984
rect 42208 4972 42214 5024
rect 43165 5015 43223 5021
rect 43165 4981 43177 5015
rect 43211 5012 43223 5015
rect 43530 5012 43536 5024
rect 43211 4984 43536 5012
rect 43211 4981 43223 4984
rect 43165 4975 43223 4981
rect 43530 4972 43536 4984
rect 43588 4972 43594 5024
rect 44913 5015 44971 5021
rect 44913 4981 44925 5015
rect 44959 5012 44971 5015
rect 45370 5012 45376 5024
rect 44959 4984 45376 5012
rect 44959 4981 44971 4984
rect 44913 4975 44971 4981
rect 45370 4972 45376 4984
rect 45428 4972 45434 5024
rect 46124 5012 46152 5111
rect 46198 5108 46204 5160
rect 46256 5108 46262 5160
rect 47121 5151 47179 5157
rect 47121 5117 47133 5151
rect 47167 5148 47179 5151
rect 47670 5148 47676 5160
rect 47167 5120 47676 5148
rect 47167 5117 47179 5120
rect 47121 5111 47179 5117
rect 47670 5108 47676 5120
rect 47728 5108 47734 5160
rect 46216 5080 46244 5108
rect 48516 5089 48544 5324
rect 50004 5287 50062 5293
rect 50004 5253 50016 5287
rect 50050 5284 50062 5287
rect 50430 5284 50436 5296
rect 50050 5256 50436 5284
rect 50050 5253 50062 5256
rect 50004 5247 50062 5253
rect 50430 5244 50436 5256
rect 50488 5244 50494 5296
rect 50724 5284 50752 5324
rect 51074 5312 51080 5364
rect 51132 5312 51138 5364
rect 52546 5312 52552 5364
rect 52604 5352 52610 5364
rect 52733 5355 52791 5361
rect 52733 5352 52745 5355
rect 52604 5324 52745 5352
rect 52604 5312 52610 5324
rect 52733 5321 52745 5324
rect 52779 5321 52791 5355
rect 52733 5315 52791 5321
rect 54018 5312 54024 5364
rect 54076 5312 54082 5364
rect 54938 5312 54944 5364
rect 54996 5312 55002 5364
rect 55674 5312 55680 5364
rect 55732 5312 55738 5364
rect 56873 5355 56931 5361
rect 56873 5321 56885 5355
rect 56919 5352 56931 5355
rect 57514 5352 57520 5364
rect 56919 5324 57520 5352
rect 56919 5321 56931 5324
rect 56873 5315 56931 5321
rect 57514 5312 57520 5324
rect 57572 5312 57578 5364
rect 57606 5312 57612 5364
rect 57664 5312 57670 5364
rect 52638 5284 52644 5296
rect 50724 5256 52644 5284
rect 52638 5244 52644 5256
rect 52696 5244 52702 5296
rect 53098 5244 53104 5296
rect 53156 5284 53162 5296
rect 54297 5287 54355 5293
rect 54297 5284 54309 5287
rect 53156 5256 54309 5284
rect 53156 5244 53162 5256
rect 54297 5253 54309 5256
rect 54343 5284 54355 5287
rect 55217 5287 55275 5293
rect 54343 5256 54800 5284
rect 54343 5253 54355 5256
rect 54297 5247 54355 5253
rect 50154 5176 50160 5228
rect 50212 5216 50218 5228
rect 50249 5219 50307 5225
rect 50249 5216 50261 5219
rect 50212 5188 50261 5216
rect 50212 5176 50218 5188
rect 50249 5185 50261 5188
rect 50295 5216 50307 5219
rect 50525 5219 50583 5225
rect 50525 5216 50537 5219
rect 50295 5188 50537 5216
rect 50295 5185 50307 5188
rect 50249 5179 50307 5185
rect 50525 5185 50537 5188
rect 50571 5185 50583 5219
rect 50525 5179 50583 5185
rect 50890 5176 50896 5228
rect 50948 5176 50954 5228
rect 53374 5176 53380 5228
rect 53432 5176 53438 5228
rect 53561 5219 53619 5225
rect 53561 5185 53573 5219
rect 53607 5185 53619 5219
rect 53561 5179 53619 5185
rect 54481 5219 54539 5225
rect 54481 5185 54493 5219
rect 54527 5185 54539 5219
rect 54772 5216 54800 5256
rect 55217 5253 55229 5287
rect 55263 5284 55275 5287
rect 57330 5284 57336 5296
rect 55263 5256 57336 5284
rect 55263 5253 55275 5256
rect 55217 5247 55275 5253
rect 57330 5244 57336 5256
rect 57388 5244 57394 5296
rect 55585 5219 55643 5225
rect 54772 5188 55352 5216
rect 54481 5179 54539 5185
rect 50338 5108 50344 5160
rect 50396 5148 50402 5160
rect 50709 5151 50767 5157
rect 50709 5148 50721 5151
rect 50396 5120 50721 5148
rect 50396 5108 50402 5120
rect 50709 5117 50721 5120
rect 50755 5117 50767 5151
rect 51629 5151 51687 5157
rect 51629 5148 51641 5151
rect 50709 5111 50767 5117
rect 51046 5120 51641 5148
rect 48501 5083 48559 5089
rect 48501 5080 48513 5083
rect 46216 5052 48513 5080
rect 48501 5049 48513 5052
rect 48547 5049 48559 5083
rect 51046 5080 51074 5120
rect 51629 5117 51641 5120
rect 51675 5117 51687 5151
rect 51629 5111 51687 5117
rect 53006 5108 53012 5160
rect 53064 5148 53070 5160
rect 53576 5148 53604 5179
rect 53064 5120 53604 5148
rect 53064 5108 53070 5120
rect 48501 5043 48559 5049
rect 50264 5052 51074 5080
rect 54496 5080 54524 5179
rect 55214 5080 55220 5092
rect 54496 5052 55220 5080
rect 46198 5012 46204 5024
rect 46124 4984 46204 5012
rect 46198 4972 46204 4984
rect 46256 4972 46262 5024
rect 46474 4972 46480 5024
rect 46532 4972 46538 5024
rect 48866 4972 48872 5024
rect 48924 5012 48930 5024
rect 50264 5012 50292 5052
rect 55214 5040 55220 5052
rect 55272 5040 55278 5092
rect 55324 5080 55352 5188
rect 55585 5185 55597 5219
rect 55631 5185 55643 5219
rect 55585 5179 55643 5185
rect 55600 5148 55628 5179
rect 55950 5176 55956 5228
rect 56008 5216 56014 5228
rect 56229 5219 56287 5225
rect 56229 5216 56241 5219
rect 56008 5188 56241 5216
rect 56008 5176 56014 5188
rect 56229 5185 56241 5188
rect 56275 5185 56287 5219
rect 56229 5179 56287 5185
rect 56962 5176 56968 5228
rect 57020 5176 57026 5228
rect 57146 5176 57152 5228
rect 57204 5216 57210 5228
rect 57425 5219 57483 5225
rect 57425 5216 57437 5219
rect 57204 5188 57437 5216
rect 57204 5176 57210 5188
rect 57425 5185 57437 5188
rect 57471 5185 57483 5219
rect 57425 5179 57483 5185
rect 56134 5148 56140 5160
rect 55600 5120 56140 5148
rect 56134 5108 56140 5120
rect 56192 5108 56198 5160
rect 56594 5108 56600 5160
rect 56652 5148 56658 5160
rect 56689 5151 56747 5157
rect 56689 5148 56701 5151
rect 56652 5120 56701 5148
rect 56652 5108 56658 5120
rect 56689 5117 56701 5120
rect 56735 5117 56747 5151
rect 56689 5111 56747 5117
rect 56980 5080 57008 5176
rect 58437 5151 58495 5157
rect 58437 5117 58449 5151
rect 58483 5117 58495 5151
rect 58437 5111 58495 5117
rect 55324 5052 57008 5080
rect 57333 5083 57391 5089
rect 57333 5049 57345 5083
rect 57379 5080 57391 5083
rect 58452 5080 58480 5111
rect 57379 5052 58480 5080
rect 57379 5049 57391 5052
rect 57333 5043 57391 5049
rect 48924 4984 50292 5012
rect 48924 4972 48930 4984
rect 51166 4972 51172 5024
rect 51224 5012 51230 5024
rect 51997 5015 52055 5021
rect 51997 5012 52009 5015
rect 51224 4984 52009 5012
rect 51224 4972 51230 4984
rect 51997 4981 52009 4984
rect 52043 4981 52055 5015
rect 51997 4975 52055 4981
rect 52457 5015 52515 5021
rect 52457 4981 52469 5015
rect 52503 5012 52515 5015
rect 52546 5012 52552 5024
rect 52503 4984 52552 5012
rect 52503 4981 52515 4984
rect 52457 4975 52515 4981
rect 52546 4972 52552 4984
rect 52604 4972 52610 5024
rect 53742 4972 53748 5024
rect 53800 4972 53806 5024
rect 53834 4972 53840 5024
rect 53892 5012 53898 5024
rect 55125 5015 55183 5021
rect 55125 5012 55137 5015
rect 53892 4984 55137 5012
rect 53892 4972 53898 4984
rect 55125 4981 55137 4984
rect 55171 4981 55183 5015
rect 55125 4975 55183 4981
rect 55398 4972 55404 5024
rect 55456 4972 55462 5024
rect 57790 4972 57796 5024
rect 57848 5012 57854 5024
rect 57885 5015 57943 5021
rect 57885 5012 57897 5015
rect 57848 4984 57897 5012
rect 57848 4972 57854 4984
rect 57885 4981 57897 4984
rect 57931 4981 57943 5015
rect 57885 4975 57943 4981
rect 1104 4922 58880 4944
rect 1104 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 22616 4922
rect 22668 4870 22680 4922
rect 22732 4870 22744 4922
rect 22796 4870 22808 4922
rect 22860 4870 22872 4922
rect 22924 4870 37060 4922
rect 37112 4870 37124 4922
rect 37176 4870 37188 4922
rect 37240 4870 37252 4922
rect 37304 4870 37316 4922
rect 37368 4870 51504 4922
rect 51556 4870 51568 4922
rect 51620 4870 51632 4922
rect 51684 4870 51696 4922
rect 51748 4870 51760 4922
rect 51812 4870 58880 4922
rect 1104 4848 58880 4870
rect 1762 4768 1768 4820
rect 1820 4768 1826 4820
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 2648 4780 2774 4808
rect 2648 4768 2654 4780
rect 2746 4740 2774 4780
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 6086 4808 6092 4820
rect 4672 4780 6092 4808
rect 4672 4768 4678 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6178 4768 6184 4820
rect 6236 4768 6242 4820
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6420 4780 7205 4808
rect 6420 4768 6426 4780
rect 7193 4777 7205 4780
rect 7239 4808 7251 4811
rect 8938 4808 8944 4820
rect 7239 4780 8944 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9398 4808 9404 4820
rect 9355 4780 9404 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9824 4780 9965 4808
rect 9824 4768 9830 4780
rect 9953 4777 9965 4780
rect 9999 4808 10011 4811
rect 9999 4780 13400 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 4982 4740 4988 4752
rect 2746 4712 4988 4740
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 5997 4743 6055 4749
rect 5997 4709 6009 4743
rect 6043 4740 6055 4743
rect 6196 4740 6224 4768
rect 6043 4712 6224 4740
rect 6733 4743 6791 4749
rect 6043 4709 6055 4712
rect 5997 4703 6055 4709
rect 6733 4709 6745 4743
rect 6779 4740 6791 4743
rect 8294 4740 8300 4752
rect 6779 4712 8300 4740
rect 6779 4709 6791 4712
rect 6733 4703 6791 4709
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 6012 4672 6040 4703
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8956 4740 8984 4768
rect 9585 4743 9643 4749
rect 9585 4740 9597 4743
rect 8956 4712 9597 4740
rect 9585 4709 9597 4712
rect 9631 4740 9643 4743
rect 9674 4740 9680 4752
rect 9631 4712 9680 4740
rect 9631 4709 9643 4712
rect 9585 4703 9643 4709
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 7742 4672 7748 4684
rect 3292 4644 6040 4672
rect 7116 4644 7748 4672
rect 3292 4632 3298 4644
rect 7116 4616 7144 4644
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 8754 4672 8760 4684
rect 8711 4644 8760 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9030 4632 9036 4684
rect 9088 4632 9094 4684
rect 2866 4564 2872 4616
rect 2924 4564 2930 4616
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3142 4604 3148 4616
rect 3099 4576 3148 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4672 4576 4905 4604
rect 4672 4564 4678 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 5902 4604 5908 4616
rect 5767 4576 5908 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6546 4564 6552 4616
rect 6604 4564 6610 4616
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 8389 4607 8447 4613
rect 7607 4576 7696 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 2133 4539 2191 4545
rect 2133 4505 2145 4539
rect 2179 4536 2191 4539
rect 5166 4536 5172 4548
rect 2179 4508 5172 4536
rect 2179 4505 2191 4508
rect 2133 4499 2191 4505
rect 5166 4496 5172 4508
rect 5224 4496 5230 4548
rect 2222 4428 2228 4480
rect 2280 4428 2286 4480
rect 3602 4428 3608 4480
rect 3660 4428 3666 4480
rect 4246 4428 4252 4480
rect 4304 4428 4310 4480
rect 4338 4428 4344 4480
rect 4396 4428 4402 4480
rect 5074 4428 5080 4480
rect 5132 4428 5138 4480
rect 7374 4428 7380 4480
rect 7432 4428 7438 4480
rect 7668 4468 7696 4576
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 9048 4604 9076 4632
rect 8435 4576 9076 4604
rect 9692 4604 9720 4700
rect 10502 4604 10508 4616
rect 9692 4576 10508 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 10502 4564 10508 4576
rect 10560 4604 10566 4616
rect 13372 4613 13400 4780
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16080 4780 18644 4808
rect 16080 4768 16086 4780
rect 14829 4743 14887 4749
rect 14829 4709 14841 4743
rect 14875 4740 14887 4743
rect 15194 4740 15200 4752
rect 14875 4712 15200 4740
rect 14875 4709 14887 4712
rect 14829 4703 14887 4709
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 17497 4743 17555 4749
rect 17497 4709 17509 4743
rect 17543 4709 17555 4743
rect 18616 4740 18644 4780
rect 19242 4768 19248 4820
rect 19300 4768 19306 4820
rect 20070 4768 20076 4820
rect 20128 4768 20134 4820
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 21821 4811 21879 4817
rect 21821 4808 21833 4811
rect 20496 4780 21833 4808
rect 20496 4768 20502 4780
rect 21821 4777 21833 4780
rect 21867 4777 21879 4811
rect 21821 4771 21879 4777
rect 23385 4811 23443 4817
rect 23385 4777 23397 4811
rect 23431 4808 23443 4811
rect 24118 4808 24124 4820
rect 23431 4780 24124 4808
rect 23431 4777 23443 4780
rect 23385 4771 23443 4777
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24210 4768 24216 4820
rect 24268 4768 24274 4820
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 26421 4811 26479 4817
rect 24360 4780 25820 4808
rect 24360 4768 24366 4780
rect 20088 4740 20116 4768
rect 18616 4712 20116 4740
rect 17497 4703 17555 4709
rect 14277 4675 14335 4681
rect 14277 4641 14289 4675
rect 14323 4672 14335 4675
rect 15838 4672 15844 4684
rect 14323 4644 15844 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 17512 4672 17540 4703
rect 19889 4675 19947 4681
rect 17512 4644 17816 4672
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 10560 4576 11529 4604
rect 10560 4564 10566 4576
rect 11517 4573 11529 4576
rect 11563 4604 11575 4607
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11563 4576 11621 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 13449 4607 13507 4613
rect 13449 4573 13461 4607
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 11146 4536 11152 4548
rect 7800 4508 11152 4536
rect 7800 4496 7806 4508
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11272 4539 11330 4545
rect 11272 4505 11284 4539
rect 11318 4536 11330 4539
rect 11422 4536 11428 4548
rect 11318 4508 11428 4536
rect 11318 4505 11330 4508
rect 11272 4499 11330 4505
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 13078 4496 13084 4548
rect 13136 4536 13142 4548
rect 13464 4536 13492 4567
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13964 4576 14473 4604
rect 13964 4564 13970 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16206 4604 16212 4616
rect 16163 4576 16212 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16206 4564 16212 4576
rect 16264 4604 16270 4616
rect 17681 4607 17739 4613
rect 17681 4604 17693 4607
rect 16264 4576 17693 4604
rect 16264 4564 16270 4576
rect 17681 4573 17693 4576
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 15197 4539 15255 4545
rect 15197 4536 15209 4539
rect 13136 4508 13492 4536
rect 13556 4508 15209 4536
rect 13136 4496 13142 4508
rect 7926 4468 7932 4480
rect 7668 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8018 4428 8024 4480
rect 8076 4428 8082 4480
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 9122 4468 9128 4480
rect 8527 4440 9128 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 11054 4468 11060 4480
rect 10183 4440 11060 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 11054 4428 11060 4440
rect 11112 4468 11118 4480
rect 11514 4468 11520 4480
rect 11112 4440 11520 4468
rect 11112 4428 11118 4440
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 12986 4468 12992 4480
rect 11756 4440 12992 4468
rect 11756 4428 11762 4440
rect 12986 4428 12992 4440
rect 13044 4468 13050 4480
rect 13556 4468 13584 4508
rect 15197 4505 15209 4508
rect 15243 4536 15255 4539
rect 15286 4536 15292 4548
rect 15243 4508 15292 4536
rect 15243 4505 15255 4508
rect 15197 4499 15255 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15473 4539 15531 4545
rect 15473 4505 15485 4539
rect 15519 4536 15531 4539
rect 15746 4536 15752 4548
rect 15519 4508 15752 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 16384 4539 16442 4545
rect 16384 4505 16396 4539
rect 16430 4536 16442 4539
rect 16666 4536 16672 4548
rect 16430 4508 16672 4536
rect 16430 4505 16442 4508
rect 16384 4499 16442 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 17788 4536 17816 4644
rect 19889 4641 19901 4675
rect 19935 4672 19947 4675
rect 20088 4672 20116 4712
rect 19935 4644 20116 4672
rect 19935 4641 19947 4644
rect 19889 4635 19947 4641
rect 21358 4632 21364 4684
rect 21416 4672 21422 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21416 4644 22017 4672
rect 21416 4632 21422 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 24026 4632 24032 4684
rect 24084 4632 24090 4684
rect 17948 4607 18006 4613
rect 17948 4573 17960 4607
rect 17994 4604 18006 4607
rect 18506 4604 18512 4616
rect 17994 4576 18512 4604
rect 17994 4573 18006 4576
rect 17948 4567 18006 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 19444 4576 20729 4604
rect 18046 4536 18052 4548
rect 17788 4508 18052 4536
rect 18046 4496 18052 4508
rect 18104 4536 18110 4548
rect 19242 4536 19248 4548
rect 18104 4508 19248 4536
rect 18104 4496 18110 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 19444 4480 19472 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20717 4567 20775 4573
rect 20806 4564 20812 4616
rect 20864 4564 20870 4616
rect 21910 4564 21916 4616
rect 21968 4604 21974 4616
rect 22261 4607 22319 4613
rect 22261 4604 22273 4607
rect 21968 4576 22273 4604
rect 21968 4564 21974 4576
rect 22261 4573 22273 4576
rect 22307 4573 22319 4607
rect 22261 4567 22319 4573
rect 23845 4607 23903 4613
rect 23845 4573 23857 4607
rect 23891 4604 23903 4607
rect 24228 4604 24256 4768
rect 25593 4743 25651 4749
rect 25593 4709 25605 4743
rect 25639 4740 25651 4743
rect 25682 4740 25688 4752
rect 25639 4712 25688 4740
rect 25639 4709 25651 4712
rect 25593 4703 25651 4709
rect 25682 4700 25688 4712
rect 25740 4700 25746 4752
rect 25792 4740 25820 4780
rect 26421 4777 26433 4811
rect 26467 4808 26479 4811
rect 26510 4808 26516 4820
rect 26467 4780 26516 4808
rect 26467 4777 26479 4780
rect 26421 4771 26479 4777
rect 26510 4768 26516 4780
rect 26568 4768 26574 4820
rect 27614 4768 27620 4820
rect 27672 4768 27678 4820
rect 27706 4768 27712 4820
rect 27764 4808 27770 4820
rect 35069 4811 35127 4817
rect 35069 4808 35081 4811
rect 27764 4780 35081 4808
rect 27764 4768 27770 4780
rect 35069 4777 35081 4780
rect 35115 4777 35127 4811
rect 35069 4771 35127 4777
rect 35529 4811 35587 4817
rect 35529 4777 35541 4811
rect 35575 4808 35587 4811
rect 37645 4811 37703 4817
rect 35575 4780 37412 4808
rect 35575 4777 35587 4780
rect 35529 4771 35587 4777
rect 28810 4740 28816 4752
rect 25792 4712 28816 4740
rect 28810 4700 28816 4712
rect 28868 4740 28874 4752
rect 28868 4712 29316 4740
rect 28868 4700 28874 4712
rect 24670 4672 24676 4684
rect 24320 4644 24676 4672
rect 24320 4616 24348 4644
rect 24670 4632 24676 4644
rect 24728 4672 24734 4684
rect 25179 4675 25237 4681
rect 25179 4672 25191 4675
rect 24728 4644 25191 4672
rect 24728 4632 24734 4644
rect 25179 4641 25191 4644
rect 25225 4641 25237 4675
rect 25179 4635 25237 4641
rect 25314 4632 25320 4684
rect 25372 4632 25378 4684
rect 26237 4675 26295 4681
rect 26237 4641 26249 4675
rect 26283 4672 26295 4675
rect 26970 4672 26976 4684
rect 26283 4644 26976 4672
rect 26283 4641 26295 4644
rect 26237 4635 26295 4641
rect 26970 4632 26976 4644
rect 27028 4632 27034 4684
rect 23891 4576 24256 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 24302 4564 24308 4616
rect 24360 4564 24366 4616
rect 25038 4564 25044 4616
rect 25096 4564 25102 4616
rect 26050 4564 26056 4616
rect 26108 4564 26114 4616
rect 26602 4564 26608 4616
rect 26660 4564 26666 4616
rect 26697 4607 26755 4613
rect 26697 4573 26709 4607
rect 26743 4573 26755 4607
rect 26697 4567 26755 4573
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27985 4607 28043 4613
rect 27985 4604 27997 4607
rect 27295 4576 27997 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 27985 4573 27997 4576
rect 28031 4604 28043 4607
rect 28258 4604 28264 4616
rect 28031 4576 28264 4604
rect 28031 4573 28043 4576
rect 27985 4567 28043 4573
rect 19610 4496 19616 4548
rect 19668 4536 19674 4548
rect 20254 4536 20260 4548
rect 19668 4508 20260 4536
rect 19668 4496 19674 4508
rect 20254 4496 20260 4508
rect 20312 4496 20318 4548
rect 26326 4496 26332 4548
rect 26384 4536 26390 4548
rect 26712 4536 26740 4567
rect 28258 4564 28264 4576
rect 28316 4564 28322 4616
rect 28350 4564 28356 4616
rect 28408 4564 28414 4616
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 28460 4576 28825 4604
rect 26384 4508 26740 4536
rect 26384 4496 26390 4508
rect 28074 4496 28080 4548
rect 28132 4536 28138 4548
rect 28460 4536 28488 4576
rect 28813 4573 28825 4576
rect 28859 4573 28871 4607
rect 29288 4604 29316 4712
rect 30742 4700 30748 4752
rect 30800 4740 30806 4752
rect 31021 4743 31079 4749
rect 31021 4740 31033 4743
rect 30800 4712 31033 4740
rect 30800 4700 30806 4712
rect 31021 4709 31033 4712
rect 31067 4740 31079 4743
rect 31478 4740 31484 4752
rect 31067 4712 31484 4740
rect 31067 4709 31079 4712
rect 31021 4703 31079 4709
rect 31478 4700 31484 4712
rect 31536 4700 31542 4752
rect 32582 4700 32588 4752
rect 32640 4740 32646 4752
rect 36170 4740 36176 4752
rect 32640 4712 36176 4740
rect 32640 4700 32646 4712
rect 36170 4700 36176 4712
rect 36228 4700 36234 4752
rect 36446 4700 36452 4752
rect 36504 4700 36510 4752
rect 37384 4740 37412 4780
rect 37645 4777 37657 4811
rect 37691 4808 37703 4811
rect 37734 4808 37740 4820
rect 37691 4780 37740 4808
rect 37691 4777 37703 4780
rect 37645 4771 37703 4777
rect 37734 4768 37740 4780
rect 37792 4768 37798 4820
rect 37918 4768 37924 4820
rect 37976 4768 37982 4820
rect 38010 4768 38016 4820
rect 38068 4768 38074 4820
rect 38838 4768 38844 4820
rect 38896 4768 38902 4820
rect 39577 4811 39635 4817
rect 39577 4777 39589 4811
rect 39623 4808 39635 4811
rect 39666 4808 39672 4820
rect 39623 4780 39672 4808
rect 39623 4777 39635 4780
rect 39577 4771 39635 4777
rect 39666 4768 39672 4780
rect 39724 4768 39730 4820
rect 41874 4808 41880 4820
rect 40420 4780 41880 4808
rect 37936 4740 37964 4768
rect 40420 4740 40448 4780
rect 41874 4768 41880 4780
rect 41932 4768 41938 4820
rect 42429 4811 42487 4817
rect 42429 4777 42441 4811
rect 42475 4808 42487 4811
rect 42702 4808 42708 4820
rect 42475 4780 42708 4808
rect 42475 4777 42487 4780
rect 42429 4771 42487 4777
rect 42702 4768 42708 4780
rect 42760 4768 42766 4820
rect 46014 4768 46020 4820
rect 46072 4768 46078 4820
rect 46474 4768 46480 4820
rect 46532 4768 46538 4820
rect 48498 4768 48504 4820
rect 48556 4808 48562 4820
rect 48777 4811 48835 4817
rect 48777 4808 48789 4811
rect 48556 4780 48789 4808
rect 48556 4768 48562 4780
rect 48777 4777 48789 4780
rect 48823 4808 48835 4811
rect 50154 4808 50160 4820
rect 48823 4780 50160 4808
rect 48823 4777 48835 4780
rect 48777 4771 48835 4777
rect 50154 4768 50160 4780
rect 50212 4768 50218 4820
rect 51350 4768 51356 4820
rect 51408 4808 51414 4820
rect 51721 4811 51779 4817
rect 51721 4808 51733 4811
rect 51408 4780 51733 4808
rect 51408 4768 51414 4780
rect 51721 4777 51733 4780
rect 51767 4777 51779 4811
rect 51721 4771 51779 4777
rect 52546 4768 52552 4820
rect 52604 4768 52610 4820
rect 55125 4811 55183 4817
rect 55125 4777 55137 4811
rect 55171 4808 55183 4811
rect 57146 4808 57152 4820
rect 55171 4780 57152 4808
rect 55171 4777 55183 4780
rect 55125 4771 55183 4777
rect 57146 4768 57152 4780
rect 57204 4768 57210 4820
rect 57698 4768 57704 4820
rect 57756 4808 57762 4820
rect 57756 4780 57928 4808
rect 57756 4768 57762 4780
rect 41046 4740 41052 4752
rect 37384 4712 37964 4740
rect 39408 4712 40448 4740
rect 40604 4712 41052 4740
rect 29365 4675 29423 4681
rect 29365 4641 29377 4675
rect 29411 4672 29423 4675
rect 31294 4672 31300 4684
rect 29411 4644 31300 4672
rect 29411 4641 29423 4644
rect 29365 4635 29423 4641
rect 31294 4632 31300 4644
rect 31352 4632 31358 4684
rect 33321 4675 33379 4681
rect 33321 4672 33333 4675
rect 32416 4644 33333 4672
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29288 4576 29561 4604
rect 28813 4567 28871 4573
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 28132 4508 28488 4536
rect 28537 4539 28595 4545
rect 28132 4496 28138 4508
rect 28537 4505 28549 4539
rect 28583 4536 28595 4539
rect 29178 4536 29184 4548
rect 28583 4508 29184 4536
rect 28583 4505 28595 4508
rect 28537 4499 28595 4505
rect 29178 4496 29184 4508
rect 29236 4496 29242 4548
rect 30190 4496 30196 4548
rect 30248 4536 30254 4548
rect 30377 4539 30435 4545
rect 30377 4536 30389 4539
rect 30248 4508 30389 4536
rect 30248 4496 30254 4508
rect 30377 4505 30389 4508
rect 30423 4505 30435 4539
rect 32030 4536 32036 4548
rect 30377 4499 30435 4505
rect 30484 4508 32036 4536
rect 13044 4440 13584 4468
rect 13633 4471 13691 4477
rect 13044 4428 13050 4440
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 14090 4468 14096 4480
rect 13679 4440 14096 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14366 4428 14372 4480
rect 14424 4428 14430 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15381 4471 15439 4477
rect 15381 4468 15393 4471
rect 14608 4440 15393 4468
rect 14608 4428 14614 4440
rect 15381 4437 15393 4440
rect 15427 4437 15439 4471
rect 15381 4431 15439 4437
rect 16114 4428 16120 4480
rect 16172 4468 16178 4480
rect 18874 4468 18880 4480
rect 16172 4440 18880 4468
rect 16172 4428 16178 4440
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19061 4471 19119 4477
rect 19061 4437 19073 4471
rect 19107 4468 19119 4471
rect 19426 4468 19432 4480
rect 19107 4440 19432 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 20073 4471 20131 4477
rect 20073 4468 20085 4471
rect 19751 4440 20085 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 20073 4437 20085 4440
rect 20119 4437 20131 4471
rect 20073 4431 20131 4437
rect 21082 4428 21088 4480
rect 21140 4468 21146 4480
rect 21453 4471 21511 4477
rect 21453 4468 21465 4471
rect 21140 4440 21465 4468
rect 21140 4428 21146 4440
rect 21453 4437 21465 4440
rect 21499 4437 21511 4471
rect 21453 4431 21511 4437
rect 23474 4428 23480 4480
rect 23532 4428 23538 4480
rect 23934 4428 23940 4480
rect 23992 4428 23998 4480
rect 24394 4428 24400 4480
rect 24452 4428 24458 4480
rect 26878 4428 26884 4480
rect 26936 4428 26942 4480
rect 28626 4428 28632 4480
rect 28684 4428 28690 4480
rect 28718 4428 28724 4480
rect 28776 4468 28782 4480
rect 30484 4468 30512 4508
rect 32030 4496 32036 4508
rect 32088 4496 32094 4548
rect 32248 4539 32306 4545
rect 32248 4505 32260 4539
rect 32294 4536 32306 4539
rect 32416 4536 32444 4644
rect 33321 4641 33333 4644
rect 33367 4641 33379 4675
rect 33321 4635 33379 4641
rect 33778 4632 33784 4684
rect 33836 4672 33842 4684
rect 34425 4675 34483 4681
rect 34425 4672 34437 4675
rect 33836 4644 34437 4672
rect 33836 4632 33842 4644
rect 34425 4641 34437 4644
rect 34471 4672 34483 4675
rect 34471 4644 35572 4672
rect 34471 4641 34483 4644
rect 34425 4635 34483 4641
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4604 32551 4607
rect 32539 4576 32628 4604
rect 32539 4573 32551 4576
rect 32493 4567 32551 4573
rect 32294 4508 32444 4536
rect 32600 4536 32628 4576
rect 32858 4564 32864 4616
rect 32916 4604 32922 4616
rect 33137 4607 33195 4613
rect 33137 4604 33149 4607
rect 32916 4576 33149 4604
rect 32916 4564 32922 4576
rect 33137 4573 33149 4576
rect 33183 4573 33195 4607
rect 33137 4567 33195 4573
rect 33502 4564 33508 4616
rect 33560 4564 33566 4616
rect 33870 4564 33876 4616
rect 33928 4564 33934 4616
rect 35345 4607 35403 4613
rect 35345 4573 35357 4607
rect 35391 4573 35403 4607
rect 35544 4604 35572 4644
rect 35618 4632 35624 4684
rect 35676 4672 35682 4684
rect 35805 4675 35863 4681
rect 35805 4672 35817 4675
rect 35676 4644 35817 4672
rect 35676 4632 35682 4644
rect 35805 4641 35817 4644
rect 35851 4641 35863 4675
rect 35805 4635 35863 4641
rect 36538 4632 36544 4684
rect 36596 4672 36602 4684
rect 36725 4675 36783 4681
rect 36725 4672 36737 4675
rect 36596 4644 36737 4672
rect 36596 4632 36602 4644
rect 36725 4641 36737 4644
rect 36771 4641 36783 4675
rect 36725 4635 36783 4641
rect 36998 4632 37004 4684
rect 37056 4632 37062 4684
rect 35710 4604 35716 4616
rect 35544 4576 35716 4604
rect 35345 4567 35403 4573
rect 32766 4536 32772 4548
rect 32600 4508 32772 4536
rect 32294 4505 32306 4508
rect 32248 4499 32306 4505
rect 32766 4496 32772 4508
rect 32824 4536 32830 4548
rect 33520 4536 33548 4564
rect 32824 4508 33548 4536
rect 32824 4496 32830 4508
rect 34146 4496 34152 4548
rect 34204 4536 34210 4548
rect 34204 4508 34376 4536
rect 34204 4496 34210 4508
rect 28776 4440 30512 4468
rect 31113 4471 31171 4477
rect 28776 4428 28782 4440
rect 31113 4437 31125 4471
rect 31159 4468 31171 4471
rect 31938 4468 31944 4480
rect 31159 4440 31944 4468
rect 31159 4437 31171 4440
rect 31113 4431 31171 4437
rect 31938 4428 31944 4440
rect 31996 4428 32002 4480
rect 32582 4428 32588 4480
rect 32640 4428 32646 4480
rect 34348 4468 34376 4508
rect 35158 4496 35164 4548
rect 35216 4496 35222 4548
rect 35360 4536 35388 4567
rect 35710 4564 35716 4576
rect 35768 4564 35774 4616
rect 35989 4607 36047 4613
rect 35989 4573 36001 4607
rect 36035 4604 36047 4607
rect 36170 4604 36176 4616
rect 36035 4576 36176 4604
rect 36035 4573 36047 4576
rect 35989 4567 36047 4573
rect 36170 4564 36176 4576
rect 36228 4564 36234 4616
rect 36814 4564 36820 4616
rect 36872 4613 36878 4616
rect 39408 4613 39436 4712
rect 40218 4632 40224 4684
rect 40276 4672 40282 4684
rect 40604 4681 40632 4712
rect 41046 4700 41052 4712
rect 41104 4700 41110 4752
rect 41230 4700 41236 4752
rect 41288 4700 41294 4752
rect 40589 4675 40647 4681
rect 40589 4672 40601 4675
rect 40276 4644 40601 4672
rect 40276 4632 40282 4644
rect 40589 4641 40601 4644
rect 40635 4641 40647 4675
rect 40589 4635 40647 4641
rect 41322 4632 41328 4684
rect 41380 4672 41386 4684
rect 41509 4675 41567 4681
rect 41509 4672 41521 4675
rect 41380 4644 41521 4672
rect 41380 4632 41386 4644
rect 41509 4641 41521 4644
rect 41555 4641 41567 4675
rect 41509 4635 41567 4641
rect 41647 4675 41705 4681
rect 41647 4641 41659 4675
rect 41693 4672 41705 4675
rect 41966 4672 41972 4684
rect 41693 4644 41972 4672
rect 41693 4641 41705 4644
rect 41647 4635 41705 4641
rect 41966 4632 41972 4644
rect 42024 4632 42030 4684
rect 43901 4675 43959 4681
rect 43901 4641 43913 4675
rect 43947 4672 43959 4675
rect 44174 4672 44180 4684
rect 43947 4644 44180 4672
rect 43947 4641 43959 4644
rect 43901 4635 43959 4641
rect 44174 4632 44180 4644
rect 44232 4632 44238 4684
rect 44818 4632 44824 4684
rect 44876 4672 44882 4684
rect 46492 4672 46520 4768
rect 47673 4743 47731 4749
rect 47673 4709 47685 4743
rect 47719 4740 47731 4743
rect 48682 4740 48688 4752
rect 47719 4712 48688 4740
rect 47719 4709 47731 4712
rect 47673 4703 47731 4709
rect 48682 4700 48688 4712
rect 48740 4700 48746 4752
rect 49145 4743 49203 4749
rect 49145 4709 49157 4743
rect 49191 4740 49203 4743
rect 49418 4740 49424 4752
rect 49191 4712 49424 4740
rect 49191 4709 49203 4712
rect 49145 4703 49203 4709
rect 49418 4700 49424 4712
rect 49476 4700 49482 4752
rect 49513 4743 49571 4749
rect 49513 4709 49525 4743
rect 49559 4740 49571 4743
rect 50798 4740 50804 4752
rect 49559 4712 50804 4740
rect 49559 4709 49571 4712
rect 49513 4703 49571 4709
rect 46569 4675 46627 4681
rect 46569 4672 46581 4675
rect 44876 4644 46060 4672
rect 46492 4644 46581 4672
rect 44876 4632 44882 4644
rect 36872 4607 36900 4613
rect 36888 4573 36900 4607
rect 36872 4567 36900 4573
rect 39025 4607 39083 4613
rect 39025 4573 39037 4607
rect 39071 4573 39083 4607
rect 39025 4567 39083 4573
rect 39393 4607 39451 4613
rect 39393 4573 39405 4607
rect 39439 4573 39451 4607
rect 39393 4567 39451 4573
rect 36872 4564 36878 4567
rect 35894 4536 35900 4548
rect 35360 4508 35900 4536
rect 35894 4496 35900 4508
rect 35952 4496 35958 4548
rect 38657 4539 38715 4545
rect 38657 4536 38669 4539
rect 37476 4508 38669 4536
rect 37476 4468 37504 4508
rect 38657 4505 38669 4508
rect 38703 4505 38715 4539
rect 39040 4536 39068 4567
rect 40402 4564 40408 4616
rect 40460 4564 40466 4616
rect 40773 4607 40831 4613
rect 40773 4573 40785 4607
rect 40819 4573 40831 4607
rect 40773 4567 40831 4573
rect 40586 4536 40592 4548
rect 39040 4508 40592 4536
rect 38657 4499 38715 4505
rect 40586 4496 40592 4508
rect 40644 4496 40650 4548
rect 34348 4440 37504 4468
rect 38286 4428 38292 4480
rect 38344 4428 38350 4480
rect 39850 4428 39856 4480
rect 39908 4428 39914 4480
rect 40788 4468 40816 4567
rect 41782 4564 41788 4616
rect 41840 4564 41846 4616
rect 42610 4564 42616 4616
rect 42668 4604 42674 4616
rect 44082 4604 44088 4616
rect 42668 4576 44088 4604
rect 42668 4564 42674 4576
rect 44082 4564 44088 4576
rect 44140 4564 44146 4616
rect 44634 4564 44640 4616
rect 44692 4564 44698 4616
rect 44910 4564 44916 4616
rect 44968 4604 44974 4616
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 44968 4576 45201 4604
rect 44968 4564 44974 4576
rect 45189 4573 45201 4576
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 45922 4564 45928 4616
rect 45980 4564 45986 4616
rect 46032 4604 46060 4644
rect 46569 4641 46581 4644
rect 46615 4641 46627 4675
rect 48041 4675 48099 4681
rect 48041 4672 48053 4675
rect 46569 4635 46627 4641
rect 46676 4644 48053 4672
rect 46676 4604 46704 4644
rect 48041 4641 48053 4644
rect 48087 4672 48099 4675
rect 48409 4675 48467 4681
rect 48409 4672 48421 4675
rect 48087 4644 48421 4672
rect 48087 4641 48099 4644
rect 48041 4635 48099 4641
rect 48409 4641 48421 4644
rect 48455 4672 48467 4675
rect 49528 4672 49556 4703
rect 50798 4700 50804 4712
rect 50856 4740 50862 4752
rect 52564 4740 52592 4768
rect 50856 4712 52592 4740
rect 50856 4700 50862 4712
rect 55950 4700 55956 4752
rect 56008 4740 56014 4752
rect 56502 4740 56508 4752
rect 56008 4712 56508 4740
rect 56008 4700 56014 4712
rect 56502 4700 56508 4712
rect 56560 4700 56566 4752
rect 51166 4672 51172 4684
rect 48455 4644 49556 4672
rect 49620 4644 51172 4672
rect 48455 4641 48467 4644
rect 48409 4635 48467 4641
rect 46032 4576 46704 4604
rect 47302 4564 47308 4616
rect 47360 4564 47366 4616
rect 47486 4564 47492 4616
rect 47544 4564 47550 4616
rect 48961 4607 49019 4613
rect 48961 4573 48973 4607
rect 49007 4604 49019 4607
rect 49620 4604 49648 4644
rect 51166 4632 51172 4644
rect 51224 4632 51230 4684
rect 52454 4632 52460 4684
rect 52512 4672 52518 4684
rect 53285 4675 53343 4681
rect 53285 4672 53297 4675
rect 52512 4644 53297 4672
rect 52512 4632 52518 4644
rect 53285 4641 53297 4644
rect 53331 4641 53343 4675
rect 53285 4635 53343 4641
rect 54018 4632 54024 4684
rect 54076 4672 54082 4684
rect 57900 4681 57928 4780
rect 55309 4675 55367 4681
rect 55309 4672 55321 4675
rect 54076 4644 55321 4672
rect 54076 4632 54082 4644
rect 55309 4641 55321 4644
rect 55355 4672 55367 4675
rect 57885 4675 57943 4681
rect 55355 4644 55904 4672
rect 55355 4641 55367 4644
rect 55309 4635 55367 4641
rect 49007 4576 49648 4604
rect 49007 4573 49019 4576
rect 48961 4567 49019 4573
rect 49694 4564 49700 4616
rect 49752 4604 49758 4616
rect 50157 4607 50215 4613
rect 50157 4604 50169 4607
rect 49752 4576 50169 4604
rect 49752 4564 49758 4576
rect 50157 4573 50169 4576
rect 50203 4573 50215 4607
rect 50157 4567 50215 4573
rect 51442 4564 51448 4616
rect 51500 4564 51506 4616
rect 51905 4607 51963 4613
rect 51905 4573 51917 4607
rect 51951 4604 51963 4607
rect 51994 4604 52000 4616
rect 51951 4576 52000 4604
rect 51951 4573 51963 4576
rect 51905 4567 51963 4573
rect 51994 4564 52000 4576
rect 52052 4564 52058 4616
rect 52086 4564 52092 4616
rect 52144 4564 52150 4616
rect 53098 4564 53104 4616
rect 53156 4564 53162 4616
rect 54110 4564 54116 4616
rect 54168 4564 54174 4616
rect 54573 4607 54631 4613
rect 54573 4573 54585 4607
rect 54619 4573 54631 4607
rect 54573 4567 54631 4573
rect 43656 4539 43714 4545
rect 43656 4505 43668 4539
rect 43702 4536 43714 4539
rect 43993 4539 44051 4545
rect 43993 4536 44005 4539
rect 43702 4508 44005 4536
rect 43702 4505 43714 4508
rect 43656 4499 43714 4505
rect 43993 4505 44005 4508
rect 44039 4505 44051 4539
rect 43993 4499 44051 4505
rect 49881 4539 49939 4545
rect 49881 4505 49893 4539
rect 49927 4536 49939 4539
rect 51350 4536 51356 4548
rect 49927 4508 51356 4536
rect 49927 4505 49939 4508
rect 49881 4499 49939 4505
rect 51350 4496 51356 4508
rect 51408 4496 51414 4548
rect 54588 4536 54616 4567
rect 55490 4564 55496 4616
rect 55548 4564 55554 4616
rect 55674 4564 55680 4616
rect 55732 4564 55738 4616
rect 55766 4564 55772 4616
rect 55824 4564 55830 4616
rect 55876 4604 55904 4644
rect 57885 4641 57897 4675
rect 57931 4641 57943 4675
rect 57885 4635 57943 4641
rect 57629 4607 57687 4613
rect 55876 4576 57468 4604
rect 57440 4548 57468 4576
rect 57629 4573 57641 4607
rect 57675 4604 57687 4607
rect 57790 4604 57796 4616
rect 57675 4576 57796 4604
rect 57675 4573 57687 4576
rect 57629 4567 57687 4573
rect 57790 4564 57796 4576
rect 57848 4564 57854 4616
rect 58158 4564 58164 4616
rect 58216 4564 58222 4616
rect 58253 4607 58311 4613
rect 58253 4573 58265 4607
rect 58299 4573 58311 4607
rect 58253 4567 58311 4573
rect 56594 4536 56600 4548
rect 52656 4508 54524 4536
rect 54588 4508 56600 4536
rect 42521 4471 42579 4477
rect 42521 4468 42533 4471
rect 40788 4440 42533 4468
rect 42521 4437 42533 4440
rect 42567 4468 42579 4471
rect 43806 4468 43812 4480
rect 42567 4440 43812 4468
rect 42567 4437 42579 4440
rect 42521 4431 42579 4437
rect 43806 4428 43812 4440
rect 43864 4428 43870 4480
rect 45002 4428 45008 4480
rect 45060 4428 45066 4480
rect 45278 4428 45284 4480
rect 45336 4428 45342 4480
rect 46750 4428 46756 4480
rect 46808 4428 46814 4480
rect 49602 4428 49608 4480
rect 49660 4468 49666 4480
rect 49789 4471 49847 4477
rect 49789 4468 49801 4471
rect 49660 4440 49801 4468
rect 49660 4428 49666 4440
rect 49789 4437 49801 4440
rect 49835 4468 49847 4471
rect 50522 4468 50528 4480
rect 49835 4440 50528 4468
rect 49835 4437 49847 4440
rect 49789 4431 49847 4437
rect 50522 4428 50528 4440
rect 50580 4428 50586 4480
rect 50798 4428 50804 4480
rect 50856 4428 50862 4480
rect 50890 4428 50896 4480
rect 50948 4428 50954 4480
rect 52656 4477 52684 4508
rect 52641 4471 52699 4477
rect 52641 4437 52653 4471
rect 52687 4437 52699 4471
rect 52641 4431 52699 4437
rect 52730 4428 52736 4480
rect 52788 4428 52794 4480
rect 53190 4428 53196 4480
rect 53248 4428 53254 4480
rect 53558 4428 53564 4480
rect 53616 4428 53622 4480
rect 54496 4468 54524 4508
rect 56594 4496 56600 4508
rect 56652 4496 56658 4548
rect 57422 4496 57428 4548
rect 57480 4536 57486 4548
rect 58268 4536 58296 4567
rect 57480 4508 58296 4536
rect 57480 4496 57486 4508
rect 56042 4468 56048 4480
rect 54496 4440 56048 4468
rect 56042 4428 56048 4440
rect 56100 4428 56106 4480
rect 56410 4428 56416 4480
rect 56468 4428 56474 4480
rect 57054 4428 57060 4480
rect 57112 4468 57118 4480
rect 57977 4471 58035 4477
rect 57977 4468 57989 4471
rect 57112 4440 57989 4468
rect 57112 4428 57118 4440
rect 57977 4437 57989 4440
rect 58023 4437 58035 4471
rect 57977 4431 58035 4437
rect 1104 4378 59040 4400
rect 1104 4326 15394 4378
rect 15446 4326 15458 4378
rect 15510 4326 15522 4378
rect 15574 4326 15586 4378
rect 15638 4326 15650 4378
rect 15702 4326 29838 4378
rect 29890 4326 29902 4378
rect 29954 4326 29966 4378
rect 30018 4326 30030 4378
rect 30082 4326 30094 4378
rect 30146 4326 44282 4378
rect 44334 4326 44346 4378
rect 44398 4326 44410 4378
rect 44462 4326 44474 4378
rect 44526 4326 44538 4378
rect 44590 4326 58726 4378
rect 58778 4326 58790 4378
rect 58842 4326 58854 4378
rect 58906 4326 58918 4378
rect 58970 4326 58982 4378
rect 59034 4326 59040 4378
rect 1104 4304 59040 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 2924 4236 3249 4264
rect 2924 4224 2930 4236
rect 3237 4233 3249 4236
rect 3283 4233 3295 4267
rect 3237 4227 3295 4233
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 3697 4267 3755 4273
rect 3697 4264 3709 4267
rect 3660 4236 3709 4264
rect 3660 4224 3666 4236
rect 3697 4233 3709 4236
rect 3743 4233 3755 4267
rect 3697 4227 3755 4233
rect 4341 4267 4399 4273
rect 4341 4233 4353 4267
rect 4387 4264 4399 4267
rect 4614 4264 4620 4276
rect 4387 4236 4620 4264
rect 4387 4233 4399 4236
rect 4341 4227 4399 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 4801 4267 4859 4273
rect 4801 4233 4813 4267
rect 4847 4264 4859 4267
rect 5074 4264 5080 4276
rect 4847 4236 5080 4264
rect 4847 4233 4859 4236
rect 4801 4227 4859 4233
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4233 7527 4267
rect 7469 4227 7527 4233
rect 2032 4199 2090 4205
rect 2032 4165 2044 4199
rect 2078 4196 2090 4199
rect 2222 4196 2228 4208
rect 2078 4168 2228 4196
rect 2078 4165 2090 4168
rect 2032 4159 2090 4165
rect 2222 4156 2228 4168
rect 2280 4156 2286 4208
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 4709 4199 4767 4205
rect 4709 4196 4721 4199
rect 3568 4168 4721 4196
rect 3568 4156 3574 4168
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 3620 4137 3648 4168
rect 4709 4165 4721 4168
rect 4755 4196 4767 4199
rect 5626 4196 5632 4208
rect 4755 4168 5632 4196
rect 4755 4165 4767 4168
rect 4709 4159 4767 4165
rect 5626 4156 5632 4168
rect 5684 4156 5690 4208
rect 7098 4196 7104 4208
rect 6012 4168 7104 4196
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4246 4128 4252 4140
rect 4111 4100 4252 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 6012 4128 6040 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 4908 4100 6040 4128
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3786 4060 3792 4072
rect 3016 4032 3792 4060
rect 3016 4020 3022 4032
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4908 4060 4936 4100
rect 6086 4088 6092 4140
rect 6144 4088 6150 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6822 4128 6828 4140
rect 6595 4100 6828 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7484 4128 7512 4227
rect 7558 4224 7564 4276
rect 7616 4224 7622 4276
rect 7926 4224 7932 4276
rect 7984 4224 7990 4276
rect 9398 4224 9404 4276
rect 9456 4224 9462 4276
rect 9858 4224 9864 4276
rect 9916 4224 9922 4276
rect 10134 4224 10140 4276
rect 10192 4224 10198 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 11480 4236 11529 4264
rect 11480 4224 11486 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11517 4227 11575 4233
rect 11698 4224 11704 4276
rect 11756 4224 11762 4276
rect 14093 4267 14151 4273
rect 14093 4233 14105 4267
rect 14139 4264 14151 4267
rect 14366 4264 14372 4276
rect 14139 4236 14372 4264
rect 14139 4233 14151 4236
rect 14093 4227 14151 4233
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 16390 4264 16396 4276
rect 15896 4236 16396 4264
rect 15896 4224 15902 4236
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16945 4267 17003 4273
rect 16945 4233 16957 4267
rect 16991 4264 17003 4267
rect 17218 4264 17224 4276
rect 16991 4236 17224 4264
rect 16991 4233 17003 4236
rect 16945 4227 17003 4233
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 17313 4267 17371 4273
rect 17313 4233 17325 4267
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 17405 4267 17463 4273
rect 17405 4233 17417 4267
rect 17451 4264 17463 4267
rect 17494 4264 17500 4276
rect 17451 4236 17500 4264
rect 17451 4233 17463 4236
rect 17405 4227 17463 4233
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 8021 4199 8079 4205
rect 8021 4196 8033 4199
rect 7708 4168 8033 4196
rect 7708 4156 7714 4168
rect 8021 4165 8033 4168
rect 8067 4165 8079 4199
rect 8021 4159 8079 4165
rect 8757 4199 8815 4205
rect 8757 4165 8769 4199
rect 8803 4196 8815 4199
rect 9030 4196 9036 4208
rect 8803 4168 9036 4196
rect 8803 4165 8815 4168
rect 8757 4159 8815 4165
rect 9030 4156 9036 4168
rect 9088 4196 9094 4208
rect 9416 4196 9444 4224
rect 9088 4168 9444 4196
rect 9088 4156 9094 4168
rect 10594 4156 10600 4208
rect 10652 4196 10658 4208
rect 11716 4196 11744 4224
rect 10652 4168 11744 4196
rect 10652 4156 10658 4168
rect 13998 4156 14004 4208
rect 14056 4156 14062 4208
rect 15286 4156 15292 4208
rect 15344 4156 15350 4208
rect 17328 4196 17356 4227
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 19610 4264 19616 4276
rect 18524 4236 19616 4264
rect 18524 4196 18552 4236
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 20625 4267 20683 4273
rect 20625 4233 20637 4267
rect 20671 4264 20683 4267
rect 20898 4264 20904 4276
rect 20671 4236 20904 4264
rect 20671 4233 20683 4236
rect 20625 4227 20683 4233
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 23385 4267 23443 4273
rect 23385 4233 23397 4267
rect 23431 4264 23443 4267
rect 24302 4264 24308 4276
rect 23431 4236 24308 4264
rect 23431 4233 23443 4236
rect 23385 4227 23443 4233
rect 24302 4224 24308 4236
rect 24360 4224 24366 4276
rect 24394 4224 24400 4276
rect 24452 4264 24458 4276
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24452 4236 24777 4264
rect 24452 4224 24458 4236
rect 24765 4233 24777 4236
rect 24811 4233 24823 4267
rect 24765 4227 24823 4233
rect 27614 4224 27620 4276
rect 27672 4224 27678 4276
rect 29825 4267 29883 4273
rect 29825 4233 29837 4267
rect 29871 4233 29883 4267
rect 29825 4227 29883 4233
rect 32401 4267 32459 4273
rect 32401 4233 32413 4267
rect 32447 4264 32459 4267
rect 32582 4264 32588 4276
rect 32447 4236 32588 4264
rect 32447 4233 32459 4236
rect 32401 4227 32459 4233
rect 17328 4168 18552 4196
rect 20530 4156 20536 4208
rect 20588 4156 20594 4208
rect 22204 4168 22416 4196
rect 7064 4100 7512 4128
rect 7064 4088 7070 4100
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7742 4128 7748 4140
rect 7616 4100 7748 4128
rect 7616 4088 7622 4100
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8570 4128 8576 4140
rect 8435 4100 8576 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9364 4100 9413 4128
rect 9364 4088 9370 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9677 4131 9735 4137
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 9858 4128 9864 4140
rect 9723 4100 9864 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 9968 4100 10885 4128
rect 4212 4032 4936 4060
rect 4212 4020 4218 4032
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5810 4060 5816 4072
rect 5040 4032 5816 4060
rect 5040 4020 5046 4032
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6236 4032 6745 4060
rect 6236 4020 6242 4032
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 7098 4020 7104 4072
rect 7156 4020 7162 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7248 4032 7389 4060
rect 7248 4020 7254 4032
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 9968 4060 9996 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13446 4088 13452 4140
rect 13504 4088 13510 4140
rect 14016 4128 14044 4156
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14016 4100 15117 4128
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15304 4128 15332 4156
rect 15304 4100 17540 4128
rect 15105 4091 15163 4097
rect 7423 4032 9996 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 12158 4020 12164 4072
rect 12216 4020 12222 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12802 4060 12808 4072
rect 12483 4032 12808 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12894 4020 12900 4072
rect 12952 4020 12958 4072
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 13004 4032 13185 4060
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 5074 3992 5080 4004
rect 3200 3964 5080 3992
rect 3200 3952 3206 3964
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 8205 3995 8263 4001
rect 5684 3964 6500 3992
rect 5684 3952 5690 3964
rect 1670 3884 1676 3936
rect 1728 3884 1734 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 6362 3924 6368 3936
rect 4295 3896 6368 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6472 3933 6500 3964
rect 7024 3964 8156 3992
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 7024 3924 7052 3964
rect 6503 3896 7052 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 7616 3896 8033 3924
rect 7616 3884 7622 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8128 3924 8156 3964
rect 8205 3961 8217 3995
rect 8251 3992 8263 3995
rect 10594 3992 10600 4004
rect 8251 3964 10600 3992
rect 8251 3961 8263 3964
rect 8205 3955 8263 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 9122 3924 9128 3936
rect 8128 3896 9128 3924
rect 8021 3887 8079 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 13004 3924 13032 4032
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 13311 4063 13369 4069
rect 13311 4029 13323 4063
rect 13357 4060 13369 4063
rect 13630 4060 13636 4072
rect 13357 4032 13636 4060
rect 13357 4029 13369 4032
rect 13311 4023 13369 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 13832 4032 14749 4060
rect 11572 3896 13032 3924
rect 11572 3884 11578 3896
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 13832 3924 13860 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4060 15347 4063
rect 15378 4060 15384 4072
rect 15335 4032 15384 4060
rect 15335 4029 15347 4032
rect 15289 4023 15347 4029
rect 15378 4020 15384 4032
rect 15436 4060 15442 4072
rect 15930 4060 15936 4072
rect 15436 4032 15936 4060
rect 15436 4020 15442 4032
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 17512 4069 17540 4100
rect 17954 4088 17960 4140
rect 18012 4088 18018 4140
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4128 20039 4131
rect 20806 4128 20812 4140
rect 20027 4100 20812 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 21634 4088 21640 4140
rect 21692 4088 21698 4140
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22204 4128 22232 4168
rect 22278 4137 22284 4140
rect 22112 4100 22232 4128
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 19058 4020 19064 4072
rect 19116 4069 19122 4072
rect 19116 4063 19165 4069
rect 19116 4029 19119 4063
rect 19153 4029 19165 4063
rect 19116 4023 19165 4029
rect 19116 4020 19122 4023
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 19484 4032 20177 4060
rect 19484 4020 19490 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 20165 4023 20223 4029
rect 20364 4032 20453 4060
rect 20364 4004 20392 4032
rect 20441 4029 20453 4032
rect 20487 4060 20499 4063
rect 21269 4063 21327 4069
rect 21269 4060 21281 4063
rect 20487 4032 21281 4060
rect 20487 4029 20499 4032
rect 20441 4023 20499 4029
rect 21269 4029 21281 4032
rect 21315 4060 21327 4063
rect 22112 4060 22140 4100
rect 22272 4091 22284 4137
rect 22278 4088 22284 4091
rect 22336 4088 22342 4140
rect 22388 4128 22416 4168
rect 23934 4156 23940 4208
rect 23992 4196 23998 4208
rect 23992 4168 25084 4196
rect 23992 4156 23998 4168
rect 22388 4100 24992 4128
rect 21315 4032 22140 4060
rect 23753 4063 23811 4069
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 23753 4029 23765 4063
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 13964 3964 15669 3992
rect 13964 3952 13970 3964
rect 15657 3961 15669 3964
rect 15703 3961 15715 3995
rect 16850 3992 16856 4004
rect 15657 3955 15715 3961
rect 16546 3964 16856 3992
rect 13688 3896 13860 3924
rect 13688 3884 13694 3896
rect 14182 3884 14188 3936
rect 14240 3884 14246 3936
rect 14918 3884 14924 3936
rect 14976 3884 14982 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15068 3896 16037 3924
rect 15068 3884 15074 3896
rect 16025 3893 16037 3896
rect 16071 3924 16083 3927
rect 16546 3924 16574 3964
rect 16850 3952 16856 3964
rect 16908 3992 16914 4004
rect 17862 3992 17868 4004
rect 16908 3964 17868 3992
rect 16908 3952 16914 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 19521 3995 19579 4001
rect 19521 3961 19533 3995
rect 19567 3992 19579 3995
rect 19886 3992 19892 4004
rect 19567 3964 19892 3992
rect 19567 3961 19579 3964
rect 19521 3955 19579 3961
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 20346 3952 20352 4004
rect 20404 3952 20410 4004
rect 20530 3952 20536 4004
rect 20588 3952 20594 4004
rect 20993 3995 21051 4001
rect 20993 3961 21005 3995
rect 21039 3992 21051 3995
rect 21818 3992 21824 4004
rect 21039 3964 21824 3992
rect 21039 3961 21051 3964
rect 20993 3955 21051 3961
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 23768 3992 23796 4023
rect 24486 4020 24492 4072
rect 24544 4060 24550 4072
rect 24964 4069 24992 4100
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 24544 4032 24869 4060
rect 24544 4020 24550 4032
rect 24857 4029 24869 4032
rect 24903 4029 24915 4063
rect 24857 4023 24915 4029
rect 24949 4063 25007 4069
rect 24949 4029 24961 4063
rect 24995 4029 25007 4063
rect 25056 4060 25084 4168
rect 27338 4156 27344 4208
rect 27396 4156 27402 4208
rect 27632 4196 27660 4224
rect 29840 4196 29868 4227
rect 32582 4224 32588 4236
rect 32640 4224 32646 4276
rect 32674 4224 32680 4276
rect 32732 4264 32738 4276
rect 33321 4267 33379 4273
rect 33321 4264 33333 4267
rect 32732 4236 33333 4264
rect 32732 4224 32738 4236
rect 33321 4233 33333 4236
rect 33367 4233 33379 4267
rect 37458 4264 37464 4276
rect 33321 4227 33379 4233
rect 33704 4236 37464 4264
rect 33704 4196 33732 4236
rect 37458 4224 37464 4236
rect 37516 4264 37522 4276
rect 38286 4264 38292 4276
rect 37516 4236 38292 4264
rect 37516 4224 37522 4236
rect 38286 4224 38292 4236
rect 38344 4224 38350 4276
rect 40037 4267 40095 4273
rect 40037 4233 40049 4267
rect 40083 4264 40095 4267
rect 40402 4264 40408 4276
rect 40083 4236 40408 4264
rect 40083 4233 40095 4236
rect 40037 4227 40095 4233
rect 40402 4224 40408 4236
rect 40460 4224 40466 4276
rect 40494 4224 40500 4276
rect 40552 4224 40558 4276
rect 42797 4267 42855 4273
rect 42797 4233 42809 4267
rect 42843 4264 42855 4267
rect 43257 4267 43315 4273
rect 43257 4264 43269 4267
rect 42843 4236 43269 4264
rect 42843 4233 42855 4236
rect 42797 4227 42855 4233
rect 43257 4233 43269 4236
rect 43303 4233 43315 4267
rect 43257 4227 43315 4233
rect 44174 4224 44180 4276
rect 44232 4224 44238 4276
rect 44266 4224 44272 4276
rect 44324 4264 44330 4276
rect 44818 4264 44824 4276
rect 44324 4236 44824 4264
rect 44324 4224 44330 4236
rect 44818 4224 44824 4236
rect 44876 4224 44882 4276
rect 45922 4224 45928 4276
rect 45980 4264 45986 4276
rect 46109 4267 46167 4273
rect 46109 4264 46121 4267
rect 45980 4236 46121 4264
rect 45980 4224 45986 4236
rect 46109 4233 46121 4236
rect 46155 4233 46167 4267
rect 46109 4227 46167 4233
rect 46569 4267 46627 4273
rect 46569 4233 46581 4267
rect 46615 4264 46627 4267
rect 46750 4264 46756 4276
rect 46615 4236 46756 4264
rect 46615 4233 46627 4236
rect 46569 4227 46627 4233
rect 46750 4224 46756 4236
rect 46808 4224 46814 4276
rect 47946 4224 47952 4276
rect 48004 4224 48010 4276
rect 49053 4267 49111 4273
rect 49053 4233 49065 4267
rect 49099 4264 49111 4267
rect 49694 4264 49700 4276
rect 49099 4236 49700 4264
rect 49099 4233 49111 4236
rect 49053 4227 49111 4233
rect 49694 4224 49700 4236
rect 49752 4264 49758 4276
rect 49878 4264 49884 4276
rect 49752 4236 49884 4264
rect 49752 4224 49758 4236
rect 49878 4224 49884 4236
rect 49936 4224 49942 4276
rect 50798 4224 50804 4276
rect 50856 4224 50862 4276
rect 50890 4224 50896 4276
rect 50948 4224 50954 4276
rect 51261 4267 51319 4273
rect 51261 4233 51273 4267
rect 51307 4264 51319 4267
rect 51442 4264 51448 4276
rect 51307 4236 51448 4264
rect 51307 4233 51319 4236
rect 51261 4227 51319 4233
rect 51442 4224 51448 4236
rect 51500 4224 51506 4276
rect 55306 4264 55312 4276
rect 54220 4236 55312 4264
rect 27632 4168 28028 4196
rect 25593 4131 25651 4137
rect 25593 4097 25605 4131
rect 25639 4128 25651 4131
rect 26053 4131 26111 4137
rect 26053 4128 26065 4131
rect 25639 4100 26065 4128
rect 25639 4097 25651 4100
rect 25593 4091 25651 4097
rect 26053 4097 26065 4100
rect 26099 4097 26111 4131
rect 26053 4091 26111 4097
rect 27246 4088 27252 4140
rect 27304 4088 27310 4140
rect 27522 4088 27528 4140
rect 27580 4128 27586 4140
rect 28000 4137 28028 4168
rect 29380 4168 29868 4196
rect 32324 4168 33732 4196
rect 35621 4199 35679 4205
rect 27617 4131 27675 4137
rect 27617 4128 27629 4131
rect 27580 4100 27629 4128
rect 27580 4088 27586 4100
rect 27617 4097 27629 4100
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 27985 4131 28043 4137
rect 27985 4097 27997 4131
rect 28031 4097 28043 4131
rect 27985 4091 28043 4097
rect 28252 4131 28310 4137
rect 28252 4097 28264 4131
rect 28298 4128 28310 4131
rect 28718 4128 28724 4140
rect 28298 4100 28724 4128
rect 28298 4097 28310 4100
rect 28252 4091 28310 4097
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 29380 4128 29408 4168
rect 28868 4100 29408 4128
rect 28868 4088 28874 4100
rect 29454 4088 29460 4140
rect 29512 4088 29518 4140
rect 29638 4088 29644 4140
rect 29696 4128 29702 4140
rect 30009 4131 30067 4137
rect 30009 4128 30021 4131
rect 29696 4100 30021 4128
rect 29696 4088 29702 4100
rect 30009 4097 30021 4100
rect 30055 4097 30067 4131
rect 30009 4091 30067 4097
rect 30742 4088 30748 4140
rect 30800 4088 30806 4140
rect 25685 4063 25743 4069
rect 25685 4060 25697 4063
rect 25056 4032 25697 4060
rect 24949 4023 25007 4029
rect 25685 4029 25697 4032
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 25225 3995 25283 4001
rect 25225 3992 25237 3995
rect 23768 3964 25237 3992
rect 25225 3961 25237 3964
rect 25271 3961 25283 3995
rect 25225 3955 25283 3961
rect 16071 3896 16574 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 18138 3884 18144 3936
rect 18196 3884 18202 3936
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 20548 3924 20576 3952
rect 18371 3896 20576 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 21450 3884 21456 3936
rect 21508 3884 21514 3936
rect 24302 3884 24308 3936
rect 24360 3884 24366 3936
rect 24394 3884 24400 3936
rect 24452 3884 24458 3936
rect 25700 3924 25728 4023
rect 25774 4020 25780 4072
rect 25832 4020 25838 4072
rect 26605 4063 26663 4069
rect 26605 4060 26617 4063
rect 26068 4032 26617 4060
rect 26068 4004 26096 4032
rect 26605 4029 26617 4032
rect 26651 4029 26663 4063
rect 26605 4023 26663 4029
rect 27430 4020 27436 4072
rect 27488 4020 27494 4072
rect 29730 4060 29736 4072
rect 29656 4032 29736 4060
rect 26050 3952 26056 4004
rect 26108 3952 26114 4004
rect 29656 4001 29684 4032
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 30101 4063 30159 4069
rect 30101 4029 30113 4063
rect 30147 4060 30159 4063
rect 30374 4060 30380 4072
rect 30147 4032 30380 4060
rect 30147 4029 30159 4032
rect 30101 4023 30159 4029
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 30834 4020 30840 4072
rect 30892 4069 30898 4072
rect 30892 4063 30941 4069
rect 30892 4029 30895 4063
rect 30929 4029 30941 4063
rect 30892 4023 30941 4029
rect 31021 4063 31079 4069
rect 31021 4029 31033 4063
rect 31067 4060 31079 4063
rect 31067 4032 31248 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 30892 4020 30898 4023
rect 29641 3995 29699 4001
rect 29641 3961 29653 3995
rect 29687 3961 29699 3995
rect 29641 3955 29699 3961
rect 29748 3964 30420 3992
rect 26694 3924 26700 3936
rect 25700 3896 26700 3924
rect 26694 3884 26700 3896
rect 26752 3884 26758 3936
rect 27062 3884 27068 3936
rect 27120 3884 27126 3936
rect 27338 3884 27344 3936
rect 27396 3884 27402 3936
rect 27798 3884 27804 3936
rect 27856 3884 27862 3936
rect 29365 3927 29423 3933
rect 29365 3893 29377 3927
rect 29411 3924 29423 3927
rect 29748 3924 29776 3964
rect 29411 3896 29776 3924
rect 30392 3924 30420 3964
rect 30926 3924 30932 3936
rect 30392 3896 30932 3924
rect 29411 3893 29423 3896
rect 29365 3887 29423 3893
rect 30926 3884 30932 3896
rect 30984 3924 30990 3936
rect 31220 3924 31248 4032
rect 31294 4020 31300 4072
rect 31352 4020 31358 4072
rect 31754 4020 31760 4072
rect 31812 4020 31818 4072
rect 31938 4020 31944 4072
rect 31996 4020 32002 4072
rect 32324 4069 32352 4168
rect 35621 4165 35633 4199
rect 35667 4196 35679 4199
rect 36081 4199 36139 4205
rect 36081 4196 36093 4199
rect 35667 4168 36093 4196
rect 35667 4165 35679 4168
rect 35621 4159 35679 4165
rect 36081 4165 36093 4168
rect 36127 4165 36139 4199
rect 36081 4159 36139 4165
rect 32490 4088 32496 4140
rect 32548 4088 32554 4140
rect 32858 4088 32864 4140
rect 32916 4088 32922 4140
rect 33226 4088 33232 4140
rect 33284 4088 33290 4140
rect 33778 4088 33784 4140
rect 33836 4088 33842 4140
rect 33962 4088 33968 4140
rect 34020 4088 34026 4140
rect 35713 4131 35771 4137
rect 35713 4097 35725 4131
rect 35759 4128 35771 4131
rect 35986 4128 35992 4140
rect 35759 4100 35992 4128
rect 35759 4097 35771 4100
rect 35713 4091 35771 4097
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 36262 4088 36268 4140
rect 36320 4128 36326 4140
rect 36320 4100 36952 4128
rect 36320 4088 36326 4100
rect 32309 4063 32367 4069
rect 32309 4029 32321 4063
rect 32355 4029 32367 4063
rect 32876 4060 32904 4088
rect 32309 4023 32367 4029
rect 32416 4032 32904 4060
rect 33137 4063 33195 4069
rect 31956 3992 31984 4020
rect 32416 3992 32444 4032
rect 33137 4029 33149 4063
rect 33183 4060 33195 4063
rect 33594 4060 33600 4072
rect 33183 4032 33600 4060
rect 33183 4029 33195 4032
rect 33137 4023 33195 4029
rect 33594 4020 33600 4032
rect 33652 4020 33658 4072
rect 33870 4020 33876 4072
rect 33928 4020 33934 4072
rect 34149 4063 34207 4069
rect 34149 4029 34161 4063
rect 34195 4060 34207 4063
rect 34698 4060 34704 4072
rect 34195 4032 34704 4060
rect 34195 4029 34207 4032
rect 34149 4023 34207 4029
rect 34698 4020 34704 4032
rect 34756 4020 34762 4072
rect 35161 4063 35219 4069
rect 35161 4029 35173 4063
rect 35207 4029 35219 4063
rect 35161 4023 35219 4029
rect 31956 3964 32444 3992
rect 32861 3995 32919 4001
rect 32861 3961 32873 3995
rect 32907 3992 32919 3995
rect 33888 3992 33916 4020
rect 32907 3964 33916 3992
rect 35176 3992 35204 4023
rect 35342 4020 35348 4072
rect 35400 4060 35406 4072
rect 35805 4063 35863 4069
rect 35805 4060 35817 4063
rect 35400 4032 35817 4060
rect 35400 4020 35406 4032
rect 35805 4029 35817 4032
rect 35851 4029 35863 4063
rect 35805 4023 35863 4029
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 36633 4063 36691 4069
rect 36633 4060 36645 4063
rect 36136 4032 36645 4060
rect 36136 4020 36142 4032
rect 36633 4029 36645 4032
rect 36679 4060 36691 4063
rect 36814 4060 36820 4072
rect 36679 4032 36820 4060
rect 36679 4029 36691 4032
rect 36633 4023 36691 4029
rect 36814 4020 36820 4032
rect 36872 4020 36878 4072
rect 36924 4060 36952 4100
rect 37090 4088 37096 4140
rect 37148 4088 37154 4140
rect 38197 4131 38255 4137
rect 38197 4128 38209 4131
rect 37200 4100 38209 4128
rect 37200 4060 37228 4100
rect 38197 4097 38209 4100
rect 38243 4097 38255 4131
rect 38197 4091 38255 4097
rect 36924 4032 37228 4060
rect 37826 4020 37832 4072
rect 37884 4020 37890 4072
rect 35253 3995 35311 4001
rect 35253 3992 35265 3995
rect 35176 3964 35265 3992
rect 32907 3961 32919 3964
rect 32861 3955 32919 3961
rect 35253 3961 35265 3964
rect 35299 3961 35311 3995
rect 35253 3955 35311 3961
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 38013 3995 38071 4001
rect 38013 3992 38025 3995
rect 35676 3964 38025 3992
rect 35676 3952 35682 3964
rect 38013 3961 38025 3964
rect 38059 3961 38071 3995
rect 38013 3955 38071 3961
rect 30984 3896 31248 3924
rect 33689 3927 33747 3933
rect 30984 3884 30990 3896
rect 33689 3893 33701 3927
rect 33735 3924 33747 3927
rect 34054 3924 34060 3936
rect 33735 3896 34060 3924
rect 33735 3893 33747 3896
rect 33689 3887 33747 3893
rect 34054 3884 34060 3896
rect 34112 3884 34118 3936
rect 34514 3884 34520 3936
rect 34572 3884 34578 3936
rect 36630 3884 36636 3936
rect 36688 3924 36694 3936
rect 36909 3927 36967 3933
rect 36909 3924 36921 3927
rect 36688 3896 36921 3924
rect 36688 3884 36694 3896
rect 36909 3893 36921 3896
rect 36955 3893 36967 3927
rect 36909 3887 36967 3893
rect 37277 3927 37335 3933
rect 37277 3893 37289 3927
rect 37323 3924 37335 3927
rect 37458 3924 37464 3936
rect 37323 3896 37464 3924
rect 37323 3893 37335 3896
rect 37277 3887 37335 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 38304 3924 38332 4224
rect 38832 4199 38890 4205
rect 38832 4165 38844 4199
rect 38878 4196 38890 4199
rect 39850 4196 39856 4208
rect 38878 4168 39856 4196
rect 38878 4165 38890 4168
rect 38832 4159 38890 4165
rect 39850 4156 39856 4168
rect 39908 4156 39914 4208
rect 40126 4156 40132 4208
rect 40184 4156 40190 4208
rect 41230 4196 41236 4208
rect 40420 4168 41236 4196
rect 38565 4131 38623 4137
rect 38565 4097 38577 4131
rect 38611 4128 38623 4131
rect 38654 4128 38660 4140
rect 38611 4100 38660 4128
rect 38611 4097 38623 4100
rect 38565 4091 38623 4097
rect 38654 4088 38660 4100
rect 38712 4088 38718 4140
rect 40144 4128 40172 4156
rect 40420 4137 40448 4168
rect 41230 4156 41236 4168
rect 41288 4156 41294 4208
rect 41417 4199 41475 4205
rect 41417 4165 41429 4199
rect 41463 4196 41475 4199
rect 42978 4196 42984 4208
rect 41463 4168 42984 4196
rect 41463 4165 41475 4168
rect 41417 4159 41475 4165
rect 42978 4156 42984 4168
rect 43036 4156 43042 4208
rect 44192 4196 44220 4224
rect 44904 4199 44962 4205
rect 44192 4168 44680 4196
rect 44652 4140 44680 4168
rect 44904 4165 44916 4199
rect 44950 4196 44962 4199
rect 45278 4196 45284 4208
rect 44950 4168 45284 4196
rect 44950 4165 44962 4168
rect 44904 4159 44962 4165
rect 45278 4156 45284 4168
rect 45336 4156 45342 4208
rect 48869 4199 48927 4205
rect 46492 4168 47348 4196
rect 40405 4131 40463 4137
rect 40405 4128 40417 4131
rect 40144 4100 40417 4128
rect 40405 4097 40417 4100
rect 40451 4097 40463 4131
rect 40405 4091 40463 4097
rect 40512 4100 41414 4128
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 40512 4060 40540 4100
rect 39632 4032 40540 4060
rect 40589 4063 40647 4069
rect 39632 4020 39638 4032
rect 40589 4029 40601 4063
rect 40635 4029 40647 4063
rect 40589 4023 40647 4029
rect 39945 3995 40003 4001
rect 39945 3961 39957 3995
rect 39991 3992 40003 3995
rect 40218 3992 40224 4004
rect 39991 3964 40224 3992
rect 39991 3961 40003 3964
rect 39945 3955 40003 3961
rect 40218 3952 40224 3964
rect 40276 3952 40282 4004
rect 40604 3992 40632 4023
rect 41046 4020 41052 4072
rect 41104 4020 41110 4072
rect 41386 4060 41414 4100
rect 41598 4088 41604 4140
rect 41656 4128 41662 4140
rect 41785 4131 41843 4137
rect 41785 4128 41797 4131
rect 41656 4100 41797 4128
rect 41656 4088 41662 4100
rect 41785 4097 41797 4100
rect 41831 4097 41843 4131
rect 42061 4131 42119 4137
rect 42061 4128 42073 4131
rect 41785 4091 41843 4097
rect 41892 4100 42073 4128
rect 41892 4060 41920 4100
rect 42061 4097 42073 4100
rect 42107 4097 42119 4131
rect 42061 4091 42119 4097
rect 42444 4100 43760 4128
rect 41386 4032 41920 4060
rect 41969 4063 42027 4069
rect 41969 4029 41981 4063
rect 42015 4060 42027 4063
rect 42150 4060 42156 4072
rect 42015 4032 42156 4060
rect 42015 4029 42027 4032
rect 41969 4023 42027 4029
rect 42150 4020 42156 4032
rect 42208 4060 42214 4072
rect 42444 4060 42472 4100
rect 42208 4032 42472 4060
rect 42208 4020 42214 4032
rect 42610 4020 42616 4072
rect 42668 4020 42674 4072
rect 42705 4063 42763 4069
rect 42705 4029 42717 4063
rect 42751 4029 42763 4063
rect 43732 4060 43760 4100
rect 43806 4088 43812 4140
rect 43864 4088 43870 4140
rect 44266 4088 44272 4140
rect 44324 4088 44330 4140
rect 44361 4131 44419 4137
rect 44361 4097 44373 4131
rect 44407 4097 44419 4131
rect 44361 4091 44419 4097
rect 44284 4060 44312 4088
rect 43732 4032 44312 4060
rect 44376 4060 44404 4091
rect 44634 4088 44640 4140
rect 44692 4088 44698 4140
rect 45186 4128 45192 4140
rect 44744 4100 45192 4128
rect 44744 4060 44772 4100
rect 45186 4088 45192 4100
rect 45244 4088 45250 4140
rect 46198 4088 46204 4140
rect 46256 4128 46262 4140
rect 46492 4137 46520 4168
rect 46477 4131 46535 4137
rect 46477 4128 46489 4131
rect 46256 4100 46489 4128
rect 46256 4088 46262 4100
rect 46477 4097 46489 4100
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 46584 4100 46796 4128
rect 44376 4032 44772 4060
rect 42705 4023 42763 4029
rect 42720 3992 42748 4023
rect 45738 4020 45744 4072
rect 45796 4060 45802 4072
rect 46584 4060 46612 4100
rect 45796 4032 46612 4060
rect 45796 4020 45802 4032
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 46768 4060 46796 4100
rect 47210 4088 47216 4140
rect 47268 4088 47274 4140
rect 47320 4128 47348 4168
rect 48869 4165 48881 4199
rect 48915 4196 48927 4199
rect 49786 4196 49792 4208
rect 48915 4168 49792 4196
rect 48915 4165 48927 4168
rect 48869 4159 48927 4165
rect 49786 4156 49792 4168
rect 49844 4156 49850 4208
rect 50188 4199 50246 4205
rect 50188 4165 50200 4199
rect 50234 4196 50246 4199
rect 50908 4196 50936 4224
rect 50234 4168 50936 4196
rect 53101 4199 53159 4205
rect 50234 4165 50246 4168
rect 50188 4159 50246 4165
rect 53101 4165 53113 4199
rect 53147 4196 53159 4199
rect 53926 4196 53932 4208
rect 53147 4168 53932 4196
rect 53147 4165 53159 4168
rect 53101 4159 53159 4165
rect 53926 4156 53932 4168
rect 53984 4156 53990 4208
rect 48406 4128 48412 4140
rect 47320 4100 48412 4128
rect 48406 4088 48412 4100
rect 48464 4088 48470 4140
rect 48590 4088 48596 4140
rect 48648 4088 48654 4140
rect 49602 4128 49608 4140
rect 48700 4100 49608 4128
rect 46768 4032 47440 4060
rect 40512 3964 40632 3992
rect 41386 3964 42748 3992
rect 43165 3995 43223 4001
rect 40310 3924 40316 3936
rect 38304 3896 40316 3924
rect 40310 3884 40316 3896
rect 40368 3924 40374 3936
rect 40512 3924 40540 3964
rect 40368 3896 40540 3924
rect 40368 3884 40374 3896
rect 41230 3884 41236 3936
rect 41288 3924 41294 3936
rect 41386 3924 41414 3964
rect 43165 3961 43177 3995
rect 43211 3992 43223 3995
rect 44450 3992 44456 4004
rect 43211 3964 44456 3992
rect 43211 3961 43223 3964
rect 43165 3955 43223 3961
rect 44450 3952 44456 3964
rect 44508 3952 44514 4004
rect 45830 3952 45836 4004
rect 45888 3952 45894 4004
rect 46017 3995 46075 4001
rect 46017 3961 46029 3995
rect 46063 3992 46075 3995
rect 47302 3992 47308 4004
rect 46063 3964 47308 3992
rect 46063 3961 46075 3964
rect 46017 3955 46075 3961
rect 47302 3952 47308 3964
rect 47360 3952 47366 4004
rect 47412 3992 47440 4032
rect 47578 4020 47584 4072
rect 47636 4060 47642 4072
rect 47673 4063 47731 4069
rect 47673 4060 47685 4063
rect 47636 4032 47685 4060
rect 47636 4020 47642 4032
rect 47673 4029 47685 4032
rect 47719 4029 47731 4063
rect 47673 4023 47731 4029
rect 47854 4020 47860 4072
rect 47912 4020 47918 4072
rect 48424 4060 48452 4088
rect 48700 4060 48728 4100
rect 49602 4088 49608 4100
rect 49660 4088 49666 4140
rect 50338 4088 50344 4140
rect 50396 4128 50402 4140
rect 50433 4131 50491 4137
rect 50433 4128 50445 4131
rect 50396 4100 50445 4128
rect 50396 4088 50402 4100
rect 50433 4097 50445 4100
rect 50479 4097 50491 4131
rect 50433 4091 50491 4097
rect 50522 4088 50528 4140
rect 50580 4128 50586 4140
rect 50893 4131 50951 4137
rect 50893 4128 50905 4131
rect 50580 4100 50905 4128
rect 50580 4088 50586 4100
rect 50893 4097 50905 4100
rect 50939 4097 50951 4131
rect 50893 4091 50951 4097
rect 51258 4088 51264 4140
rect 51316 4128 51322 4140
rect 51629 4131 51687 4137
rect 51629 4128 51641 4131
rect 51316 4100 51641 4128
rect 51316 4088 51322 4100
rect 51629 4097 51641 4100
rect 51675 4097 51687 4131
rect 51629 4091 51687 4097
rect 52549 4131 52607 4137
rect 52549 4097 52561 4131
rect 52595 4128 52607 4131
rect 52730 4128 52736 4140
rect 52595 4100 52736 4128
rect 52595 4097 52607 4100
rect 52549 4091 52607 4097
rect 52730 4088 52736 4100
rect 52788 4088 52794 4140
rect 53837 4131 53895 4137
rect 53837 4097 53849 4131
rect 53883 4128 53895 4131
rect 54220 4128 54248 4236
rect 55306 4224 55312 4236
rect 55364 4224 55370 4276
rect 55490 4224 55496 4276
rect 55548 4264 55554 4276
rect 56045 4267 56103 4273
rect 56045 4264 56057 4267
rect 55548 4236 56057 4264
rect 55548 4224 55554 4236
rect 56045 4233 56057 4236
rect 56091 4233 56103 4267
rect 56045 4227 56103 4233
rect 56410 4224 56416 4276
rect 56468 4264 56474 4276
rect 57241 4267 57299 4273
rect 57241 4264 57253 4267
rect 56468 4236 57253 4264
rect 56468 4224 56474 4236
rect 57241 4233 57253 4236
rect 57287 4233 57299 4267
rect 57241 4227 57299 4233
rect 55858 4156 55864 4208
rect 55916 4196 55922 4208
rect 55916 4168 56456 4196
rect 55916 4156 55922 4168
rect 53883 4100 54248 4128
rect 53883 4097 53895 4100
rect 53837 4091 53895 4097
rect 54754 4088 54760 4140
rect 54812 4088 54818 4140
rect 55950 4088 55956 4140
rect 56008 4088 56014 4140
rect 56428 4137 56456 4168
rect 56962 4156 56968 4208
rect 57020 4196 57026 4208
rect 57149 4199 57207 4205
rect 57149 4196 57161 4199
rect 57020 4168 57161 4196
rect 57020 4156 57026 4168
rect 57149 4165 57161 4168
rect 57195 4165 57207 4199
rect 57149 4159 57207 4165
rect 56413 4131 56471 4137
rect 56413 4097 56425 4131
rect 56459 4097 56471 4131
rect 56413 4091 56471 4097
rect 48424 4032 48728 4060
rect 48777 4063 48835 4069
rect 48777 4029 48789 4063
rect 48823 4029 48835 4063
rect 48777 4023 48835 4029
rect 50709 4063 50767 4069
rect 50709 4029 50721 4063
rect 50755 4060 50767 4063
rect 51074 4060 51080 4072
rect 50755 4032 51080 4060
rect 50755 4029 50767 4032
rect 50709 4023 50767 4029
rect 48409 3995 48467 4001
rect 48409 3992 48421 3995
rect 47412 3964 48421 3992
rect 48409 3961 48421 3964
rect 48455 3961 48467 3995
rect 48792 3992 48820 4023
rect 51074 4020 51080 4032
rect 51132 4020 51138 4072
rect 51445 4063 51503 4069
rect 51445 4029 51457 4063
rect 51491 4029 51503 4063
rect 51445 4023 51503 4029
rect 51813 4063 51871 4069
rect 51813 4029 51825 4063
rect 51859 4060 51871 4063
rect 52638 4060 52644 4072
rect 51859 4032 52644 4060
rect 51859 4029 51871 4032
rect 51813 4023 51871 4029
rect 51460 3992 51488 4023
rect 52638 4020 52644 4032
rect 52696 4020 52702 4072
rect 52914 4020 52920 4072
rect 52972 4020 52978 4072
rect 53009 4063 53067 4069
rect 53009 4029 53021 4063
rect 53055 4060 53067 4063
rect 53098 4060 53104 4072
rect 53055 4032 53104 4060
rect 53055 4029 53067 4032
rect 53009 4023 53067 4029
rect 53098 4020 53104 4032
rect 53156 4020 53162 4072
rect 53653 4063 53711 4069
rect 53653 4060 53665 4063
rect 53208 4032 53665 4060
rect 52546 3992 52552 4004
rect 48792 3964 49556 3992
rect 51460 3964 52552 3992
rect 48409 3955 48467 3961
rect 41288 3896 41414 3924
rect 41288 3884 41294 3896
rect 41598 3884 41604 3936
rect 41656 3884 41662 3936
rect 42242 3884 42248 3936
rect 42300 3884 42306 3936
rect 44545 3927 44603 3933
rect 44545 3893 44557 3927
rect 44591 3924 44603 3927
rect 45278 3924 45284 3936
rect 44591 3896 45284 3924
rect 44591 3893 44603 3896
rect 44545 3887 44603 3893
rect 45278 3884 45284 3896
rect 45336 3884 45342 3936
rect 45848 3924 45876 3952
rect 47029 3927 47087 3933
rect 47029 3924 47041 3927
rect 45848 3896 47041 3924
rect 47029 3893 47041 3896
rect 47075 3893 47087 3927
rect 47029 3887 47087 3893
rect 48314 3884 48320 3936
rect 48372 3884 48378 3936
rect 48682 3884 48688 3936
rect 48740 3884 48746 3936
rect 49528 3924 49556 3964
rect 52546 3952 52552 3964
rect 52604 3992 52610 4004
rect 53208 3992 53236 4032
rect 53653 4029 53665 4032
rect 53699 4060 53711 4063
rect 54018 4060 54024 4072
rect 53699 4032 54024 4060
rect 53699 4029 53711 4032
rect 53653 4023 53711 4029
rect 54018 4020 54024 4032
rect 54076 4020 54082 4072
rect 54110 4020 54116 4072
rect 54168 4020 54174 4072
rect 54846 4020 54852 4072
rect 54904 4069 54910 4072
rect 54904 4063 54953 4069
rect 54904 4029 54907 4063
rect 54941 4029 54953 4063
rect 54904 4023 54953 4029
rect 54904 4020 54910 4023
rect 55030 4020 55036 4072
rect 55088 4020 55094 4072
rect 55309 4063 55367 4069
rect 55309 4029 55321 4063
rect 55355 4060 55367 4063
rect 55582 4060 55588 4072
rect 55355 4032 55588 4060
rect 55355 4029 55367 4032
rect 55309 4023 55367 4029
rect 55582 4020 55588 4032
rect 55640 4020 55646 4072
rect 55766 4020 55772 4072
rect 55824 4060 55830 4072
rect 56505 4063 56563 4069
rect 55824 4032 55996 4060
rect 55824 4020 55830 4032
rect 52604 3964 53236 3992
rect 53469 3995 53527 4001
rect 52604 3952 52610 3964
rect 53469 3961 53481 3995
rect 53515 3992 53527 3995
rect 54128 3992 54156 4020
rect 55968 4004 55996 4032
rect 56505 4029 56517 4063
rect 56551 4029 56563 4063
rect 56505 4023 56563 4029
rect 53515 3964 54156 3992
rect 53515 3961 53527 3964
rect 53469 3955 53527 3961
rect 55950 3952 55956 4004
rect 56008 3952 56014 4004
rect 49694 3924 49700 3936
rect 49528 3896 49700 3924
rect 49694 3884 49700 3896
rect 49752 3884 49758 3936
rect 51902 3884 51908 3936
rect 51960 3884 51966 3936
rect 54018 3884 54024 3936
rect 54076 3884 54082 3936
rect 54113 3927 54171 3933
rect 54113 3893 54125 3927
rect 54159 3924 54171 3927
rect 56520 3924 56548 4023
rect 56686 4020 56692 4072
rect 56744 4020 56750 4072
rect 57057 4063 57115 4069
rect 57057 4029 57069 4063
rect 57103 4060 57115 4063
rect 57238 4060 57244 4072
rect 57103 4032 57244 4060
rect 57103 4029 57115 4032
rect 57057 4023 57115 4029
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 58437 4063 58495 4069
rect 58437 4029 58449 4063
rect 58483 4029 58495 4063
rect 58437 4023 58495 4029
rect 57609 3995 57667 4001
rect 57609 3961 57621 3995
rect 57655 3992 57667 3995
rect 58452 3992 58480 4023
rect 57655 3964 58480 3992
rect 57655 3961 57667 3964
rect 57609 3955 57667 3961
rect 54159 3896 56548 3924
rect 54159 3893 54171 3896
rect 54113 3887 54171 3893
rect 57514 3884 57520 3936
rect 57572 3924 57578 3936
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 57572 3896 57897 3924
rect 57572 3884 57578 3896
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 1104 3834 58880 3856
rect 1104 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 22616 3834
rect 22668 3782 22680 3834
rect 22732 3782 22744 3834
rect 22796 3782 22808 3834
rect 22860 3782 22872 3834
rect 22924 3782 37060 3834
rect 37112 3782 37124 3834
rect 37176 3782 37188 3834
rect 37240 3782 37252 3834
rect 37304 3782 37316 3834
rect 37368 3782 51504 3834
rect 51556 3782 51568 3834
rect 51620 3782 51632 3834
rect 51684 3782 51696 3834
rect 51748 3782 51760 3834
rect 51812 3782 58880 3834
rect 1104 3760 58880 3782
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3559 3692 6684 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3652 2007 3655
rect 4154 3652 4160 3664
rect 1995 3624 4160 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 5350 3612 5356 3664
rect 5408 3612 5414 3664
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 6089 3655 6147 3661
rect 6089 3652 6101 3655
rect 5500 3624 6101 3652
rect 5500 3612 5506 3624
rect 6089 3621 6101 3624
rect 6135 3621 6147 3655
rect 6089 3615 6147 3621
rect 2130 3544 2136 3596
rect 2188 3544 2194 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3142 3584 3148 3596
rect 3007 3556 3148 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 4614 3584 4620 3596
rect 3292 3556 4620 3584
rect 3292 3544 3298 3556
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4798 3544 4804 3596
rect 4856 3544 4862 3596
rect 4890 3544 4896 3596
rect 4948 3593 4954 3596
rect 5074 3593 5080 3596
rect 4948 3587 4997 3593
rect 4948 3553 4951 3587
rect 4985 3553 4997 3587
rect 4948 3547 4997 3553
rect 5058 3587 5080 3593
rect 5058 3553 5070 3587
rect 5058 3547 5080 3553
rect 4948 3544 4954 3547
rect 5074 3544 5080 3547
rect 5132 3544 5138 3596
rect 6656 3593 6684 3692
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 6880 3692 7849 3720
rect 6880 3680 6886 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 8220 3692 10548 3720
rect 6748 3652 6776 3680
rect 8220 3664 8248 3692
rect 7009 3655 7067 3661
rect 7009 3652 7021 3655
rect 6748 3624 7021 3652
rect 7009 3621 7021 3624
rect 7055 3621 7067 3655
rect 7009 3615 7067 3621
rect 7098 3612 7104 3664
rect 7156 3652 7162 3664
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 7156 3624 7481 3652
rect 7156 3612 7162 3624
rect 7469 3621 7481 3624
rect 7515 3652 7527 3655
rect 8202 3652 8208 3664
rect 7515 3624 8208 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 10520 3652 10548 3692
rect 10594 3680 10600 3732
rect 10652 3680 10658 3732
rect 13538 3680 13544 3732
rect 13596 3680 13602 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 15657 3723 15715 3729
rect 14148 3692 15608 3720
rect 14148 3680 14154 3692
rect 11238 3652 11244 3664
rect 9723 3624 10364 3652
rect 10520 3624 11244 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 6641 3587 6699 3593
rect 5859 3556 6592 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3510 3516 3516 3528
rect 3099 3488 3516 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 5902 3476 5908 3528
rect 5960 3516 5966 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5960 3488 6009 3516
rect 5960 3476 5966 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 6564 3516 6592 3556
rect 6641 3553 6653 3587
rect 6687 3553 6699 3587
rect 7926 3584 7932 3596
rect 6641 3547 6699 3553
rect 7300 3556 7932 3584
rect 7300 3516 7328 3556
rect 7926 3544 7932 3556
rect 7984 3584 7990 3596
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7984 3556 8125 3584
rect 7984 3544 7990 3556
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 9030 3544 9036 3596
rect 9088 3544 9094 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 10336 3593 10364 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 13556 3652 13584 3680
rect 12406 3624 13584 3652
rect 15013 3655 15071 3661
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 9180 3556 9229 3584
rect 9180 3544 9186 3556
rect 9217 3553 9229 3556
rect 9263 3553 9275 3587
rect 9217 3547 9275 3553
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3553 10379 3587
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 10321 3547 10379 3553
rect 11348 3556 12265 3584
rect 6564 3488 7328 3516
rect 5997 3479 6055 3485
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 10778 3476 10784 3528
rect 10836 3476 10842 3528
rect 2685 3451 2743 3457
rect 2685 3417 2697 3451
rect 2731 3448 2743 3451
rect 3145 3451 3203 3457
rect 3145 3448 3157 3451
rect 2731 3420 3157 3448
rect 2731 3417 2743 3420
rect 2685 3411 2743 3417
rect 3145 3417 3157 3420
rect 3191 3417 3203 3451
rect 3145 3411 3203 3417
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3476 3420 3893 3448
rect 3476 3408 3482 3420
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 7282 3408 7288 3460
rect 7340 3408 7346 3460
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 8803 3420 9321 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 11348 3392 11376 3556
rect 12253 3553 12265 3556
rect 12299 3584 12311 3587
rect 12406 3584 12434 3624
rect 15013 3621 15025 3655
rect 15059 3621 15071 3655
rect 15580 3652 15608 3692
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 15746 3720 15752 3732
rect 15703 3692 15752 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16209 3723 16267 3729
rect 16209 3689 16221 3723
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 16224 3652 16252 3683
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16448 3692 17356 3720
rect 16448 3680 16454 3692
rect 17328 3652 17356 3692
rect 17402 3680 17408 3732
rect 17460 3680 17466 3732
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 17920 3692 20852 3720
rect 17920 3680 17926 3692
rect 20346 3652 20352 3664
rect 15580 3624 16252 3652
rect 16408 3624 17264 3652
rect 17328 3624 20352 3652
rect 15013 3615 15071 3621
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 12299 3556 12434 3584
rect 12820 3556 13277 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12820 3528 12848 3556
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 15028 3584 15056 3615
rect 16408 3593 16436 3624
rect 16393 3587 16451 3593
rect 15028 3556 16252 3584
rect 13265 3547 13323 3553
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 12802 3476 12808 3528
rect 12860 3476 12866 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 13004 3448 13032 3479
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14056 3488 14657 3516
rect 14056 3476 14062 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 15252 3488 15301 3516
rect 15252 3476 15258 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 15838 3476 15844 3528
rect 15896 3476 15902 3528
rect 16224 3525 16252 3556
rect 16393 3553 16405 3587
rect 16439 3553 16451 3587
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16393 3547 16451 3553
rect 16500 3556 16865 3584
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16500 3516 16528 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 17236 3584 17264 3624
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 18782 3584 18788 3596
rect 17236 3556 18788 3584
rect 16853 3547 16911 3553
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 20824 3593 20852 3692
rect 22278 3680 22284 3732
rect 22336 3720 22342 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 22336 3692 22937 3720
rect 22336 3680 22342 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 24762 3720 24768 3732
rect 22925 3683 22983 3689
rect 24596 3692 24768 3720
rect 21453 3655 21511 3661
rect 21453 3621 21465 3655
rect 21499 3652 21511 3655
rect 21499 3624 22140 3652
rect 21499 3621 21511 3624
rect 21453 3615 21511 3621
rect 22112 3593 22140 3624
rect 22480 3624 23796 3652
rect 19705 3587 19763 3593
rect 19705 3584 19717 3587
rect 19208 3556 19717 3584
rect 19208 3544 19214 3556
rect 19705 3553 19717 3556
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 22097 3587 22155 3593
rect 22097 3553 22109 3587
rect 22143 3553 22155 3587
rect 22097 3547 22155 3553
rect 16209 3479 16267 3485
rect 16408 3488 16528 3516
rect 15396 3448 15424 3476
rect 16408 3448 16436 3488
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16632 3488 16773 3516
rect 16632 3476 16638 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 18322 3476 18328 3528
rect 18380 3476 18386 3528
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 19058 3516 19064 3528
rect 19015 3488 19064 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 11480 3420 13032 3448
rect 13832 3420 16436 3448
rect 16485 3451 16543 3457
rect 11480 3408 11486 3420
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4062 3380 4068 3392
rect 4019 3352 4068 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 6914 3380 6920 3392
rect 4203 3352 6920 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 9766 3340 9772 3392
rect 9824 3340 9830 3392
rect 10870 3340 10876 3392
rect 10928 3340 10934 3392
rect 11330 3340 11336 3392
rect 11388 3340 11394 3392
rect 11698 3340 11704 3392
rect 11756 3340 11762 3392
rect 12434 3340 12440 3392
rect 12492 3340 12498 3392
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 13832 3380 13860 3420
rect 16485 3417 16497 3451
rect 16531 3417 16543 3451
rect 18984 3448 19012 3479
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 19334 3476 19340 3528
rect 19392 3476 19398 3528
rect 20254 3476 20260 3528
rect 20312 3516 20318 3528
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20312 3488 21005 3516
rect 20312 3476 20318 3488
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 20993 3479 21051 3485
rect 21082 3476 21088 3528
rect 21140 3476 21146 3528
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 22281 3519 22339 3525
rect 21416 3512 22232 3516
rect 22281 3512 22293 3519
rect 21416 3488 22293 3512
rect 21416 3476 21422 3488
rect 22204 3485 22293 3488
rect 22327 3485 22339 3519
rect 22204 3484 22339 3485
rect 22281 3479 22339 3484
rect 16485 3411 16543 3417
rect 18248 3420 19012 3448
rect 12768 3352 13860 3380
rect 12768 3340 12774 3352
rect 13906 3340 13912 3392
rect 13964 3340 13970 3392
rect 14090 3340 14096 3392
rect 14148 3340 14154 3392
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15194 3380 15200 3392
rect 15151 3352 15200 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 16022 3340 16028 3392
rect 16080 3340 16086 3392
rect 16500 3380 16528 3411
rect 18248 3392 18276 3420
rect 21450 3408 21456 3460
rect 21508 3448 21514 3460
rect 22480 3448 22508 3624
rect 23474 3544 23480 3596
rect 23532 3544 23538 3596
rect 23768 3593 23796 3624
rect 24596 3593 24624 3692
rect 24762 3680 24768 3692
rect 24820 3680 24826 3732
rect 25961 3723 26019 3729
rect 25961 3689 25973 3723
rect 26007 3720 26019 3723
rect 26050 3720 26056 3732
rect 26007 3692 26056 3720
rect 26007 3689 26019 3692
rect 25961 3683 26019 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 26694 3720 26700 3732
rect 26283 3692 26700 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 26694 3680 26700 3692
rect 26752 3680 26758 3732
rect 28718 3680 28724 3732
rect 28776 3680 28782 3732
rect 29454 3720 29460 3732
rect 28828 3692 29460 3720
rect 27893 3655 27951 3661
rect 27893 3621 27905 3655
rect 27939 3652 27951 3655
rect 28828 3652 28856 3692
rect 29454 3680 29460 3692
rect 29512 3680 29518 3732
rect 30926 3680 30932 3732
rect 30984 3680 30990 3732
rect 36078 3680 36084 3732
rect 36136 3680 36142 3732
rect 36170 3680 36176 3732
rect 36228 3720 36234 3732
rect 37645 3723 37703 3729
rect 36228 3692 37596 3720
rect 36228 3680 36234 3692
rect 29549 3655 29607 3661
rect 29549 3652 29561 3655
rect 27939 3624 28856 3652
rect 29380 3624 29561 3652
rect 27939 3621 27951 3624
rect 27893 3615 27951 3621
rect 29380 3593 29408 3624
rect 29549 3621 29561 3624
rect 29595 3621 29607 3655
rect 29549 3615 29607 3621
rect 23753 3587 23811 3593
rect 23753 3553 23765 3587
rect 23799 3584 23811 3587
rect 24581 3587 24639 3593
rect 23799 3556 24532 3584
rect 23799 3553 23811 3556
rect 23753 3547 23811 3553
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 23014 3516 23020 3528
rect 22603 3488 23020 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23937 3519 23995 3525
rect 23937 3485 23949 3519
rect 23983 3516 23995 3519
rect 24394 3516 24400 3528
rect 23983 3488 24400 3516
rect 23983 3485 23995 3488
rect 23937 3479 23995 3485
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 24504 3516 24532 3556
rect 24581 3553 24593 3587
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3584 26755 3587
rect 29365 3587 29423 3593
rect 26743 3556 29316 3584
rect 26743 3553 26755 3556
rect 26697 3547 26755 3553
rect 25222 3516 25228 3528
rect 24504 3488 25228 3516
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 27157 3519 27215 3525
rect 27157 3485 27169 3519
rect 27203 3485 27215 3519
rect 27157 3479 27215 3485
rect 27341 3519 27399 3525
rect 27341 3485 27353 3519
rect 27387 3485 27399 3519
rect 27341 3479 27399 3485
rect 28077 3519 28135 3525
rect 28077 3485 28089 3519
rect 28123 3516 28135 3519
rect 29288 3516 29316 3556
rect 29365 3553 29377 3587
rect 29411 3553 29423 3587
rect 29365 3547 29423 3553
rect 30098 3544 30104 3596
rect 30156 3544 30162 3596
rect 30944 3593 30972 3680
rect 31754 3612 31760 3664
rect 31812 3652 31818 3664
rect 37568 3652 37596 3692
rect 37645 3689 37657 3723
rect 37691 3720 37703 3723
rect 37826 3720 37832 3732
rect 37691 3692 37832 3720
rect 37691 3689 37703 3692
rect 37645 3683 37703 3689
rect 37826 3680 37832 3692
rect 37884 3680 37890 3732
rect 37918 3680 37924 3732
rect 37976 3720 37982 3732
rect 42150 3720 42156 3732
rect 37976 3692 42156 3720
rect 37976 3680 37982 3692
rect 42150 3680 42156 3692
rect 42208 3680 42214 3732
rect 42886 3680 42892 3732
rect 42944 3680 42950 3732
rect 42978 3680 42984 3732
rect 43036 3680 43042 3732
rect 45738 3720 45744 3732
rect 43548 3692 45744 3720
rect 40589 3655 40647 3661
rect 31812 3624 33548 3652
rect 37568 3624 39068 3652
rect 31812 3612 31818 3624
rect 30929 3587 30987 3593
rect 30929 3553 30941 3587
rect 30975 3553 30987 3587
rect 30929 3547 30987 3553
rect 32030 3544 32036 3596
rect 32088 3584 32094 3596
rect 32217 3587 32275 3593
rect 32217 3584 32229 3587
rect 32088 3556 32229 3584
rect 32088 3544 32094 3556
rect 32217 3553 32229 3556
rect 32263 3553 32275 3587
rect 32217 3547 32275 3553
rect 32490 3544 32496 3596
rect 32548 3544 32554 3596
rect 33520 3593 33548 3624
rect 33505 3587 33563 3593
rect 33505 3553 33517 3587
rect 33551 3553 33563 3587
rect 33505 3547 33563 3553
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 33965 3587 34023 3593
rect 33965 3584 33977 3587
rect 33652 3556 33977 3584
rect 33652 3544 33658 3556
rect 33965 3553 33977 3556
rect 34011 3584 34023 3587
rect 34011 3556 34744 3584
rect 34011 3553 34023 3556
rect 33965 3547 34023 3553
rect 30116 3516 30144 3544
rect 28123 3488 29132 3516
rect 29288 3488 30144 3516
rect 28123 3485 28135 3488
rect 28077 3479 28135 3485
rect 21508 3420 22508 3448
rect 22756 3420 24256 3448
rect 21508 3408 21514 3420
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16500 3352 16589 3380
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 17218 3340 17224 3392
rect 17276 3340 17282 3392
rect 17678 3340 17684 3392
rect 17736 3340 17742 3392
rect 18230 3340 18236 3392
rect 18288 3340 18294 3392
rect 18414 3340 18420 3392
rect 18472 3340 18478 3392
rect 21542 3340 21548 3392
rect 21600 3340 21606 3392
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3380 22523 3383
rect 22646 3380 22652 3392
rect 22511 3352 22652 3380
rect 22511 3349 22523 3352
rect 22465 3343 22523 3349
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 22756 3389 22784 3420
rect 22741 3383 22799 3389
rect 22741 3349 22753 3383
rect 22787 3349 22799 3383
rect 22741 3343 22799 3349
rect 24118 3340 24124 3392
rect 24176 3340 24182 3392
rect 24228 3380 24256 3420
rect 24302 3408 24308 3460
rect 24360 3448 24366 3460
rect 24826 3451 24884 3457
rect 24826 3448 24838 3451
rect 24360 3420 24838 3448
rect 24360 3408 24366 3420
rect 24826 3417 24838 3420
rect 24872 3417 24884 3451
rect 26145 3451 26203 3457
rect 26145 3448 26157 3451
rect 24826 3411 24884 3417
rect 24964 3420 26157 3448
rect 24964 3380 24992 3420
rect 26145 3417 26157 3420
rect 26191 3417 26203 3451
rect 27172 3448 27200 3479
rect 26145 3411 26203 3417
rect 26252 3420 27200 3448
rect 27356 3448 27384 3479
rect 29104 3460 29132 3488
rect 31294 3476 31300 3528
rect 31352 3476 31358 3528
rect 31938 3476 31944 3528
rect 31996 3476 32002 3528
rect 32401 3519 32459 3525
rect 32401 3485 32413 3519
rect 32447 3516 32459 3519
rect 32508 3516 32536 3544
rect 34057 3519 34115 3525
rect 34057 3516 34069 3519
rect 32447 3488 34069 3516
rect 32447 3485 32459 3488
rect 32401 3479 32459 3485
rect 34057 3485 34069 3488
rect 34103 3485 34115 3519
rect 34057 3479 34115 3485
rect 28534 3448 28540 3460
rect 27356 3420 28540 3448
rect 24228 3352 24992 3380
rect 25222 3340 25228 3392
rect 25280 3380 25286 3392
rect 25774 3380 25780 3392
rect 25280 3352 25780 3380
rect 25280 3340 25286 3352
rect 25774 3340 25780 3352
rect 25832 3380 25838 3392
rect 26252 3380 26280 3420
rect 25832 3352 26280 3380
rect 25832 3340 25838 3352
rect 26786 3340 26792 3392
rect 26844 3340 26850 3392
rect 27172 3380 27200 3420
rect 28534 3408 28540 3420
rect 28592 3408 28598 3460
rect 29086 3408 29092 3460
rect 29144 3408 29150 3460
rect 29917 3451 29975 3457
rect 29917 3417 29929 3451
rect 29963 3448 29975 3451
rect 32416 3448 32444 3479
rect 34514 3476 34520 3528
rect 34572 3476 34578 3528
rect 34716 3525 34744 3556
rect 38102 3544 38108 3596
rect 38160 3544 38166 3596
rect 38289 3587 38347 3593
rect 38289 3553 38301 3587
rect 38335 3584 38347 3587
rect 38378 3584 38384 3596
rect 38335 3556 38384 3584
rect 38335 3553 38347 3556
rect 38289 3547 38347 3553
rect 38378 3544 38384 3556
rect 38436 3544 38442 3596
rect 38470 3544 38476 3596
rect 38528 3584 38534 3596
rect 39040 3593 39068 3624
rect 40589 3621 40601 3655
rect 40635 3652 40647 3655
rect 42058 3652 42064 3664
rect 40635 3624 41276 3652
rect 40635 3621 40647 3624
rect 40589 3615 40647 3621
rect 39025 3587 39083 3593
rect 38528 3556 38792 3584
rect 38528 3544 38534 3556
rect 34701 3519 34759 3525
rect 34701 3485 34713 3519
rect 34747 3516 34759 3519
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 34747 3488 37565 3516
rect 34747 3485 34759 3488
rect 34701 3479 34759 3485
rect 37553 3485 37565 3488
rect 37599 3516 37611 3519
rect 37642 3516 37648 3528
rect 37599 3488 37648 3516
rect 37599 3485 37611 3488
rect 37553 3479 37611 3485
rect 37642 3476 37648 3488
rect 37700 3516 37706 3528
rect 38654 3516 38660 3528
rect 37700 3488 38660 3516
rect 37700 3476 37706 3488
rect 38654 3476 38660 3488
rect 38712 3476 38718 3528
rect 38764 3516 38792 3556
rect 39025 3553 39037 3587
rect 39071 3553 39083 3587
rect 39025 3547 39083 3553
rect 39942 3544 39948 3596
rect 40000 3544 40006 3596
rect 40126 3544 40132 3596
rect 40184 3544 40190 3596
rect 41248 3593 41276 3624
rect 41386 3624 42064 3652
rect 41233 3587 41291 3593
rect 41233 3553 41245 3587
rect 41279 3553 41291 3587
rect 41233 3547 41291 3553
rect 39209 3519 39267 3525
rect 39209 3516 39221 3519
rect 38764 3488 39221 3516
rect 39209 3485 39221 3488
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 29963 3420 32444 3448
rect 32493 3451 32551 3457
rect 29963 3417 29975 3420
rect 29917 3411 29975 3417
rect 32493 3417 32505 3451
rect 32539 3448 32551 3451
rect 32953 3451 33011 3457
rect 32953 3448 32965 3451
rect 32539 3420 32965 3448
rect 32539 3417 32551 3420
rect 32493 3411 32551 3417
rect 32953 3417 32965 3420
rect 32999 3417 33011 3451
rect 32953 3411 33011 3417
rect 28258 3380 28264 3392
rect 27172 3352 28264 3380
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 28629 3383 28687 3389
rect 28629 3349 28641 3383
rect 28675 3380 28687 3383
rect 29270 3380 29276 3392
rect 28675 3352 29276 3380
rect 28675 3349 28687 3352
rect 28629 3343 28687 3349
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 29730 3380 29736 3392
rect 29420 3352 29736 3380
rect 29420 3340 29426 3352
rect 29730 3340 29736 3352
rect 29788 3380 29794 3392
rect 29932 3380 29960 3411
rect 33226 3408 33232 3460
rect 33284 3448 33290 3460
rect 34241 3451 34299 3457
rect 34241 3448 34253 3451
rect 33284 3420 34253 3448
rect 33284 3408 33290 3420
rect 34241 3417 34253 3420
rect 34287 3417 34299 3451
rect 34532 3448 34560 3476
rect 34946 3451 35004 3457
rect 34946 3448 34958 3451
rect 34532 3420 34958 3448
rect 34241 3411 34299 3417
rect 34946 3417 34958 3420
rect 34992 3417 35004 3451
rect 34946 3411 35004 3417
rect 37308 3451 37366 3457
rect 37308 3417 37320 3451
rect 37354 3448 37366 3451
rect 37458 3448 37464 3460
rect 37354 3420 37464 3448
rect 37354 3417 37366 3420
rect 37308 3411 37366 3417
rect 37458 3408 37464 3420
rect 37516 3408 37522 3460
rect 38013 3451 38071 3457
rect 38013 3417 38025 3451
rect 38059 3448 38071 3451
rect 38473 3451 38531 3457
rect 38473 3448 38485 3451
rect 38059 3420 38485 3448
rect 38059 3417 38071 3420
rect 38013 3411 38071 3417
rect 38473 3417 38485 3420
rect 38519 3417 38531 3451
rect 39224 3448 39252 3479
rect 39390 3476 39396 3528
rect 39448 3476 39454 3528
rect 41386 3516 41414 3624
rect 42058 3612 42064 3624
rect 42116 3612 42122 3664
rect 42996 3652 43024 3680
rect 43441 3655 43499 3661
rect 43441 3652 43453 3655
rect 42996 3624 43453 3652
rect 43441 3621 43453 3624
rect 43487 3621 43499 3655
rect 43441 3615 43499 3621
rect 43070 3544 43076 3596
rect 43128 3544 43134 3596
rect 43165 3587 43223 3593
rect 43165 3553 43177 3587
rect 43211 3584 43223 3587
rect 43548 3584 43576 3692
rect 45738 3680 45744 3692
rect 45796 3680 45802 3732
rect 46201 3723 46259 3729
rect 46201 3689 46213 3723
rect 46247 3720 46259 3723
rect 47854 3720 47860 3732
rect 46247 3692 47860 3720
rect 46247 3689 46259 3692
rect 46201 3683 46259 3689
rect 47854 3680 47860 3692
rect 47912 3680 47918 3732
rect 48317 3723 48375 3729
rect 48317 3689 48329 3723
rect 48363 3720 48375 3723
rect 48590 3720 48596 3732
rect 48363 3692 48596 3720
rect 48363 3689 48375 3692
rect 48317 3683 48375 3689
rect 48590 3680 48596 3692
rect 48648 3680 48654 3732
rect 49050 3680 49056 3732
rect 49108 3720 49114 3732
rect 49108 3692 49280 3720
rect 49108 3680 49114 3692
rect 45281 3655 45339 3661
rect 45281 3652 45293 3655
rect 44284 3624 45293 3652
rect 43211 3556 43576 3584
rect 43717 3587 43775 3593
rect 43211 3553 43223 3556
rect 43165 3547 43223 3553
rect 43717 3553 43729 3587
rect 43763 3584 43775 3587
rect 44174 3584 44180 3596
rect 43763 3556 44180 3584
rect 43763 3553 43775 3556
rect 43717 3547 43775 3553
rect 44174 3544 44180 3556
rect 44232 3544 44238 3596
rect 44284 3593 44312 3624
rect 45281 3621 45293 3624
rect 45327 3621 45339 3655
rect 45281 3615 45339 3621
rect 47397 3655 47455 3661
rect 47397 3621 47409 3655
rect 47443 3652 47455 3655
rect 47762 3652 47768 3664
rect 47443 3624 47768 3652
rect 47443 3621 47455 3624
rect 47397 3615 47455 3621
rect 47762 3612 47768 3624
rect 47820 3612 47826 3664
rect 49145 3655 49203 3661
rect 49145 3652 49157 3655
rect 48516 3624 49157 3652
rect 44269 3587 44327 3593
rect 44269 3553 44281 3587
rect 44315 3553 44327 3587
rect 44269 3547 44327 3553
rect 45002 3544 45008 3596
rect 45060 3544 45066 3596
rect 45094 3544 45100 3596
rect 45152 3584 45158 3596
rect 45370 3584 45376 3596
rect 45152 3556 45376 3584
rect 45152 3544 45158 3556
rect 45370 3544 45376 3556
rect 45428 3584 45434 3596
rect 45833 3587 45891 3593
rect 45833 3584 45845 3587
rect 45428 3556 45845 3584
rect 45428 3544 45434 3556
rect 45833 3553 45845 3556
rect 45879 3553 45891 3587
rect 45833 3547 45891 3553
rect 46842 3544 46848 3596
rect 46900 3544 46906 3596
rect 47121 3587 47179 3593
rect 47121 3553 47133 3587
rect 47167 3584 47179 3587
rect 47302 3584 47308 3596
rect 47167 3556 47308 3584
rect 47167 3553 47179 3556
rect 47121 3547 47179 3553
rect 47302 3544 47308 3556
rect 47360 3544 47366 3596
rect 48516 3593 48544 3624
rect 49145 3621 49157 3624
rect 49191 3621 49203 3655
rect 49145 3615 49203 3621
rect 48041 3587 48099 3593
rect 48041 3553 48053 3587
rect 48087 3584 48099 3587
rect 48501 3587 48559 3593
rect 48087 3556 48452 3584
rect 48087 3553 48099 3556
rect 48041 3547 48099 3553
rect 40144 3488 41414 3516
rect 40144 3448 40172 3488
rect 41966 3476 41972 3528
rect 42024 3476 42030 3528
rect 42153 3519 42211 3525
rect 42153 3485 42165 3519
rect 42199 3485 42211 3519
rect 42153 3479 42211 3485
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3516 42855 3519
rect 43625 3519 43683 3525
rect 43625 3516 43637 3519
rect 42843 3488 43637 3516
rect 42843 3485 42855 3488
rect 42797 3479 42855 3485
rect 43625 3485 43637 3488
rect 43671 3485 43683 3519
rect 43625 3479 43683 3485
rect 39224 3420 40172 3448
rect 40221 3451 40279 3457
rect 38473 3411 38531 3417
rect 40221 3417 40233 3451
rect 40267 3448 40279 3451
rect 41417 3451 41475 3457
rect 41417 3448 41429 3451
rect 40267 3420 41429 3448
rect 40267 3417 40279 3420
rect 40221 3411 40279 3417
rect 41417 3417 41429 3420
rect 41463 3417 41475 3451
rect 41417 3411 41475 3417
rect 41782 3408 41788 3460
rect 41840 3448 41846 3460
rect 42168 3448 42196 3479
rect 43898 3476 43904 3528
rect 43956 3476 43962 3528
rect 43990 3476 43996 3528
rect 44048 3516 44054 3528
rect 45020 3516 45048 3544
rect 44048 3488 45048 3516
rect 45189 3519 45247 3525
rect 44048 3476 44054 3488
rect 45189 3485 45201 3519
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45741 3519 45799 3525
rect 45741 3485 45753 3519
rect 45787 3516 45799 3519
rect 46198 3516 46204 3528
rect 45787 3488 46204 3516
rect 45787 3485 45799 3488
rect 45741 3479 45799 3485
rect 41840 3420 42196 3448
rect 41840 3408 41846 3420
rect 42886 3408 42892 3460
rect 42944 3408 42950 3460
rect 43257 3451 43315 3457
rect 43257 3417 43269 3451
rect 43303 3448 43315 3451
rect 43806 3448 43812 3460
rect 43303 3420 43812 3448
rect 43303 3417 43315 3420
rect 43257 3411 43315 3417
rect 43806 3408 43812 3420
rect 43864 3408 43870 3460
rect 45204 3448 45232 3479
rect 46198 3476 46204 3488
rect 46256 3476 46262 3528
rect 47026 3525 47032 3528
rect 47004 3519 47032 3525
rect 47004 3485 47016 3519
rect 47004 3479 47032 3485
rect 47026 3476 47032 3479
rect 47084 3476 47090 3528
rect 47857 3519 47915 3525
rect 47857 3485 47869 3519
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 43916 3420 45232 3448
rect 47872 3448 47900 3479
rect 48130 3476 48136 3528
rect 48188 3476 48194 3528
rect 48424 3516 48452 3556
rect 48501 3553 48513 3587
rect 48547 3553 48559 3587
rect 48501 3547 48559 3553
rect 48866 3544 48872 3596
rect 48924 3584 48930 3596
rect 49053 3587 49111 3593
rect 49053 3584 49065 3587
rect 48924 3556 49065 3584
rect 48924 3544 48930 3556
rect 49053 3553 49065 3556
rect 49099 3553 49111 3587
rect 49252 3584 49280 3692
rect 51350 3680 51356 3732
rect 51408 3680 51414 3732
rect 51629 3723 51687 3729
rect 51629 3689 51641 3723
rect 51675 3720 51687 3723
rect 51994 3720 52000 3732
rect 51675 3692 52000 3720
rect 51675 3689 51687 3692
rect 51629 3683 51687 3689
rect 51994 3680 52000 3692
rect 52052 3680 52058 3732
rect 53190 3680 53196 3732
rect 53248 3720 53254 3732
rect 53561 3723 53619 3729
rect 53561 3720 53573 3723
rect 53248 3692 53573 3720
rect 53248 3680 53254 3692
rect 53561 3689 53573 3692
rect 53607 3689 53619 3723
rect 53561 3683 53619 3689
rect 53926 3680 53932 3732
rect 53984 3720 53990 3732
rect 54297 3723 54355 3729
rect 54297 3720 54309 3723
rect 53984 3692 54309 3720
rect 53984 3680 53990 3692
rect 54297 3689 54309 3692
rect 54343 3689 54355 3723
rect 54297 3683 54355 3689
rect 55030 3680 55036 3732
rect 55088 3680 55094 3732
rect 55214 3680 55220 3732
rect 55272 3720 55278 3732
rect 55401 3723 55459 3729
rect 55401 3720 55413 3723
rect 55272 3692 55413 3720
rect 55272 3680 55278 3692
rect 55401 3689 55413 3692
rect 55447 3689 55459 3723
rect 55401 3683 55459 3689
rect 51368 3652 51396 3680
rect 51813 3655 51871 3661
rect 51813 3652 51825 3655
rect 51368 3624 51825 3652
rect 51813 3621 51825 3624
rect 51859 3621 51871 3655
rect 51813 3615 51871 3621
rect 53469 3655 53527 3661
rect 53469 3621 53481 3655
rect 53515 3621 53527 3655
rect 53469 3615 53527 3621
rect 49697 3587 49755 3593
rect 49697 3584 49709 3587
rect 49252 3556 49709 3584
rect 49053 3547 49111 3553
rect 49697 3553 49709 3556
rect 49743 3553 49755 3587
rect 49697 3547 49755 3553
rect 49878 3544 49884 3596
rect 49936 3544 49942 3596
rect 50338 3544 50344 3596
rect 50396 3584 50402 3596
rect 53484 3584 53512 3615
rect 54205 3587 54263 3593
rect 54205 3584 54217 3587
rect 50396 3556 52132 3584
rect 53484 3556 54217 3584
rect 50396 3544 50402 3556
rect 49896 3516 49924 3544
rect 48424 3488 49924 3516
rect 50706 3476 50712 3528
rect 50764 3476 50770 3528
rect 50985 3519 51043 3525
rect 50985 3485 50997 3519
rect 51031 3485 51043 3519
rect 50985 3479 51043 3485
rect 49418 3448 49424 3460
rect 47872 3420 49424 3448
rect 29788 3352 29960 3380
rect 30009 3383 30067 3389
rect 29788 3340 29794 3352
rect 30009 3349 30021 3383
rect 30055 3380 30067 3383
rect 30377 3383 30435 3389
rect 30377 3380 30389 3383
rect 30055 3352 30389 3380
rect 30055 3349 30067 3352
rect 30009 3343 30067 3349
rect 30377 3349 30389 3352
rect 30423 3349 30435 3383
rect 30377 3343 30435 3349
rect 31110 3340 31116 3392
rect 31168 3340 31174 3392
rect 31386 3340 31392 3392
rect 31444 3340 31450 3392
rect 32861 3383 32919 3389
rect 32861 3349 32873 3383
rect 32907 3380 32919 3383
rect 33502 3380 33508 3392
rect 32907 3352 33508 3380
rect 32907 3349 32919 3352
rect 32861 3343 32919 3349
rect 33502 3340 33508 3352
rect 33560 3340 33566 3392
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 37550 3380 37556 3392
rect 36044 3352 37556 3380
rect 36044 3340 36050 3352
rect 37550 3340 37556 3352
rect 37608 3340 37614 3392
rect 39577 3383 39635 3389
rect 39577 3349 39589 3383
rect 39623 3380 39635 3383
rect 39850 3380 39856 3392
rect 39623 3352 39856 3380
rect 39623 3349 39635 3352
rect 39577 3343 39635 3349
rect 39850 3340 39856 3352
rect 39908 3340 39914 3392
rect 40678 3340 40684 3392
rect 40736 3340 40742 3392
rect 43162 3340 43168 3392
rect 43220 3380 43226 3392
rect 43916 3380 43944 3420
rect 49418 3408 49424 3420
rect 49476 3408 49482 3460
rect 49513 3451 49571 3457
rect 49513 3417 49525 3451
rect 49559 3448 49571 3451
rect 50157 3451 50215 3457
rect 50157 3448 50169 3451
rect 49559 3420 50169 3448
rect 49559 3417 49571 3420
rect 49513 3411 49571 3417
rect 50157 3417 50169 3420
rect 50203 3417 50215 3451
rect 50157 3411 50215 3417
rect 50246 3408 50252 3460
rect 50304 3448 50310 3460
rect 51000 3448 51028 3479
rect 51902 3476 51908 3528
rect 51960 3476 51966 3528
rect 51994 3476 52000 3528
rect 52052 3476 52058 3528
rect 52104 3525 52132 3556
rect 54205 3553 54217 3556
rect 54251 3584 54263 3587
rect 55048 3584 55076 3680
rect 58526 3652 58532 3664
rect 56612 3624 58532 3652
rect 56612 3593 56640 3624
rect 58526 3612 58532 3624
rect 58584 3612 58590 3664
rect 54251 3556 55076 3584
rect 56597 3587 56655 3593
rect 54251 3553 54263 3556
rect 54205 3547 54263 3553
rect 56597 3553 56609 3587
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 57238 3544 57244 3596
rect 57296 3584 57302 3596
rect 57609 3587 57667 3593
rect 57609 3584 57621 3587
rect 57296 3556 57621 3584
rect 57296 3544 57302 3556
rect 57609 3553 57621 3556
rect 57655 3553 57667 3587
rect 57609 3547 57667 3553
rect 52089 3519 52147 3525
rect 52089 3485 52101 3519
rect 52135 3516 52147 3519
rect 52822 3516 52828 3528
rect 52135 3488 52828 3516
rect 52135 3485 52147 3488
rect 52089 3479 52147 3485
rect 52822 3476 52828 3488
rect 52880 3476 52886 3528
rect 54846 3476 54852 3528
rect 54904 3476 54910 3528
rect 55585 3519 55643 3525
rect 55585 3485 55597 3519
rect 55631 3516 55643 3519
rect 55631 3488 57008 3516
rect 55631 3485 55643 3488
rect 55585 3479 55643 3485
rect 50304 3420 51028 3448
rect 51920 3448 51948 3476
rect 52334 3451 52392 3457
rect 52334 3448 52346 3451
rect 51920 3420 52346 3448
rect 50304 3408 50310 3420
rect 52334 3417 52346 3420
rect 52380 3417 52392 3451
rect 54864 3448 54892 3476
rect 52334 3411 52392 3417
rect 54128 3420 54892 3448
rect 56980 3448 57008 3488
rect 57054 3476 57060 3528
rect 57112 3476 57118 3528
rect 57146 3476 57152 3528
rect 57204 3476 57210 3528
rect 57882 3448 57888 3460
rect 56980 3420 57888 3448
rect 54128 3392 54156 3420
rect 57882 3408 57888 3420
rect 57940 3408 57946 3460
rect 43220 3352 43944 3380
rect 44085 3383 44143 3389
rect 43220 3340 43226 3352
rect 44085 3349 44097 3383
rect 44131 3380 44143 3383
rect 44174 3380 44180 3392
rect 44131 3352 44180 3380
rect 44131 3349 44143 3352
rect 44085 3343 44143 3349
rect 44174 3340 44180 3352
rect 44232 3340 44238 3392
rect 44818 3340 44824 3392
rect 44876 3340 44882 3392
rect 45002 3340 45008 3392
rect 45060 3340 45066 3392
rect 45646 3340 45652 3392
rect 45704 3340 45710 3392
rect 46198 3340 46204 3392
rect 46256 3380 46262 3392
rect 47486 3380 47492 3392
rect 46256 3352 47492 3380
rect 46256 3340 46262 3352
rect 47486 3340 47492 3352
rect 47544 3340 47550 3392
rect 48406 3340 48412 3392
rect 48464 3380 48470 3392
rect 49605 3383 49663 3389
rect 49605 3380 49617 3383
rect 48464 3352 49617 3380
rect 48464 3340 48470 3352
rect 49605 3349 49617 3352
rect 49651 3349 49663 3383
rect 49605 3343 49663 3349
rect 49694 3340 49700 3392
rect 49752 3380 49758 3392
rect 51718 3380 51724 3392
rect 49752 3352 51724 3380
rect 49752 3340 49758 3352
rect 51718 3340 51724 3352
rect 51776 3340 51782 3392
rect 54110 3340 54116 3392
rect 54168 3340 54174 3392
rect 1104 3290 59040 3312
rect 1104 3238 15394 3290
rect 15446 3238 15458 3290
rect 15510 3238 15522 3290
rect 15574 3238 15586 3290
rect 15638 3238 15650 3290
rect 15702 3238 29838 3290
rect 29890 3238 29902 3290
rect 29954 3238 29966 3290
rect 30018 3238 30030 3290
rect 30082 3238 30094 3290
rect 30146 3238 44282 3290
rect 44334 3238 44346 3290
rect 44398 3238 44410 3290
rect 44462 3238 44474 3290
rect 44526 3238 44538 3290
rect 44590 3238 58726 3290
rect 58778 3238 58790 3290
rect 58842 3238 58854 3290
rect 58906 3238 58918 3290
rect 58970 3238 58982 3290
rect 59034 3238 59040 3290
rect 1104 3216 59040 3238
rect 1854 3136 1860 3188
rect 1912 3136 1918 3188
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2130 3176 2136 3188
rect 1995 3148 2136 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4120 3148 4476 3176
rect 4120 3136 4126 3148
rect 4240 3111 4298 3117
rect 1780 3080 4016 3108
rect 1780 3052 1808 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 1688 2972 1716 3003
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 3073 3043 3131 3049
rect 3073 3009 3085 3043
rect 3119 3040 3131 3043
rect 3234 3040 3240 3052
rect 3119 3012 3240 3040
rect 3119 3009 3131 3012
rect 3073 3003 3131 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3344 3049 3372 3080
rect 3988 3049 4016 3080
rect 4240 3077 4252 3111
rect 4286 3108 4298 3111
rect 4338 3108 4344 3120
rect 4286 3080 4344 3108
rect 4286 3077 4298 3080
rect 4240 3071 4298 3077
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4448 3108 4476 3148
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 5258 3176 5264 3188
rect 4672 3148 5264 3176
rect 4672 3136 4678 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5902 3176 5908 3188
rect 5399 3148 5908 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 6972 3148 7389 3176
rect 6972 3136 6978 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 7558 3136 7564 3188
rect 7616 3136 7622 3188
rect 7926 3136 7932 3188
rect 7984 3136 7990 3188
rect 9766 3176 9772 3188
rect 9232 3148 9772 3176
rect 4448 3080 6132 3108
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 3973 3003 4031 3009
rect 4080 3012 5457 3040
rect 2314 2972 2320 2984
rect 1688 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 3620 2972 3648 3003
rect 4080 2972 4108 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 3620 2944 4108 2972
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5040 2944 6009 2972
rect 5040 2932 5046 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 5534 2864 5540 2916
rect 5592 2864 5598 2916
rect 6104 2904 6132 3080
rect 6380 3049 6408 3136
rect 6733 3111 6791 3117
rect 6733 3077 6745 3111
rect 6779 3108 6791 3111
rect 7576 3108 7604 3136
rect 6779 3080 7604 3108
rect 9064 3111 9122 3117
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 9064 3077 9076 3111
rect 9110 3108 9122 3111
rect 9232 3108 9260 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 11330 3136 11336 3188
rect 11388 3136 11394 3188
rect 11514 3136 11520 3188
rect 11572 3136 11578 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11756 3148 11897 3176
rect 11756 3136 11762 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 11977 3179 12035 3185
rect 11977 3145 11989 3179
rect 12023 3176 12035 3179
rect 14550 3176 14556 3188
rect 12023 3148 14556 3176
rect 12023 3145 12035 3148
rect 11977 3139 12035 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 15896 3148 16405 3176
rect 15896 3136 15902 3148
rect 16393 3145 16405 3148
rect 16439 3145 16451 3179
rect 16393 3139 16451 3145
rect 17678 3136 17684 3188
rect 17736 3136 17742 3188
rect 17954 3136 17960 3188
rect 18012 3136 18018 3188
rect 18230 3136 18236 3188
rect 18288 3136 18294 3188
rect 18322 3136 18328 3188
rect 18380 3136 18386 3188
rect 18414 3136 18420 3188
rect 18472 3176 18478 3188
rect 18693 3179 18751 3185
rect 18693 3176 18705 3179
rect 18472 3148 18705 3176
rect 18472 3136 18478 3148
rect 18693 3145 18705 3148
rect 18739 3145 18751 3179
rect 18693 3139 18751 3145
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19889 3179 19947 3185
rect 19889 3176 19901 3179
rect 18840 3148 19901 3176
rect 18840 3136 18846 3148
rect 19889 3145 19901 3148
rect 19935 3145 19947 3179
rect 19889 3139 19947 3145
rect 20165 3179 20223 3185
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20806 3176 20812 3188
rect 20211 3148 20812 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 21542 3136 21548 3188
rect 21600 3136 21606 3188
rect 21818 3136 21824 3188
rect 21876 3176 21882 3188
rect 22925 3179 22983 3185
rect 21876 3148 22600 3176
rect 21876 3136 21882 3148
rect 9674 3108 9680 3120
rect 9110 3080 9260 3108
rect 9324 3080 9680 3108
rect 9110 3077 9122 3080
rect 9064 3071 9122 3077
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6512 3012 6837 3040
rect 6512 3000 6518 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 7282 3040 7288 3052
rect 7147 3012 7288 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 9324 3049 9352 3080
rect 9674 3068 9680 3080
rect 9732 3108 9738 3120
rect 10220 3111 10278 3117
rect 9732 3080 10180 3108
rect 9732 3068 9738 3080
rect 9968 3049 9996 3080
rect 9309 3043 9367 3049
rect 8260 3012 9260 3040
rect 8260 3000 8266 3012
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 7484 2972 7512 3000
rect 6696 2944 7512 2972
rect 9232 2972 9260 3012
rect 9309 3009 9321 3043
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 9416 2972 9444 3003
rect 9232 2944 9444 2972
rect 9600 2972 9628 3003
rect 10042 3000 10048 3052
rect 10100 3000 10106 3052
rect 10152 3040 10180 3080
rect 10220 3077 10232 3111
rect 10266 3108 10278 3111
rect 10888 3108 10916 3136
rect 13814 3108 13820 3120
rect 10266 3080 10916 3108
rect 11164 3080 13820 3108
rect 10266 3077 10278 3080
rect 10220 3071 10278 3077
rect 11164 3040 11192 3080
rect 13814 3068 13820 3080
rect 13872 3108 13878 3120
rect 17120 3111 17178 3117
rect 13872 3080 14228 3108
rect 13872 3068 13878 3080
rect 10152 3012 11192 3040
rect 11256 3012 12434 3040
rect 10060 2972 10088 3000
rect 11256 2984 11284 3012
rect 9600 2944 10088 2972
rect 6696 2932 6702 2944
rect 11238 2932 11244 2984
rect 11296 2932 11302 2984
rect 12066 2932 12072 2984
rect 12124 2932 12130 2984
rect 12406 2972 12434 3012
rect 12526 3000 12532 3052
rect 12584 3000 12590 3052
rect 13929 3043 13987 3049
rect 13929 3009 13941 3043
rect 13975 3040 13987 3043
rect 14090 3040 14096 3052
rect 13975 3012 14096 3040
rect 13975 3009 13987 3012
rect 13929 3003 13987 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14200 3049 14228 3080
rect 17120 3077 17132 3111
rect 17166 3108 17178 3111
rect 17696 3108 17724 3136
rect 17166 3080 17724 3108
rect 17972 3108 18000 3136
rect 19153 3111 19211 3117
rect 19153 3108 19165 3111
rect 17972 3080 19165 3108
rect 17166 3077 17178 3080
rect 17120 3071 17178 3077
rect 19153 3077 19165 3080
rect 19199 3077 19211 3111
rect 19153 3071 19211 3077
rect 21300 3111 21358 3117
rect 21300 3077 21312 3111
rect 21346 3108 21358 3111
rect 21560 3108 21588 3136
rect 21346 3080 21588 3108
rect 21346 3077 21358 3080
rect 21300 3071 21358 3077
rect 21726 3068 21732 3120
rect 21784 3108 21790 3120
rect 21784 3080 22140 3108
rect 21784 3068 21790 3080
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 14976 3012 15485 3040
rect 14976 3000 14982 3012
rect 15473 3009 15485 3012
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 18046 3000 18052 3052
rect 18104 3040 18110 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 18104 3012 20085 3040
rect 18104 3000 18110 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 21545 3043 21603 3049
rect 21545 3009 21557 3043
rect 21591 3040 21603 3043
rect 22002 3040 22008 3052
rect 21591 3012 22008 3040
rect 21591 3009 21603 3012
rect 21545 3003 21603 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 22112 3049 22140 3080
rect 22572 3049 22600 3148
rect 22925 3145 22937 3179
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3009 22155 3043
rect 22097 3003 22155 3009
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3009 22615 3043
rect 22557 3003 22615 3009
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 12710 2972 12716 2984
rect 12406 2944 12716 2972
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 14458 2932 14464 2984
rect 14516 2932 14522 2984
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15344 2944 15761 2972
rect 15344 2932 15350 2944
rect 15749 2941 15761 2944
rect 15795 2941 15807 2975
rect 15749 2935 15807 2941
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16264 2944 16865 2972
rect 16264 2932 16270 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 16853 2935 16911 2941
rect 18524 2944 18797 2972
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 6104 2876 7205 2904
rect 7193 2873 7205 2876
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 9692 2876 9996 2904
rect 3789 2839 3847 2845
rect 3789 2805 3801 2839
rect 3835 2836 3847 2839
rect 5552 2836 5580 2864
rect 3835 2808 5580 2836
rect 3835 2805 3847 2808
rect 3789 2799 3847 2805
rect 7742 2796 7748 2848
rect 7800 2796 7806 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9692 2836 9720 2876
rect 9088 2808 9720 2836
rect 9088 2796 9094 2808
rect 9766 2796 9772 2848
rect 9824 2796 9830 2848
rect 9968 2836 9996 2876
rect 10888 2876 13308 2904
rect 10888 2836 10916 2876
rect 9968 2808 10916 2836
rect 12342 2796 12348 2848
rect 12400 2796 12406 2848
rect 12802 2796 12808 2848
rect 12860 2796 12866 2848
rect 13280 2836 13308 2876
rect 14642 2836 14648 2848
rect 13280 2808 14648 2836
rect 14642 2796 14648 2808
rect 14700 2836 14706 2848
rect 15010 2836 15016 2848
rect 14700 2808 15016 2836
rect 14700 2796 14706 2808
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 18524 2836 18552 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 18874 2932 18880 2984
rect 18932 2932 18938 2984
rect 19705 2975 19763 2981
rect 19705 2941 19717 2975
rect 19751 2941 19763 2975
rect 21468 2972 21496 3000
rect 21913 2975 21971 2981
rect 21913 2972 21925 2975
rect 21468 2944 21925 2972
rect 19705 2935 19763 2941
rect 21913 2941 21925 2944
rect 21959 2972 21971 2975
rect 22664 2972 22692 3003
rect 21959 2944 22692 2972
rect 22940 2972 22968 3139
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 23477 3179 23535 3185
rect 23477 3176 23489 3179
rect 23072 3148 23489 3176
rect 23072 3136 23078 3148
rect 23477 3145 23489 3148
rect 23523 3145 23535 3179
rect 23477 3139 23535 3145
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 26789 3179 26847 3185
rect 26789 3145 26801 3179
rect 26835 3176 26847 3179
rect 27246 3176 27252 3188
rect 26835 3148 27252 3176
rect 26835 3145 26847 3148
rect 26789 3139 26847 3145
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 27522 3136 27528 3188
rect 27580 3136 27586 3188
rect 27617 3179 27675 3185
rect 27617 3145 27629 3179
rect 27663 3145 27675 3179
rect 27617 3139 27675 3145
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 23109 3043 23167 3049
rect 23109 3040 23121 3043
rect 23072 3012 23121 3040
rect 23072 3000 23078 3012
rect 23109 3009 23121 3012
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 23385 3043 23443 3049
rect 23385 3009 23397 3043
rect 23431 3040 23443 3043
rect 23750 3040 23756 3052
rect 23431 3012 23756 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24136 3040 24164 3136
rect 26234 3108 26240 3120
rect 25884 3080 26240 3108
rect 25884 3049 25912 3080
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 24136 3012 24225 3040
rect 24213 3009 24225 3012
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 25869 3043 25927 3049
rect 25869 3009 25881 3043
rect 25915 3009 25927 3043
rect 27540 3040 27568 3136
rect 27632 3108 27660 3139
rect 29086 3136 29092 3188
rect 29144 3176 29150 3188
rect 30834 3176 30840 3188
rect 29144 3148 30840 3176
rect 29144 3136 29150 3148
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 31754 3136 31760 3188
rect 31812 3176 31818 3188
rect 32125 3179 32183 3185
rect 32125 3176 32137 3179
rect 31812 3148 32137 3176
rect 31812 3136 31818 3148
rect 32125 3145 32137 3148
rect 32171 3145 32183 3179
rect 32125 3139 32183 3145
rect 33502 3136 33508 3188
rect 33560 3176 33566 3188
rect 33560 3148 33640 3176
rect 33560 3136 33566 3148
rect 27954 3111 28012 3117
rect 27954 3108 27966 3111
rect 27632 3080 27966 3108
rect 27954 3077 27966 3080
rect 28000 3077 28012 3111
rect 27954 3071 28012 3077
rect 28258 3068 28264 3120
rect 28316 3108 28322 3120
rect 28316 3080 31892 3108
rect 28316 3068 28322 3080
rect 25869 3003 25927 3009
rect 25976 3012 27568 3040
rect 23293 2975 23351 2981
rect 22940 2944 23244 2972
rect 21959 2941 21971 2944
rect 21913 2935 21971 2941
rect 18598 2864 18604 2916
rect 18656 2904 18662 2916
rect 19720 2904 19748 2935
rect 18656 2876 19748 2904
rect 18656 2864 18662 2876
rect 20254 2864 20260 2916
rect 20312 2864 20318 2916
rect 21542 2864 21548 2916
rect 21600 2904 21606 2916
rect 23216 2904 23244 2944
rect 23293 2941 23305 2975
rect 23339 2972 23351 2975
rect 23474 2972 23480 2984
rect 23339 2944 23480 2972
rect 23339 2941 23351 2944
rect 23293 2935 23351 2941
rect 23474 2932 23480 2944
rect 23532 2932 23538 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23624 2944 24041 2972
rect 23624 2932 23630 2944
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 24118 2932 24124 2984
rect 24176 2972 24182 2984
rect 24673 2975 24731 2981
rect 24673 2972 24685 2975
rect 24176 2944 24685 2972
rect 24176 2932 24182 2944
rect 24673 2941 24685 2944
rect 24719 2941 24731 2975
rect 24673 2935 24731 2941
rect 25685 2975 25743 2981
rect 25685 2941 25697 2975
rect 25731 2972 25743 2975
rect 25774 2972 25780 2984
rect 25731 2944 25780 2972
rect 25731 2941 25743 2944
rect 25685 2935 25743 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 25976 2904 26004 3012
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27672 3012 27721 3040
rect 27672 3000 27678 3012
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 28994 3040 29000 3052
rect 27709 3003 27767 3009
rect 27816 3012 29000 3040
rect 26237 2975 26295 2981
rect 26237 2941 26249 2975
rect 26283 2972 26295 2975
rect 26602 2972 26608 2984
rect 26283 2944 26608 2972
rect 26283 2941 26295 2944
rect 26237 2935 26295 2941
rect 26602 2932 26608 2944
rect 26660 2932 26666 2984
rect 27065 2975 27123 2981
rect 27065 2941 27077 2975
rect 27111 2972 27123 2975
rect 27816 2972 27844 3012
rect 28994 3000 29000 3012
rect 29052 3000 29058 3052
rect 29178 3000 29184 3052
rect 29236 3000 29242 3052
rect 31662 3000 31668 3052
rect 31720 3000 31726 3052
rect 27111 2944 27844 2972
rect 27111 2941 27123 2944
rect 27065 2935 27123 2941
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 29144 2944 29653 2972
rect 29144 2932 29150 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 30190 2932 30196 2984
rect 30248 2972 30254 2984
rect 31864 2981 31892 3080
rect 33249 3043 33307 3049
rect 33249 3009 33261 3043
rect 33295 3040 33307 3043
rect 33295 3012 33456 3040
rect 33295 3009 33307 3012
rect 33249 3003 33307 3009
rect 30745 2975 30803 2981
rect 30745 2972 30757 2975
rect 30248 2944 30757 2972
rect 30248 2932 30254 2944
rect 30745 2941 30757 2944
rect 30791 2941 30803 2975
rect 30745 2935 30803 2941
rect 31849 2975 31907 2981
rect 31849 2941 31861 2975
rect 31895 2972 31907 2975
rect 33428 2972 33456 3012
rect 33502 3000 33508 3052
rect 33560 3000 33566 3052
rect 33612 3040 33640 3148
rect 34606 3136 34612 3188
rect 34664 3176 34670 3188
rect 35069 3179 35127 3185
rect 35069 3176 35081 3179
rect 34664 3148 35081 3176
rect 34664 3136 34670 3148
rect 35069 3145 35081 3148
rect 35115 3145 35127 3179
rect 35069 3139 35127 3145
rect 36265 3179 36323 3185
rect 36265 3145 36277 3179
rect 36311 3176 36323 3179
rect 36354 3176 36360 3188
rect 36311 3148 36360 3176
rect 36311 3145 36323 3148
rect 36265 3139 36323 3145
rect 36354 3136 36360 3148
rect 36412 3136 36418 3188
rect 38470 3136 38476 3188
rect 38528 3136 38534 3188
rect 40678 3136 40684 3188
rect 40736 3136 40742 3188
rect 41598 3136 41604 3188
rect 41656 3136 41662 3188
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 42429 3179 42487 3185
rect 42429 3176 42441 3179
rect 41932 3148 42441 3176
rect 41932 3136 41938 3148
rect 42429 3145 42441 3148
rect 42475 3145 42487 3179
rect 42429 3139 42487 3145
rect 43070 3136 43076 3188
rect 43128 3176 43134 3188
rect 43165 3179 43223 3185
rect 43165 3176 43177 3179
rect 43128 3148 43177 3176
rect 43128 3136 43134 3148
rect 43165 3145 43177 3148
rect 43211 3145 43223 3179
rect 43165 3139 43223 3145
rect 43530 3136 43536 3188
rect 43588 3136 43594 3188
rect 44361 3179 44419 3185
rect 44361 3145 44373 3179
rect 44407 3176 44419 3179
rect 44726 3176 44732 3188
rect 44407 3148 44732 3176
rect 44407 3145 44419 3148
rect 44361 3139 44419 3145
rect 44726 3136 44732 3148
rect 44784 3136 44790 3188
rect 45002 3136 45008 3188
rect 45060 3136 45066 3188
rect 47210 3136 47216 3188
rect 47268 3176 47274 3188
rect 47581 3179 47639 3185
rect 47581 3176 47593 3179
rect 47268 3148 47593 3176
rect 47268 3136 47274 3148
rect 47581 3145 47593 3148
rect 47627 3145 47639 3179
rect 47581 3139 47639 3145
rect 48314 3136 48320 3188
rect 48372 3136 48378 3188
rect 49418 3136 49424 3188
rect 49476 3176 49482 3188
rect 50157 3179 50215 3185
rect 50157 3176 50169 3179
rect 49476 3148 50169 3176
rect 49476 3136 49482 3148
rect 50157 3145 50169 3148
rect 50203 3176 50215 3179
rect 50706 3176 50712 3188
rect 50203 3148 50712 3176
rect 50203 3145 50215 3148
rect 50157 3139 50215 3145
rect 50706 3136 50712 3148
rect 50764 3136 50770 3188
rect 54018 3136 54024 3188
rect 54076 3136 54082 3188
rect 54110 3136 54116 3188
rect 54168 3136 54174 3188
rect 55950 3136 55956 3188
rect 56008 3136 56014 3188
rect 57514 3176 57520 3188
rect 57256 3148 57520 3176
rect 34977 3111 35035 3117
rect 34977 3077 34989 3111
rect 35023 3108 35035 3111
rect 38488 3108 38516 3136
rect 35023 3080 36492 3108
rect 35023 3077 35035 3080
rect 34977 3071 35035 3077
rect 34149 3043 34207 3049
rect 34149 3040 34161 3043
rect 33612 3012 34161 3040
rect 34149 3009 34161 3012
rect 34195 3009 34207 3043
rect 34149 3003 34207 3009
rect 35253 3043 35311 3049
rect 35253 3009 35265 3043
rect 35299 3040 35311 3043
rect 35434 3040 35440 3052
rect 35299 3012 35440 3040
rect 35299 3009 35311 3012
rect 35253 3003 35311 3009
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35529 3043 35587 3049
rect 35529 3009 35541 3043
rect 35575 3040 35587 3043
rect 35618 3040 35624 3052
rect 35575 3012 35624 3040
rect 35575 3009 35587 3012
rect 35529 3003 35587 3009
rect 35618 3000 35624 3012
rect 35676 3000 35682 3052
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3040 35955 3043
rect 35986 3040 35992 3052
rect 35943 3012 35992 3040
rect 35943 3009 35955 3012
rect 35897 3003 35955 3009
rect 35986 3000 35992 3012
rect 36044 3000 36050 3052
rect 36081 3043 36139 3049
rect 36081 3009 36093 3043
rect 36127 3040 36139 3043
rect 36354 3040 36360 3052
rect 36127 3012 36360 3040
rect 36127 3009 36139 3012
rect 36081 3003 36139 3009
rect 36354 3000 36360 3012
rect 36412 3000 36418 3052
rect 36464 3049 36492 3080
rect 36740 3080 38516 3108
rect 39384 3111 39442 3117
rect 36740 3049 36768 3080
rect 39384 3077 39396 3111
rect 39430 3108 39442 3111
rect 40696 3108 40724 3136
rect 39430 3080 40724 3108
rect 39430 3077 39442 3080
rect 39384 3071 39442 3077
rect 36449 3043 36507 3049
rect 36449 3009 36461 3043
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 36725 3043 36783 3049
rect 36725 3009 36737 3043
rect 36771 3009 36783 3043
rect 36725 3003 36783 3009
rect 33597 2975 33655 2981
rect 33597 2972 33609 2975
rect 31895 2944 32536 2972
rect 33428 2944 33609 2972
rect 31895 2941 31907 2944
rect 31849 2935 31907 2941
rect 21600 2876 22600 2904
rect 23216 2876 26004 2904
rect 31389 2907 31447 2913
rect 21600 2864 21606 2876
rect 20272 2836 20300 2864
rect 18524 2808 20300 2836
rect 22278 2796 22284 2848
rect 22336 2796 22342 2848
rect 22370 2796 22376 2848
rect 22428 2796 22434 2848
rect 22572 2836 22600 2876
rect 31389 2873 31401 2907
rect 31435 2904 31447 2907
rect 32030 2904 32036 2916
rect 31435 2876 32036 2904
rect 31435 2873 31447 2876
rect 31389 2867 31447 2873
rect 32030 2864 32036 2876
rect 32088 2864 32094 2916
rect 23109 2839 23167 2845
rect 23109 2836 23121 2839
rect 22572 2808 23121 2836
rect 23109 2805 23121 2808
rect 23155 2805 23167 2839
rect 23109 2799 23167 2805
rect 26053 2839 26111 2845
rect 26053 2805 26065 2839
rect 26099 2836 26111 2839
rect 27706 2836 27712 2848
rect 26099 2808 27712 2836
rect 26099 2805 26111 2808
rect 26053 2799 26111 2805
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 31481 2839 31539 2845
rect 31481 2805 31493 2839
rect 31527 2836 31539 2839
rect 31754 2836 31760 2848
rect 31527 2808 31760 2836
rect 31527 2805 31539 2808
rect 31481 2799 31539 2805
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 32508 2836 32536 2944
rect 33597 2941 33609 2944
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 34333 2975 34391 2981
rect 34333 2941 34345 2975
rect 34379 2941 34391 2975
rect 34333 2935 34391 2941
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 34348 2904 34376 2935
rect 35342 2932 35348 2984
rect 35400 2932 35406 2984
rect 35710 2932 35716 2984
rect 35768 2972 35774 2984
rect 36740 2972 36768 3003
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 37001 3043 37059 3049
rect 37001 3009 37013 3043
rect 37047 3040 37059 3043
rect 37461 3043 37519 3049
rect 37461 3040 37473 3043
rect 37047 3012 37473 3040
rect 37047 3009 37059 3012
rect 37001 3003 37059 3009
rect 37461 3009 37473 3012
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 38654 3000 38660 3052
rect 38712 3040 38718 3052
rect 39117 3043 39175 3049
rect 39117 3040 39129 3043
rect 38712 3012 39129 3040
rect 38712 3000 38718 3012
rect 39117 3009 39129 3012
rect 39163 3009 39175 3043
rect 41616 3040 41644 3136
rect 41969 3043 42027 3049
rect 41969 3040 41981 3043
rect 41616 3012 41981 3040
rect 39117 3003 39175 3009
rect 41969 3009 41981 3012
rect 42015 3009 42027 3043
rect 41969 3003 42027 3009
rect 43346 3000 43352 3052
rect 43404 3000 43410 3052
rect 43548 3040 43576 3136
rect 44818 3117 44824 3120
rect 43625 3111 43683 3117
rect 43625 3077 43637 3111
rect 43671 3108 43683 3111
rect 43671 3080 44772 3108
rect 43671 3077 43683 3080
rect 43625 3071 43683 3077
rect 43901 3043 43959 3049
rect 43901 3040 43913 3043
rect 43548 3012 43913 3040
rect 43901 3009 43913 3012
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 43990 3000 43996 3052
rect 44048 3000 44054 3052
rect 44082 3000 44088 3052
rect 44140 3000 44146 3052
rect 44177 3043 44235 3049
rect 44177 3009 44189 3043
rect 44223 3040 44235 3043
rect 44450 3040 44456 3052
rect 44223 3012 44456 3040
rect 44223 3009 44235 3012
rect 44177 3003 44235 3009
rect 44450 3000 44456 3012
rect 44508 3000 44514 3052
rect 44545 3043 44603 3049
rect 44545 3009 44557 3043
rect 44591 3040 44603 3043
rect 44634 3040 44640 3052
rect 44591 3012 44640 3040
rect 44591 3009 44603 3012
rect 44545 3003 44603 3009
rect 44634 3000 44640 3012
rect 44692 3000 44698 3052
rect 44744 3040 44772 3080
rect 44812 3071 44824 3117
rect 44876 3108 44882 3120
rect 44876 3080 44912 3108
rect 44818 3068 44824 3071
rect 44876 3068 44882 3080
rect 45020 3040 45048 3136
rect 45094 3068 45100 3120
rect 45152 3108 45158 3120
rect 45152 3080 48268 3108
rect 45152 3068 45158 3080
rect 44744 3012 45048 3040
rect 45278 3000 45284 3052
rect 45336 3040 45342 3052
rect 46017 3043 46075 3049
rect 46017 3040 46029 3043
rect 45336 3012 46029 3040
rect 45336 3000 45342 3012
rect 46017 3009 46029 3012
rect 46063 3009 46075 3043
rect 46017 3003 46075 3009
rect 46934 3000 46940 3052
rect 46992 3000 46998 3052
rect 48240 3049 48268 3080
rect 48225 3043 48283 3049
rect 48225 3009 48237 3043
rect 48271 3009 48283 3043
rect 48332 3040 48360 3136
rect 50338 3108 50344 3120
rect 48792 3080 50344 3108
rect 48792 3049 48820 3080
rect 50338 3068 50344 3080
rect 50396 3068 50402 3120
rect 53000 3111 53058 3117
rect 53000 3077 53012 3111
rect 53046 3108 53058 3111
rect 53558 3108 53564 3120
rect 53046 3080 53564 3108
rect 53046 3077 53058 3080
rect 53000 3071 53058 3077
rect 53558 3068 53564 3080
rect 53616 3068 53622 3120
rect 48501 3043 48559 3049
rect 48501 3040 48513 3043
rect 48332 3012 48513 3040
rect 48225 3003 48283 3009
rect 48501 3009 48513 3012
rect 48547 3009 48559 3043
rect 48501 3003 48559 3009
rect 48777 3043 48835 3049
rect 48777 3009 48789 3043
rect 48823 3009 48835 3043
rect 48777 3003 48835 3009
rect 48866 3000 48872 3052
rect 48924 3040 48930 3052
rect 49044 3043 49102 3049
rect 49044 3040 49056 3043
rect 48924 3012 49056 3040
rect 48924 3000 48930 3012
rect 49044 3009 49056 3012
rect 49090 3009 49102 3043
rect 49044 3003 49102 3009
rect 49602 3000 49608 3052
rect 49660 3040 49666 3052
rect 50433 3043 50491 3049
rect 50433 3040 50445 3043
rect 49660 3012 50445 3040
rect 49660 3000 49666 3012
rect 50433 3009 50445 3012
rect 50479 3009 50491 3043
rect 50433 3003 50491 3009
rect 50617 3043 50675 3049
rect 50617 3009 50629 3043
rect 50663 3040 50675 3043
rect 52089 3043 52147 3049
rect 50663 3012 52040 3040
rect 50663 3009 50675 3012
rect 50617 3003 50675 3009
rect 35768 2944 36768 2972
rect 35768 2932 35774 2944
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37700 2944 37933 2972
rect 37700 2932 37706 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 38470 2932 38476 2984
rect 38528 2972 38534 2984
rect 38528 2944 38654 2972
rect 38528 2932 38534 2944
rect 33560 2876 34376 2904
rect 33560 2864 33566 2876
rect 34146 2836 34152 2848
rect 32508 2808 34152 2836
rect 34146 2796 34152 2808
rect 34204 2796 34210 2848
rect 35529 2839 35587 2845
rect 35529 2805 35541 2839
rect 35575 2836 35587 2839
rect 35986 2836 35992 2848
rect 35575 2808 35992 2836
rect 35575 2805 35587 2808
rect 35529 2799 35587 2805
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 37458 2836 37464 2848
rect 36412 2808 37464 2836
rect 36412 2796 36418 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 38626 2836 38654 2944
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 40957 2975 41015 2981
rect 40957 2972 40969 2975
rect 40736 2944 40969 2972
rect 40736 2932 40742 2944
rect 40957 2941 40969 2944
rect 41003 2941 41015 2975
rect 42981 2975 43039 2981
rect 42981 2972 42993 2975
rect 40957 2935 41015 2941
rect 41248 2944 42993 2972
rect 40126 2864 40132 2916
rect 40184 2904 40190 2916
rect 41248 2904 41276 2944
rect 42981 2941 42993 2944
rect 43027 2941 43039 2975
rect 42981 2935 43039 2941
rect 43533 2975 43591 2981
rect 43533 2941 43545 2975
rect 43579 2972 43591 2975
rect 44008 2972 44036 3000
rect 43579 2944 44036 2972
rect 43579 2941 43591 2944
rect 43533 2935 43591 2941
rect 45830 2932 45836 2984
rect 45888 2972 45894 2984
rect 46477 2975 46535 2981
rect 46477 2972 46489 2975
rect 45888 2944 46489 2972
rect 45888 2932 45894 2944
rect 46477 2941 46489 2944
rect 46523 2941 46535 2975
rect 46952 2972 46980 3000
rect 48038 2972 48044 2984
rect 46952 2944 48044 2972
rect 46477 2935 46535 2941
rect 48038 2932 48044 2944
rect 48096 2972 48102 2984
rect 48685 2975 48743 2981
rect 48685 2972 48697 2975
rect 48096 2944 48697 2972
rect 48096 2932 48102 2944
rect 48685 2941 48697 2944
rect 48731 2941 48743 2975
rect 48685 2935 48743 2941
rect 50706 2932 50712 2984
rect 50764 2972 50770 2984
rect 50893 2975 50951 2981
rect 50893 2972 50905 2975
rect 50764 2944 50905 2972
rect 50764 2932 50770 2944
rect 50893 2941 50905 2944
rect 50939 2941 50951 2975
rect 52012 2972 52040 3012
rect 52089 3009 52101 3043
rect 52135 3040 52147 3043
rect 52181 3043 52239 3049
rect 52181 3040 52193 3043
rect 52135 3012 52193 3040
rect 52135 3009 52147 3012
rect 52089 3003 52147 3009
rect 52181 3009 52193 3012
rect 52227 3009 52239 3043
rect 52181 3003 52239 3009
rect 52362 3000 52368 3052
rect 52420 3000 52426 3052
rect 52733 3043 52791 3049
rect 52733 3009 52745 3043
rect 52779 3040 52791 3043
rect 52822 3040 52828 3052
rect 52779 3012 52828 3040
rect 52779 3009 52791 3012
rect 52733 3003 52791 3009
rect 52822 3000 52828 3012
rect 52880 3000 52886 3052
rect 54036 3040 54064 3136
rect 57088 3111 57146 3117
rect 57088 3077 57100 3111
rect 57134 3108 57146 3111
rect 57256 3108 57284 3148
rect 57514 3136 57520 3148
rect 57572 3136 57578 3188
rect 57698 3136 57704 3188
rect 57756 3136 57762 3188
rect 57882 3136 57888 3188
rect 57940 3136 57946 3188
rect 57716 3108 57744 3136
rect 57134 3080 57284 3108
rect 57348 3080 57744 3108
rect 57134 3077 57146 3080
rect 57088 3071 57146 3077
rect 54205 3043 54263 3049
rect 54205 3040 54217 3043
rect 54036 3012 54217 3040
rect 54205 3009 54217 3012
rect 54251 3009 54263 3043
rect 54205 3003 54263 3009
rect 54478 3000 54484 3052
rect 54536 3040 54542 3052
rect 57348 3049 57376 3080
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 54536 3012 55873 3040
rect 54536 3000 54542 3012
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 57333 3043 57391 3049
rect 55861 3003 55919 3009
rect 55968 3012 57284 3040
rect 52546 2972 52552 2984
rect 52012 2944 52552 2972
rect 50893 2935 50951 2941
rect 52546 2932 52552 2944
rect 52604 2932 52610 2984
rect 53926 2932 53932 2984
rect 53984 2972 53990 2984
rect 54665 2975 54723 2981
rect 54665 2972 54677 2975
rect 53984 2944 54677 2972
rect 53984 2932 53990 2944
rect 54665 2941 54677 2944
rect 54711 2941 54723 2975
rect 54665 2935 54723 2941
rect 55030 2932 55036 2984
rect 55088 2972 55094 2984
rect 55968 2972 55996 3012
rect 55088 2944 55996 2972
rect 57256 2972 57284 3012
rect 57333 3009 57345 3043
rect 57379 3009 57391 3043
rect 57333 3003 57391 3009
rect 57698 3000 57704 3052
rect 57756 3000 57762 3052
rect 58437 2975 58495 2981
rect 58437 2972 58449 2975
rect 57256 2944 58449 2972
rect 55088 2932 55094 2944
rect 58437 2941 58449 2944
rect 58483 2941 58495 2975
rect 58437 2935 58495 2941
rect 40184 2876 41276 2904
rect 40184 2864 40190 2876
rect 42242 2864 42248 2916
rect 42300 2904 42306 2916
rect 52178 2904 52184 2916
rect 42300 2876 42840 2904
rect 42300 2864 42306 2876
rect 40402 2836 40408 2848
rect 38626 2808 40408 2836
rect 40402 2796 40408 2808
rect 40460 2796 40466 2848
rect 40497 2839 40555 2845
rect 40497 2805 40509 2839
rect 40543 2836 40555 2839
rect 41966 2836 41972 2848
rect 40543 2808 41972 2836
rect 40543 2805 40555 2808
rect 40497 2799 40555 2805
rect 41966 2796 41972 2808
rect 42024 2796 42030 2848
rect 42812 2836 42840 2876
rect 49712 2876 52184 2904
rect 43349 2839 43407 2845
rect 43349 2836 43361 2839
rect 42812 2808 43361 2836
rect 43349 2805 43361 2808
rect 43395 2805 43407 2839
rect 43349 2799 43407 2805
rect 43714 2796 43720 2848
rect 43772 2796 43778 2848
rect 43990 2796 43996 2848
rect 44048 2836 44054 2848
rect 45554 2836 45560 2848
rect 44048 2808 45560 2836
rect 44048 2796 44054 2808
rect 45554 2796 45560 2808
rect 45612 2796 45618 2848
rect 45925 2839 45983 2845
rect 45925 2805 45937 2839
rect 45971 2836 45983 2839
rect 47026 2836 47032 2848
rect 45971 2808 47032 2836
rect 45971 2805 45983 2808
rect 45925 2799 45983 2805
rect 47026 2796 47032 2808
rect 47084 2796 47090 2848
rect 48314 2796 48320 2848
rect 48372 2796 48378 2848
rect 48406 2796 48412 2848
rect 48464 2836 48470 2848
rect 49712 2836 49740 2876
rect 52178 2864 52184 2876
rect 52236 2864 52242 2916
rect 57974 2904 57980 2916
rect 53668 2876 55812 2904
rect 48464 2808 49740 2836
rect 48464 2796 48470 2808
rect 50246 2796 50252 2848
rect 50304 2796 50310 2848
rect 53374 2796 53380 2848
rect 53432 2836 53438 2848
rect 53668 2836 53696 2876
rect 53432 2808 53696 2836
rect 53432 2796 53438 2808
rect 55398 2796 55404 2848
rect 55456 2836 55462 2848
rect 55677 2839 55735 2845
rect 55677 2836 55689 2839
rect 55456 2808 55689 2836
rect 55456 2796 55462 2808
rect 55677 2805 55689 2808
rect 55723 2805 55735 2839
rect 55784 2836 55812 2876
rect 57348 2876 57980 2904
rect 57348 2836 57376 2876
rect 57974 2864 57980 2876
rect 58032 2864 58038 2916
rect 55784 2808 57376 2836
rect 55677 2799 55735 2805
rect 57422 2796 57428 2848
rect 57480 2836 57486 2848
rect 57517 2839 57575 2845
rect 57517 2836 57529 2839
rect 57480 2808 57529 2836
rect 57480 2796 57486 2808
rect 57517 2805 57529 2808
rect 57563 2805 57575 2839
rect 57517 2799 57575 2805
rect 1104 2746 58880 2768
rect 1104 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 22616 2746
rect 22668 2694 22680 2746
rect 22732 2694 22744 2746
rect 22796 2694 22808 2746
rect 22860 2694 22872 2746
rect 22924 2694 37060 2746
rect 37112 2694 37124 2746
rect 37176 2694 37188 2746
rect 37240 2694 37252 2746
rect 37304 2694 37316 2746
rect 37368 2694 51504 2746
rect 51556 2694 51568 2746
rect 51620 2694 51632 2746
rect 51684 2694 51696 2746
rect 51748 2694 51760 2746
rect 51812 2694 58880 2746
rect 1104 2672 58880 2694
rect 1946 2592 1952 2644
rect 2004 2592 2010 2644
rect 7742 2632 7748 2644
rect 6886 2604 7748 2632
rect 6886 2496 6914 2604
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9858 2632 9864 2644
rect 9815 2604 9864 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 12434 2592 12440 2644
rect 12492 2592 12498 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 14056 2604 14105 2632
rect 14056 2592 14062 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 14274 2592 14280 2644
rect 14332 2592 14338 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17586 2632 17592 2644
rect 17543 2604 17592 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 19429 2635 19487 2641
rect 19429 2601 19441 2635
rect 19475 2632 19487 2635
rect 21542 2632 21548 2644
rect 19475 2604 21548 2632
rect 19475 2601 19487 2604
rect 19429 2595 19487 2601
rect 21542 2592 21548 2604
rect 21600 2592 21606 2644
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21692 2604 21833 2632
rect 21692 2592 21698 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 21821 2595 21879 2601
rect 22370 2592 22376 2644
rect 22428 2592 22434 2644
rect 23474 2592 23480 2644
rect 23532 2592 23538 2644
rect 23750 2592 23756 2644
rect 23808 2632 23814 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23808 2604 24041 2632
rect 23808 2592 23814 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 25317 2635 25375 2641
rect 25317 2601 25329 2635
rect 25363 2632 25375 2635
rect 26418 2632 26424 2644
rect 25363 2604 26424 2632
rect 25363 2601 25375 2604
rect 25317 2595 25375 2601
rect 26418 2592 26424 2604
rect 26476 2592 26482 2644
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 26936 2604 26985 2632
rect 26936 2592 26942 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 26973 2595 27031 2601
rect 27430 2592 27436 2644
rect 27488 2592 27494 2644
rect 28626 2592 28632 2644
rect 28684 2592 28690 2644
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29549 2635 29607 2641
rect 29549 2632 29561 2635
rect 29052 2604 29561 2632
rect 29052 2592 29058 2604
rect 29549 2601 29561 2604
rect 29595 2601 29607 2635
rect 29549 2595 29607 2601
rect 31386 2592 31392 2644
rect 31444 2592 31450 2644
rect 32309 2635 32367 2641
rect 32309 2601 32321 2635
rect 32355 2632 32367 2635
rect 33778 2632 33784 2644
rect 32355 2604 33784 2632
rect 32355 2601 32367 2604
rect 32309 2595 32367 2601
rect 33778 2592 33784 2604
rect 33836 2592 33842 2644
rect 35710 2632 35716 2644
rect 34348 2604 35716 2632
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 8036 2564 8064 2592
rect 12452 2564 12480 2592
rect 7331 2536 8064 2564
rect 11532 2536 12480 2564
rect 13817 2567 13875 2573
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 3528 2468 6914 2496
rect 3528 2437 3556 2468
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7616 2468 7849 2496
rect 7616 2456 7622 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 10008 2468 10333 2496
rect 10008 2456 10014 2468
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4890 2428 4896 2440
rect 4111 2400 4896 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7006 2428 7012 2440
rect 6779 2400 7012 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 1670 2320 1676 2372
rect 1728 2320 1734 2372
rect 2038 2320 2044 2372
rect 2096 2360 2102 2372
rect 2317 2363 2375 2369
rect 2317 2360 2329 2363
rect 2096 2332 2329 2360
rect 2096 2320 2102 2332
rect 2317 2329 2329 2332
rect 2363 2329 2375 2363
rect 2317 2323 2375 2329
rect 5258 2320 5264 2372
rect 5316 2320 5322 2372
rect 6380 2360 6408 2391
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7374 2388 7380 2440
rect 7432 2388 7438 2440
rect 9214 2388 9220 2440
rect 9272 2388 9278 2440
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 11532 2437 11560 2536
rect 13817 2533 13829 2567
rect 13863 2564 13875 2567
rect 14292 2564 14320 2592
rect 13863 2536 14320 2564
rect 20165 2567 20223 2573
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 20714 2564 20720 2576
rect 20211 2536 20720 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12216 2468 12541 2496
rect 12216 2456 12222 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 14182 2496 14188 2508
rect 12529 2459 12587 2465
rect 13648 2468 14188 2496
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9824 2400 9873 2428
rect 9824 2388 9830 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12342 2428 12348 2440
rect 12299 2400 12348 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 13648 2437 13676 2468
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14550 2456 14556 2508
rect 14608 2456 14614 2508
rect 14642 2456 14648 2508
rect 14700 2456 14706 2508
rect 15838 2456 15844 2508
rect 15896 2456 15902 2508
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 17920 2468 18061 2496
rect 17920 2456 17926 2468
rect 18049 2465 18061 2468
rect 18095 2465 18107 2499
rect 22388 2496 22416 2592
rect 23492 2564 23520 2592
rect 24397 2567 24455 2573
rect 24397 2564 24409 2567
rect 23492 2536 24409 2564
rect 24397 2533 24409 2536
rect 24443 2533 24455 2567
rect 28644 2564 28672 2592
rect 31404 2564 31432 2592
rect 24397 2527 24455 2533
rect 27264 2536 28672 2564
rect 29104 2536 31432 2564
rect 18049 2459 18107 2465
rect 21652 2468 22416 2496
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13964 2400 14473 2428
rect 13964 2388 13970 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17276 2400 17601 2428
rect 17276 2388 17282 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19426 2428 19432 2440
rect 19291 2400 19432 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 20254 2428 20260 2440
rect 19659 2400 20260 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 21652 2437 21680 2468
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 21637 2431 21695 2437
rect 21637 2397 21649 2431
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22152 2400 22385 2428
rect 22152 2388 22158 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 8386 2360 8392 2372
rect 6380 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 14366 2320 14372 2372
rect 14424 2320 14430 2372
rect 20714 2320 20720 2372
rect 20772 2320 20778 2372
rect 22278 2320 22284 2372
rect 22336 2360 22342 2372
rect 22572 2360 22600 2391
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 23256 2400 24225 2428
rect 23256 2388 23262 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 25222 2428 25228 2440
rect 24811 2400 25228 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 26786 2388 26792 2440
rect 26844 2388 26850 2440
rect 27264 2437 27292 2536
rect 27614 2456 27620 2508
rect 27672 2496 27678 2508
rect 27985 2499 28043 2505
rect 27985 2496 27997 2499
rect 27672 2468 27997 2496
rect 27672 2456 27678 2468
rect 27985 2465 27997 2468
rect 28031 2465 28043 2499
rect 27985 2459 28043 2465
rect 27157 2431 27215 2437
rect 27157 2397 27169 2431
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2397 27307 2431
rect 27249 2391 27307 2397
rect 22336 2332 22600 2360
rect 22336 2320 22342 2332
rect 25774 2320 25780 2372
rect 25832 2320 25838 2372
rect 26973 2363 27031 2369
rect 26973 2329 26985 2363
rect 27019 2329 27031 2363
rect 27172 2360 27200 2391
rect 27706 2388 27712 2440
rect 27764 2388 27770 2440
rect 29104 2437 29132 2536
rect 29730 2456 29736 2508
rect 29788 2496 29794 2508
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29788 2468 30021 2496
rect 29788 2456 29794 2468
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 30098 2456 30104 2508
rect 30156 2456 30162 2508
rect 31110 2456 31116 2508
rect 31168 2456 31174 2508
rect 34348 2505 34376 2604
rect 35710 2592 35716 2604
rect 35768 2592 35774 2644
rect 35986 2592 35992 2644
rect 36044 2632 36050 2644
rect 36909 2635 36967 2641
rect 36909 2632 36921 2635
rect 36044 2604 36921 2632
rect 36044 2592 36050 2604
rect 36909 2601 36921 2604
rect 36955 2601 36967 2635
rect 36909 2595 36967 2601
rect 36998 2592 37004 2644
rect 37056 2632 37062 2644
rect 38749 2635 38807 2641
rect 38749 2632 38761 2635
rect 37056 2604 38761 2632
rect 37056 2592 37062 2604
rect 38749 2601 38761 2604
rect 38795 2601 38807 2635
rect 38749 2595 38807 2601
rect 38948 2604 42104 2632
rect 35434 2524 35440 2576
rect 35492 2564 35498 2576
rect 38948 2564 38976 2604
rect 42076 2573 42104 2604
rect 43346 2592 43352 2644
rect 43404 2592 43410 2644
rect 44450 2592 44456 2644
rect 44508 2632 44514 2644
rect 44545 2635 44603 2641
rect 44545 2632 44557 2635
rect 44508 2604 44557 2632
rect 44508 2592 44514 2604
rect 44545 2601 44557 2604
rect 44591 2601 44603 2635
rect 44545 2595 44603 2601
rect 45646 2592 45652 2644
rect 45704 2632 45710 2644
rect 46477 2635 46535 2641
rect 46477 2632 46489 2635
rect 45704 2604 46489 2632
rect 45704 2592 45710 2604
rect 46477 2601 46489 2604
rect 46523 2601 46535 2635
rect 46477 2595 46535 2601
rect 49786 2592 49792 2644
rect 49844 2592 49850 2644
rect 51166 2592 51172 2644
rect 51224 2632 51230 2644
rect 51629 2635 51687 2641
rect 51629 2632 51641 2635
rect 51224 2604 51641 2632
rect 51224 2592 51230 2604
rect 51629 2601 51641 2604
rect 51675 2601 51687 2635
rect 51629 2595 51687 2601
rect 51902 2592 51908 2644
rect 51960 2632 51966 2644
rect 52365 2635 52423 2641
rect 52365 2632 52377 2635
rect 51960 2604 52377 2632
rect 51960 2592 51966 2604
rect 52365 2601 52377 2604
rect 52411 2601 52423 2635
rect 52365 2595 52423 2601
rect 54573 2635 54631 2641
rect 54573 2601 54585 2635
rect 54619 2632 54631 2635
rect 55306 2632 55312 2644
rect 54619 2604 55312 2632
rect 54619 2601 54631 2604
rect 54573 2595 54631 2601
rect 55306 2592 55312 2604
rect 55364 2592 55370 2644
rect 55766 2632 55772 2644
rect 55600 2604 55772 2632
rect 35492 2536 38976 2564
rect 39485 2567 39543 2573
rect 35492 2524 35498 2536
rect 39485 2533 39497 2567
rect 39531 2533 39543 2567
rect 39485 2527 39543 2533
rect 42061 2567 42119 2573
rect 42061 2533 42073 2567
rect 42107 2533 42119 2567
rect 43364 2564 43392 2592
rect 44637 2567 44695 2573
rect 44637 2564 44649 2567
rect 43364 2536 44649 2564
rect 42061 2527 42119 2533
rect 44637 2533 44649 2536
rect 44683 2533 44695 2567
rect 54297 2567 54355 2573
rect 54297 2564 54309 2567
rect 44637 2527 44695 2533
rect 45664 2536 54309 2564
rect 34333 2499 34391 2505
rect 34333 2465 34345 2499
rect 34379 2465 34391 2499
rect 34333 2459 34391 2465
rect 34422 2456 34428 2508
rect 34480 2496 34486 2508
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 34480 2468 35173 2496
rect 34480 2456 34486 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 35161 2459 35219 2465
rect 35710 2456 35716 2508
rect 35768 2496 35774 2508
rect 39500 2496 39528 2527
rect 35768 2468 37596 2496
rect 35768 2456 35774 2468
rect 29089 2431 29147 2437
rect 29089 2397 29101 2431
rect 29135 2397 29147 2431
rect 29089 2391 29147 2397
rect 29270 2388 29276 2440
rect 29328 2428 29334 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29328 2400 29929 2428
rect 29328 2388 29334 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 31128 2428 31156 2456
rect 29917 2391 29975 2397
rect 30024 2400 31156 2428
rect 30024 2360 30052 2400
rect 31754 2388 31760 2440
rect 31812 2388 31818 2440
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 32088 2400 32137 2428
rect 32088 2388 32094 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 33226 2428 33232 2440
rect 32125 2391 32183 2397
rect 32232 2400 33232 2428
rect 27172 2332 30052 2360
rect 26973 2323 27031 2329
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 7650 2292 7656 2304
rect 6595 2264 7656 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 14384 2292 14412 2320
rect 11747 2264 14412 2292
rect 26988 2292 27016 2323
rect 30742 2320 30748 2372
rect 30800 2320 30806 2372
rect 28810 2292 28816 2304
rect 26988 2264 28816 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 28810 2252 28816 2264
rect 28868 2252 28874 2304
rect 29273 2295 29331 2301
rect 29273 2261 29285 2295
rect 29319 2292 29331 2295
rect 32232 2292 32260 2400
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 33873 2431 33931 2437
rect 33873 2397 33885 2431
rect 33919 2428 33931 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33919 2400 33977 2428
rect 33919 2397 33931 2400
rect 33873 2391 33931 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 34149 2431 34207 2437
rect 34149 2428 34161 2431
rect 34112 2400 34161 2428
rect 34112 2388 34118 2400
rect 34149 2397 34161 2400
rect 34195 2397 34207 2431
rect 34149 2391 34207 2397
rect 34698 2388 34704 2440
rect 34756 2388 34762 2440
rect 35250 2388 35256 2440
rect 35308 2428 35314 2440
rect 36725 2431 36783 2437
rect 36725 2428 36737 2431
rect 35308 2400 36737 2428
rect 35308 2388 35314 2400
rect 36725 2397 36737 2400
rect 36771 2397 36783 2431
rect 36725 2391 36783 2397
rect 37090 2388 37096 2440
rect 37148 2388 37154 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 37568 2428 37596 2468
rect 38304 2468 39528 2496
rect 40313 2499 40371 2505
rect 38197 2431 38255 2437
rect 38197 2428 38209 2431
rect 37568 2400 38209 2428
rect 38197 2397 38209 2400
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 32677 2363 32735 2369
rect 32677 2360 32689 2363
rect 32456 2332 32689 2360
rect 32456 2320 32462 2332
rect 32677 2329 32689 2332
rect 32723 2329 32735 2363
rect 32677 2323 32735 2329
rect 35618 2320 35624 2372
rect 35676 2360 35682 2372
rect 38304 2360 38332 2468
rect 40313 2465 40325 2499
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 39301 2431 39359 2437
rect 39301 2428 39313 2431
rect 35676 2332 38332 2360
rect 38488 2400 39313 2428
rect 35676 2320 35682 2332
rect 29319 2264 32260 2292
rect 29319 2261 29331 2264
rect 29273 2255 29331 2261
rect 35894 2252 35900 2304
rect 35952 2292 35958 2304
rect 36173 2295 36231 2301
rect 36173 2292 36185 2295
rect 35952 2264 36185 2292
rect 35952 2252 35958 2264
rect 36173 2261 36185 2264
rect 36219 2261 36231 2295
rect 36173 2255 36231 2261
rect 36814 2252 36820 2304
rect 36872 2292 36878 2304
rect 38488 2292 38516 2400
rect 39301 2397 39313 2400
rect 39347 2397 39359 2431
rect 39301 2391 39359 2397
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 39850 2388 39856 2440
rect 39908 2388 39914 2440
rect 39114 2320 39120 2372
rect 39172 2360 39178 2372
rect 40328 2360 40356 2459
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 41380 2468 44864 2496
rect 41380 2456 41386 2468
rect 40402 2388 40408 2440
rect 40460 2428 40466 2440
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 40460 2400 41889 2428
rect 40460 2388 40466 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 42242 2388 42248 2440
rect 42300 2388 42306 2440
rect 43714 2388 43720 2440
rect 43772 2388 43778 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 39172 2332 40356 2360
rect 39172 2320 39178 2332
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41325 2363 41383 2369
rect 41325 2360 41337 2363
rect 40644 2332 41337 2360
rect 40644 2320 40650 2332
rect 41325 2329 41337 2332
rect 41371 2329 41383 2363
rect 41325 2323 41383 2329
rect 42518 2320 42524 2372
rect 42576 2360 42582 2372
rect 42797 2363 42855 2369
rect 42797 2360 42809 2363
rect 42576 2332 42809 2360
rect 42576 2320 42582 2332
rect 42797 2329 42809 2332
rect 42843 2329 42855 2363
rect 42797 2323 42855 2329
rect 43438 2320 43444 2372
rect 43496 2360 43502 2372
rect 43916 2360 43944 2391
rect 44266 2388 44272 2440
rect 44324 2388 44330 2440
rect 44836 2437 44864 2468
rect 45554 2456 45560 2508
rect 45612 2456 45618 2508
rect 44821 2431 44879 2437
rect 44821 2397 44833 2431
rect 44867 2397 44879 2431
rect 44821 2391 44879 2397
rect 45005 2431 45063 2437
rect 45005 2397 45017 2431
rect 45051 2397 45063 2431
rect 45005 2391 45063 2397
rect 43496 2332 43944 2360
rect 44284 2360 44312 2388
rect 45020 2360 45048 2391
rect 44284 2332 45048 2360
rect 43496 2320 43502 2332
rect 36872 2264 38516 2292
rect 36872 2252 36878 2264
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 45664 2292 45692 2536
rect 54297 2533 54309 2536
rect 54343 2533 54355 2567
rect 54297 2527 54355 2533
rect 54496 2536 55536 2564
rect 47026 2456 47032 2508
rect 47084 2456 47090 2508
rect 49234 2456 49240 2508
rect 49292 2496 49298 2508
rect 50617 2499 50675 2505
rect 50617 2496 50629 2499
rect 49292 2468 50629 2496
rect 49292 2456 49298 2468
rect 50617 2465 50629 2468
rect 50663 2465 50675 2499
rect 50617 2459 50675 2465
rect 51994 2456 52000 2508
rect 52052 2456 52058 2508
rect 52454 2456 52460 2508
rect 52512 2496 52518 2508
rect 53193 2499 53251 2505
rect 53193 2496 53205 2499
rect 52512 2468 53205 2496
rect 52512 2456 52518 2468
rect 53193 2465 53205 2468
rect 53239 2465 53251 2499
rect 53193 2459 53251 2465
rect 53742 2456 53748 2508
rect 53800 2456 53806 2508
rect 48314 2388 48320 2440
rect 48372 2428 48378 2440
rect 48777 2431 48835 2437
rect 48777 2428 48789 2431
rect 48372 2400 48789 2428
rect 48372 2388 48378 2400
rect 48777 2397 48789 2400
rect 48823 2397 48835 2431
rect 48777 2391 48835 2397
rect 49053 2431 49111 2437
rect 49053 2397 49065 2431
rect 49099 2397 49111 2431
rect 49053 2391 49111 2397
rect 47302 2320 47308 2372
rect 47360 2360 47366 2372
rect 47765 2363 47823 2369
rect 47765 2360 47777 2363
rect 47360 2332 47777 2360
rect 47360 2320 47366 2332
rect 47765 2329 47777 2332
rect 47811 2329 47823 2363
rect 47765 2323 47823 2329
rect 43864 2264 45692 2292
rect 43864 2252 43870 2264
rect 46750 2252 46756 2304
rect 46808 2292 46814 2304
rect 49068 2292 49096 2391
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 49973 2431 50031 2437
rect 49973 2428 49985 2431
rect 49752 2400 49985 2428
rect 49752 2388 49758 2400
rect 49973 2397 49985 2400
rect 50019 2397 50031 2431
rect 49973 2391 50031 2397
rect 50246 2388 50252 2440
rect 50304 2388 50310 2440
rect 52012 2428 52040 2456
rect 50816 2400 52040 2428
rect 46808 2264 49096 2292
rect 49697 2295 49755 2301
rect 46808 2252 46814 2264
rect 49697 2261 49709 2295
rect 49743 2292 49755 2295
rect 50816 2292 50844 2400
rect 52178 2388 52184 2440
rect 52236 2388 52242 2440
rect 52549 2431 52607 2437
rect 52549 2397 52561 2431
rect 52595 2397 52607 2431
rect 52549 2391 52607 2397
rect 51350 2320 51356 2372
rect 51408 2360 51414 2372
rect 52564 2360 52592 2391
rect 52730 2388 52736 2440
rect 52788 2388 52794 2440
rect 51408 2332 52592 2360
rect 53760 2360 53788 2456
rect 54496 2437 54524 2536
rect 54941 2499 54999 2505
rect 54941 2465 54953 2499
rect 54987 2496 54999 2499
rect 55398 2496 55404 2508
rect 54987 2468 55404 2496
rect 54987 2465 54999 2468
rect 54941 2459 54999 2465
rect 55398 2456 55404 2468
rect 55456 2456 55462 2508
rect 54481 2431 54539 2437
rect 54481 2397 54493 2431
rect 54527 2397 54539 2431
rect 54481 2391 54539 2397
rect 54849 2431 54907 2437
rect 54849 2397 54861 2431
rect 54895 2397 54907 2431
rect 54849 2391 54907 2397
rect 54864 2360 54892 2391
rect 53760 2332 54892 2360
rect 55508 2360 55536 2536
rect 55600 2437 55628 2604
rect 55766 2592 55772 2604
rect 55824 2592 55830 2644
rect 57146 2592 57152 2644
rect 57204 2592 57210 2644
rect 57698 2592 57704 2644
rect 57756 2632 57762 2644
rect 57885 2635 57943 2641
rect 57885 2632 57897 2635
rect 57756 2604 57897 2632
rect 57756 2592 57762 2604
rect 57885 2601 57897 2604
rect 57931 2601 57943 2635
rect 57885 2595 57943 2601
rect 55766 2456 55772 2508
rect 55824 2496 55830 2508
rect 56137 2499 56195 2505
rect 56137 2496 56149 2499
rect 55824 2468 56149 2496
rect 55824 2456 55830 2468
rect 56137 2465 56149 2468
rect 56183 2465 56195 2499
rect 57606 2496 57612 2508
rect 56137 2459 56195 2465
rect 57348 2468 57612 2496
rect 55585 2431 55643 2437
rect 55585 2397 55597 2431
rect 55631 2397 55643 2431
rect 55585 2391 55643 2397
rect 55674 2388 55680 2440
rect 55732 2388 55738 2440
rect 57348 2437 57376 2468
rect 57606 2456 57612 2468
rect 57664 2456 57670 2508
rect 57974 2456 57980 2508
rect 58032 2496 58038 2508
rect 58437 2499 58495 2505
rect 58437 2496 58449 2499
rect 58032 2468 58449 2496
rect 58032 2456 58038 2468
rect 58437 2465 58449 2468
rect 58483 2465 58495 2499
rect 58437 2459 58495 2465
rect 57333 2431 57391 2437
rect 57333 2397 57345 2431
rect 57379 2397 57391 2431
rect 57333 2391 57391 2397
rect 57514 2388 57520 2440
rect 57572 2388 57578 2440
rect 58342 2360 58348 2372
rect 55508 2332 58348 2360
rect 51408 2320 51414 2332
rect 58342 2320 58348 2332
rect 58400 2320 58406 2372
rect 49743 2264 50844 2292
rect 49743 2261 49755 2264
rect 49697 2255 49755 2261
rect 50982 2252 50988 2304
rect 51040 2292 51046 2304
rect 55401 2295 55459 2301
rect 55401 2292 55413 2295
rect 51040 2264 55413 2292
rect 51040 2252 51046 2264
rect 55401 2261 55413 2264
rect 55447 2261 55459 2295
rect 55401 2255 55459 2261
rect 1104 2202 59040 2224
rect 1104 2150 15394 2202
rect 15446 2150 15458 2202
rect 15510 2150 15522 2202
rect 15574 2150 15586 2202
rect 15638 2150 15650 2202
rect 15702 2150 29838 2202
rect 29890 2150 29902 2202
rect 29954 2150 29966 2202
rect 30018 2150 30030 2202
rect 30082 2150 30094 2202
rect 30146 2150 44282 2202
rect 44334 2150 44346 2202
rect 44398 2150 44410 2202
rect 44462 2150 44474 2202
rect 44526 2150 44538 2202
rect 44590 2150 58726 2202
rect 58778 2150 58790 2202
rect 58842 2150 58854 2202
rect 58906 2150 58918 2202
rect 58970 2150 58982 2202
rect 59034 2150 59040 2202
rect 1104 2128 59040 2150
rect 34606 2048 34612 2100
rect 34664 2088 34670 2100
rect 39666 2088 39672 2100
rect 34664 2060 39672 2088
rect 34664 2048 34670 2060
rect 39666 2048 39672 2060
rect 39724 2048 39730 2100
rect 33042 1368 33048 1420
rect 33100 1408 33106 1420
rect 37090 1408 37096 1420
rect 33100 1380 37096 1408
rect 33100 1368 33106 1380
rect 37090 1368 37096 1380
rect 37148 1368 37154 1420
<< via1 >>
rect 15394 21734 15446 21786
rect 15458 21734 15510 21786
rect 15522 21734 15574 21786
rect 15586 21734 15638 21786
rect 15650 21734 15702 21786
rect 29838 21734 29890 21786
rect 29902 21734 29954 21786
rect 29966 21734 30018 21786
rect 30030 21734 30082 21786
rect 30094 21734 30146 21786
rect 44282 21734 44334 21786
rect 44346 21734 44398 21786
rect 44410 21734 44462 21786
rect 44474 21734 44526 21786
rect 44538 21734 44590 21786
rect 58726 21734 58778 21786
rect 58790 21734 58842 21786
rect 58854 21734 58906 21786
rect 58918 21734 58970 21786
rect 58982 21734 59034 21786
rect 38384 21496 38436 21548
rect 5632 21471 5684 21480
rect 5632 21437 5641 21471
rect 5641 21437 5675 21471
rect 5675 21437 5684 21471
rect 5632 21428 5684 21437
rect 9496 21471 9548 21480
rect 9496 21437 9505 21471
rect 9505 21437 9539 21471
rect 9539 21437 9548 21471
rect 9496 21428 9548 21437
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 13452 21428 13504 21480
rect 15200 21428 15252 21480
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 28356 21428 28408 21480
rect 30748 21471 30800 21480
rect 30748 21437 30757 21471
rect 30757 21437 30791 21471
rect 30791 21437 30800 21471
rect 30748 21428 30800 21437
rect 31576 21428 31628 21480
rect 32956 21428 33008 21480
rect 33416 21471 33468 21480
rect 33416 21437 33425 21471
rect 33425 21437 33459 21471
rect 33459 21437 33468 21471
rect 33416 21428 33468 21437
rect 38660 21471 38712 21480
rect 38660 21437 38669 21471
rect 38669 21437 38703 21471
rect 38703 21437 38712 21471
rect 38660 21428 38712 21437
rect 39856 21428 39908 21480
rect 43260 21471 43312 21480
rect 43260 21437 43269 21471
rect 43269 21437 43303 21471
rect 43303 21437 43312 21471
rect 43260 21428 43312 21437
rect 43996 21471 44048 21480
rect 43996 21437 44005 21471
rect 44005 21437 44039 21471
rect 44039 21437 44048 21471
rect 43996 21428 44048 21437
rect 44088 21428 44140 21480
rect 46112 21471 46164 21480
rect 46112 21437 46121 21471
rect 46121 21437 46155 21471
rect 46155 21437 46164 21471
rect 46112 21428 46164 21437
rect 48228 21471 48280 21480
rect 48228 21437 48237 21471
rect 48237 21437 48271 21471
rect 48271 21437 48280 21471
rect 48228 21428 48280 21437
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 53380 21471 53432 21480
rect 53380 21437 53389 21471
rect 53389 21437 53423 21471
rect 53423 21437 53432 21471
rect 53380 21428 53432 21437
rect 56600 21471 56652 21480
rect 56600 21437 56609 21471
rect 56609 21437 56643 21471
rect 56643 21437 56652 21471
rect 56600 21428 56652 21437
rect 31668 21360 31720 21412
rect 36912 21360 36964 21412
rect 4988 21335 5040 21344
rect 4988 21301 4997 21335
rect 4997 21301 5031 21335
rect 5031 21301 5040 21335
rect 4988 21292 5040 21301
rect 5172 21292 5224 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 11612 21292 11664 21344
rect 14832 21335 14884 21344
rect 14832 21301 14841 21335
rect 14841 21301 14875 21335
rect 14875 21301 14884 21335
rect 14832 21292 14884 21301
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 22376 21292 22428 21344
rect 25596 21292 25648 21344
rect 27252 21335 27304 21344
rect 27252 21301 27261 21335
rect 27261 21301 27295 21335
rect 27295 21301 27304 21335
rect 27252 21292 27304 21301
rect 28080 21335 28132 21344
rect 28080 21301 28089 21335
rect 28089 21301 28123 21335
rect 28123 21301 28132 21335
rect 28080 21292 28132 21301
rect 31300 21292 31352 21344
rect 31392 21335 31444 21344
rect 31392 21301 31401 21335
rect 31401 21301 31435 21335
rect 31435 21301 31444 21335
rect 31392 21292 31444 21301
rect 32956 21292 33008 21344
rect 33968 21335 34020 21344
rect 33968 21301 33977 21335
rect 33977 21301 34011 21335
rect 34011 21301 34020 21335
rect 33968 21292 34020 21301
rect 34520 21292 34572 21344
rect 36728 21292 36780 21344
rect 37648 21360 37700 21412
rect 46940 21360 46992 21412
rect 52000 21403 52052 21412
rect 52000 21369 52009 21403
rect 52009 21369 52043 21403
rect 52043 21369 52052 21403
rect 52000 21360 52052 21369
rect 38016 21335 38068 21344
rect 38016 21301 38025 21335
rect 38025 21301 38059 21335
rect 38059 21301 38068 21335
rect 38016 21292 38068 21301
rect 39212 21292 39264 21344
rect 40040 21292 40092 21344
rect 42708 21335 42760 21344
rect 42708 21301 42717 21335
rect 42717 21301 42751 21335
rect 42751 21301 42760 21335
rect 42708 21292 42760 21301
rect 43444 21335 43496 21344
rect 43444 21301 43453 21335
rect 43453 21301 43487 21335
rect 43487 21301 43496 21335
rect 43444 21292 43496 21301
rect 44824 21335 44876 21344
rect 44824 21301 44833 21335
rect 44833 21301 44867 21335
rect 44867 21301 44876 21335
rect 44824 21292 44876 21301
rect 45836 21335 45888 21344
rect 45836 21301 45845 21335
rect 45845 21301 45879 21335
rect 45879 21301 45888 21335
rect 45836 21292 45888 21301
rect 46480 21292 46532 21344
rect 46756 21335 46808 21344
rect 46756 21301 46765 21335
rect 46765 21301 46799 21335
rect 46799 21301 46808 21335
rect 46756 21292 46808 21301
rect 47584 21335 47636 21344
rect 47584 21301 47593 21335
rect 47593 21301 47627 21335
rect 47627 21301 47636 21335
rect 47584 21292 47636 21301
rect 48504 21335 48556 21344
rect 48504 21301 48513 21335
rect 48513 21301 48547 21335
rect 48547 21301 48556 21335
rect 48504 21292 48556 21301
rect 52828 21335 52880 21344
rect 52828 21301 52837 21335
rect 52837 21301 52871 21335
rect 52871 21301 52880 21335
rect 52828 21292 52880 21301
rect 54484 21292 54536 21344
rect 55956 21335 56008 21344
rect 55956 21301 55965 21335
rect 55965 21301 55999 21335
rect 55999 21301 56008 21335
rect 55956 21292 56008 21301
rect 56048 21335 56100 21344
rect 56048 21301 56057 21335
rect 56057 21301 56091 21335
rect 56091 21301 56100 21335
rect 56048 21292 56100 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 22616 21190 22668 21242
rect 22680 21190 22732 21242
rect 22744 21190 22796 21242
rect 22808 21190 22860 21242
rect 22872 21190 22924 21242
rect 37060 21190 37112 21242
rect 37124 21190 37176 21242
rect 37188 21190 37240 21242
rect 37252 21190 37304 21242
rect 37316 21190 37368 21242
rect 51504 21190 51556 21242
rect 51568 21190 51620 21242
rect 51632 21190 51684 21242
rect 51696 21190 51748 21242
rect 51760 21190 51812 21242
rect 5632 21088 5684 21140
rect 5172 20995 5224 21004
rect 5172 20961 5181 20995
rect 5181 20961 5215 20995
rect 5215 20961 5224 20995
rect 5172 20952 5224 20961
rect 5632 20884 5684 20936
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 8944 21088 8996 21140
rect 10784 21020 10836 21072
rect 13452 21088 13504 21140
rect 19156 21088 19208 21140
rect 8668 20952 8720 21004
rect 9404 20952 9456 21004
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 10876 20884 10928 20936
rect 12532 20884 12584 20936
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 13176 20884 13228 20936
rect 4160 20748 4212 20800
rect 7748 20791 7800 20800
rect 7748 20757 7757 20791
rect 7757 20757 7791 20791
rect 7791 20757 7800 20791
rect 7748 20748 7800 20757
rect 14832 20952 14884 21004
rect 22376 21020 22428 21072
rect 15752 20952 15804 21004
rect 24584 20952 24636 21004
rect 27804 21088 27856 21140
rect 28080 21088 28132 21140
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22100 20884 22152 20893
rect 22468 20884 22520 20936
rect 25228 20927 25280 20936
rect 25228 20893 25237 20927
rect 25237 20893 25271 20927
rect 25271 20893 25280 20927
rect 25228 20884 25280 20893
rect 25872 20927 25924 20936
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 31300 20952 31352 21004
rect 36728 21020 36780 21072
rect 28632 20927 28684 20936
rect 28632 20893 28641 20927
rect 28641 20893 28675 20927
rect 28675 20893 28684 20927
rect 28632 20884 28684 20893
rect 31852 20927 31904 20936
rect 31852 20893 31861 20927
rect 31861 20893 31895 20927
rect 31895 20893 31904 20927
rect 31852 20884 31904 20893
rect 25044 20816 25096 20868
rect 9036 20748 9088 20800
rect 9772 20791 9824 20800
rect 9772 20757 9781 20791
rect 9781 20757 9815 20791
rect 9815 20757 9824 20791
rect 9772 20748 9824 20757
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 14832 20791 14884 20800
rect 14832 20757 14841 20791
rect 14841 20757 14875 20791
rect 14875 20757 14884 20791
rect 14832 20748 14884 20757
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 18236 20791 18288 20800
rect 18236 20757 18245 20791
rect 18245 20757 18279 20791
rect 18279 20757 18288 20791
rect 18236 20748 18288 20757
rect 18696 20748 18748 20800
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 21548 20791 21600 20800
rect 21548 20757 21557 20791
rect 21557 20757 21591 20791
rect 21591 20757 21600 20791
rect 21548 20748 21600 20757
rect 23664 20748 23716 20800
rect 24676 20748 24728 20800
rect 27896 20816 27948 20868
rect 31484 20816 31536 20868
rect 34520 20884 34572 20936
rect 35256 20927 35308 20936
rect 35256 20893 35265 20927
rect 35265 20893 35299 20927
rect 35299 20893 35308 20927
rect 35256 20884 35308 20893
rect 37004 20952 37056 21004
rect 38016 21088 38068 21140
rect 39856 21131 39908 21140
rect 39856 21097 39865 21131
rect 39865 21097 39899 21131
rect 39899 21097 39908 21131
rect 39856 21088 39908 21097
rect 43444 21088 43496 21140
rect 46112 21088 46164 21140
rect 39212 20995 39264 21004
rect 39212 20961 39221 20995
rect 39221 20961 39255 20995
rect 39255 20961 39264 20995
rect 39212 20952 39264 20961
rect 41880 20927 41932 20936
rect 41880 20893 41889 20927
rect 41889 20893 41923 20927
rect 41923 20893 41932 20927
rect 41880 20884 41932 20893
rect 42432 20884 42484 20936
rect 44088 20952 44140 21004
rect 44180 20884 44232 20936
rect 47584 21088 47636 21140
rect 49148 21088 49200 21140
rect 52000 21088 52052 21140
rect 52828 21088 52880 21140
rect 56600 21088 56652 21140
rect 46480 20995 46532 21004
rect 46480 20961 46489 20995
rect 46489 20961 46523 20995
rect 46523 20961 46532 20995
rect 46480 20952 46532 20961
rect 46940 20995 46992 21004
rect 46940 20961 46949 20995
rect 46949 20961 46983 20995
rect 46983 20961 46992 20995
rect 46940 20952 46992 20961
rect 48780 20995 48832 21004
rect 48780 20961 48789 20995
rect 48789 20961 48823 20995
rect 48823 20961 48832 20995
rect 48780 20952 48832 20961
rect 53840 20952 53892 21004
rect 54668 20952 54720 21004
rect 33508 20816 33560 20868
rect 34612 20816 34664 20868
rect 28080 20791 28132 20800
rect 28080 20757 28089 20791
rect 28089 20757 28123 20791
rect 28123 20757 28132 20791
rect 28080 20748 28132 20757
rect 29000 20791 29052 20800
rect 29000 20757 29009 20791
rect 29009 20757 29043 20791
rect 29043 20757 29052 20791
rect 29000 20748 29052 20757
rect 29644 20791 29696 20800
rect 29644 20757 29653 20791
rect 29653 20757 29687 20791
rect 29687 20757 29696 20791
rect 29644 20748 29696 20757
rect 30840 20791 30892 20800
rect 30840 20757 30849 20791
rect 30849 20757 30883 20791
rect 30883 20757 30892 20791
rect 30840 20748 30892 20757
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 32128 20791 32180 20800
rect 32128 20757 32137 20791
rect 32137 20757 32171 20791
rect 32171 20757 32180 20791
rect 32128 20748 32180 20757
rect 33416 20748 33468 20800
rect 33784 20748 33836 20800
rect 34704 20791 34756 20800
rect 34704 20757 34713 20791
rect 34713 20757 34747 20791
rect 34747 20757 34756 20791
rect 34704 20748 34756 20757
rect 35992 20748 36044 20800
rect 37556 20748 37608 20800
rect 39948 20816 40000 20868
rect 47768 20884 47820 20936
rect 49424 20884 49476 20936
rect 51264 20884 51316 20936
rect 53472 20884 53524 20936
rect 38108 20791 38160 20800
rect 38108 20757 38117 20791
rect 38117 20757 38151 20791
rect 38151 20757 38160 20791
rect 38108 20748 38160 20757
rect 38476 20791 38528 20800
rect 38476 20757 38485 20791
rect 38485 20757 38519 20791
rect 38519 20757 38528 20791
rect 38476 20748 38528 20757
rect 38568 20791 38620 20800
rect 38568 20757 38577 20791
rect 38577 20757 38611 20791
rect 38611 20757 38620 20791
rect 38568 20748 38620 20757
rect 39028 20791 39080 20800
rect 39028 20757 39037 20791
rect 39037 20757 39071 20791
rect 39071 20757 39080 20791
rect 39028 20748 39080 20757
rect 39764 20748 39816 20800
rect 43812 20791 43864 20800
rect 43812 20757 43821 20791
rect 43821 20757 43855 20791
rect 43855 20757 43864 20791
rect 43812 20748 43864 20757
rect 45008 20748 45060 20800
rect 47492 20791 47544 20800
rect 47492 20757 47501 20791
rect 47501 20757 47535 20791
rect 47535 20757 47544 20791
rect 47492 20748 47544 20757
rect 55956 20952 56008 21004
rect 57520 20927 57572 20936
rect 57520 20893 57529 20927
rect 57529 20893 57563 20927
rect 57563 20893 57572 20927
rect 57520 20884 57572 20893
rect 49332 20748 49384 20800
rect 50896 20791 50948 20800
rect 50896 20757 50905 20791
rect 50905 20757 50939 20791
rect 50939 20757 50948 20791
rect 50896 20748 50948 20757
rect 51908 20791 51960 20800
rect 51908 20757 51917 20791
rect 51917 20757 51951 20791
rect 51951 20757 51960 20791
rect 51908 20748 51960 20757
rect 52552 20791 52604 20800
rect 52552 20757 52561 20791
rect 52561 20757 52595 20791
rect 52595 20757 52604 20791
rect 52552 20748 52604 20757
rect 52920 20791 52972 20800
rect 52920 20757 52929 20791
rect 52929 20757 52963 20791
rect 52963 20757 52972 20791
rect 52920 20748 52972 20757
rect 53012 20791 53064 20800
rect 53012 20757 53021 20791
rect 53021 20757 53055 20791
rect 53055 20757 53064 20791
rect 53012 20748 53064 20757
rect 53748 20791 53800 20800
rect 53748 20757 53757 20791
rect 53757 20757 53791 20791
rect 53791 20757 53800 20791
rect 53748 20748 53800 20757
rect 55036 20791 55088 20800
rect 55036 20757 55045 20791
rect 55045 20757 55079 20791
rect 55079 20757 55088 20791
rect 55036 20748 55088 20757
rect 55588 20748 55640 20800
rect 56140 20791 56192 20800
rect 56140 20757 56149 20791
rect 56149 20757 56183 20791
rect 56183 20757 56192 20791
rect 56140 20748 56192 20757
rect 56784 20816 56836 20868
rect 15394 20646 15446 20698
rect 15458 20646 15510 20698
rect 15522 20646 15574 20698
rect 15586 20646 15638 20698
rect 15650 20646 15702 20698
rect 29838 20646 29890 20698
rect 29902 20646 29954 20698
rect 29966 20646 30018 20698
rect 30030 20646 30082 20698
rect 30094 20646 30146 20698
rect 44282 20646 44334 20698
rect 44346 20646 44398 20698
rect 44410 20646 44462 20698
rect 44474 20646 44526 20698
rect 44538 20646 44590 20698
rect 58726 20646 58778 20698
rect 58790 20646 58842 20698
rect 58854 20646 58906 20698
rect 58918 20646 58970 20698
rect 58982 20646 59034 20698
rect 8576 20544 8628 20596
rect 4988 20476 5040 20528
rect 9128 20544 9180 20596
rect 11612 20544 11664 20596
rect 12256 20544 12308 20596
rect 4160 20340 4212 20392
rect 4252 20340 4304 20392
rect 7564 20383 7616 20392
rect 7564 20349 7573 20383
rect 7573 20349 7607 20383
rect 7607 20349 7616 20383
rect 7564 20340 7616 20349
rect 7656 20340 7708 20392
rect 6552 20272 6604 20324
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 9496 20408 9548 20460
rect 10140 20408 10192 20460
rect 10876 20476 10928 20528
rect 11060 20476 11112 20528
rect 14372 20544 14424 20596
rect 8760 20340 8812 20349
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 11704 20408 11756 20460
rect 13452 20408 13504 20460
rect 15200 20544 15252 20596
rect 16028 20544 16080 20596
rect 18604 20587 18656 20596
rect 18604 20553 18613 20587
rect 18613 20553 18647 20587
rect 18647 20553 18656 20587
rect 18604 20544 18656 20553
rect 19248 20544 19300 20596
rect 19800 20544 19852 20596
rect 20536 20544 20588 20596
rect 22100 20544 22152 20596
rect 25872 20544 25924 20596
rect 28356 20587 28408 20596
rect 18052 20476 18104 20528
rect 15936 20408 15988 20460
rect 20536 20451 20588 20460
rect 20536 20417 20554 20451
rect 20554 20417 20588 20451
rect 20536 20408 20588 20417
rect 21456 20408 21508 20460
rect 23572 20408 23624 20460
rect 25596 20451 25648 20460
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 25872 20451 25924 20460
rect 25872 20417 25881 20451
rect 25881 20417 25915 20451
rect 25915 20417 25924 20451
rect 25872 20408 25924 20417
rect 28356 20553 28365 20587
rect 28365 20553 28399 20587
rect 28399 20553 28408 20587
rect 28356 20544 28408 20553
rect 28632 20544 28684 20596
rect 30748 20544 30800 20596
rect 27252 20519 27304 20528
rect 27252 20485 27286 20519
rect 27286 20485 27304 20519
rect 27252 20476 27304 20485
rect 27896 20476 27948 20528
rect 30196 20476 30248 20528
rect 31208 20544 31260 20596
rect 31392 20544 31444 20596
rect 31852 20544 31904 20596
rect 27712 20408 27764 20460
rect 32128 20476 32180 20528
rect 35256 20544 35308 20596
rect 37648 20544 37700 20596
rect 37924 20544 37976 20596
rect 38476 20544 38528 20596
rect 38844 20544 38896 20596
rect 39948 20587 40000 20596
rect 39948 20553 39957 20587
rect 39957 20553 39991 20587
rect 39991 20553 40000 20587
rect 39948 20544 40000 20553
rect 40040 20587 40092 20596
rect 40040 20553 40049 20587
rect 40049 20553 40083 20587
rect 40083 20553 40092 20587
rect 40040 20544 40092 20553
rect 41880 20544 41932 20596
rect 44180 20544 44232 20596
rect 34520 20476 34572 20528
rect 12072 20340 12124 20392
rect 8116 20315 8168 20324
rect 8116 20281 8125 20315
rect 8125 20281 8159 20315
rect 8159 20281 8168 20315
rect 8116 20272 8168 20281
rect 13176 20340 13228 20392
rect 13360 20383 13412 20392
rect 13360 20349 13369 20383
rect 13369 20349 13403 20383
rect 13403 20349 13412 20383
rect 13360 20340 13412 20349
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 13820 20272 13872 20324
rect 14096 20272 14148 20324
rect 18696 20340 18748 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 20352 20383 20404 20392
rect 20352 20349 20363 20383
rect 20363 20349 20397 20383
rect 20397 20349 20404 20383
rect 20352 20340 20404 20349
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 21732 20340 21784 20392
rect 12164 20204 12216 20256
rect 12624 20247 12676 20256
rect 12624 20213 12633 20247
rect 12633 20213 12667 20247
rect 12667 20213 12676 20247
rect 12624 20204 12676 20213
rect 14464 20204 14516 20256
rect 19800 20272 19852 20324
rect 20812 20272 20864 20324
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 23480 20383 23532 20392
rect 23480 20349 23489 20383
rect 23489 20349 23523 20383
rect 23523 20349 23532 20383
rect 23480 20340 23532 20349
rect 25780 20383 25832 20392
rect 25780 20349 25798 20383
rect 25798 20349 25832 20383
rect 25780 20340 25832 20349
rect 26148 20315 26200 20324
rect 26148 20281 26157 20315
rect 26157 20281 26191 20315
rect 26191 20281 26200 20315
rect 26148 20272 26200 20281
rect 28908 20383 28960 20392
rect 28908 20349 28917 20383
rect 28917 20349 28951 20383
rect 28951 20349 28960 20383
rect 28908 20340 28960 20349
rect 29000 20383 29052 20392
rect 29000 20349 29009 20383
rect 29009 20349 29043 20383
rect 29043 20349 29052 20383
rect 29000 20340 29052 20349
rect 31484 20451 31536 20460
rect 31484 20417 31493 20451
rect 31493 20417 31527 20451
rect 31527 20417 31536 20451
rect 31484 20408 31536 20417
rect 31668 20408 31720 20460
rect 32956 20451 33008 20460
rect 32956 20417 32965 20451
rect 32965 20417 32999 20451
rect 32999 20417 33008 20451
rect 32956 20408 33008 20417
rect 33784 20408 33836 20460
rect 34152 20451 34204 20460
rect 34152 20417 34161 20451
rect 34161 20417 34195 20451
rect 34195 20417 34204 20451
rect 34152 20408 34204 20417
rect 28172 20272 28224 20324
rect 31576 20272 31628 20324
rect 33232 20383 33284 20392
rect 33232 20349 33241 20383
rect 33241 20349 33275 20383
rect 33275 20349 33284 20383
rect 33232 20340 33284 20349
rect 33508 20383 33560 20392
rect 33508 20349 33517 20383
rect 33517 20349 33551 20383
rect 33551 20349 33560 20383
rect 33508 20340 33560 20349
rect 33876 20340 33928 20392
rect 33600 20272 33652 20324
rect 34704 20408 34756 20460
rect 35716 20451 35768 20460
rect 35716 20417 35725 20451
rect 35725 20417 35759 20451
rect 35759 20417 35768 20451
rect 35716 20408 35768 20417
rect 35992 20451 36044 20460
rect 35992 20417 36026 20451
rect 36026 20417 36044 20451
rect 35992 20408 36044 20417
rect 42708 20519 42760 20528
rect 42708 20485 42742 20519
rect 42742 20485 42760 20519
rect 42708 20476 42760 20485
rect 43076 20476 43128 20528
rect 48228 20544 48280 20596
rect 46756 20476 46808 20528
rect 46940 20476 46992 20528
rect 50896 20476 50948 20528
rect 38384 20451 38436 20460
rect 38384 20417 38393 20451
rect 38393 20417 38427 20451
rect 38427 20417 38436 20451
rect 38384 20408 38436 20417
rect 39856 20408 39908 20460
rect 45744 20408 45796 20460
rect 48320 20408 48372 20460
rect 49424 20451 49476 20460
rect 49424 20417 49433 20451
rect 49433 20417 49467 20451
rect 49467 20417 49476 20451
rect 49424 20408 49476 20417
rect 38660 20383 38712 20392
rect 38660 20349 38669 20383
rect 38669 20349 38703 20383
rect 38703 20349 38712 20383
rect 38660 20340 38712 20349
rect 38844 20340 38896 20392
rect 35532 20272 35584 20324
rect 39764 20383 39816 20392
rect 39764 20349 39773 20383
rect 39773 20349 39807 20383
rect 39807 20349 39816 20383
rect 39764 20340 39816 20349
rect 40040 20340 40092 20392
rect 42432 20383 42484 20392
rect 42432 20349 42441 20383
rect 42441 20349 42475 20383
rect 42475 20349 42484 20383
rect 42432 20340 42484 20349
rect 45928 20383 45980 20392
rect 45928 20349 45937 20383
rect 45937 20349 45971 20383
rect 45971 20349 45980 20383
rect 45928 20340 45980 20349
rect 16120 20204 16172 20256
rect 21364 20204 21416 20256
rect 26240 20204 26292 20256
rect 26976 20204 27028 20256
rect 34704 20204 34756 20256
rect 34980 20247 35032 20256
rect 34980 20213 34989 20247
rect 34989 20213 35023 20247
rect 35023 20213 35032 20247
rect 34980 20204 35032 20213
rect 38844 20204 38896 20256
rect 39580 20204 39632 20256
rect 45008 20204 45060 20256
rect 47584 20247 47636 20256
rect 47584 20213 47593 20247
rect 47593 20213 47627 20247
rect 47627 20213 47636 20247
rect 47584 20204 47636 20213
rect 47676 20204 47728 20256
rect 47768 20204 47820 20256
rect 51908 20544 51960 20596
rect 53012 20476 53064 20528
rect 53748 20476 53800 20528
rect 52552 20408 52604 20460
rect 54668 20451 54720 20460
rect 54668 20417 54686 20451
rect 54686 20417 54720 20451
rect 54668 20408 54720 20417
rect 56048 20519 56100 20528
rect 56048 20485 56082 20519
rect 56082 20485 56100 20519
rect 56048 20476 56100 20485
rect 57520 20544 57572 20596
rect 48872 20272 48924 20324
rect 52828 20383 52880 20392
rect 52828 20349 52837 20383
rect 52837 20349 52871 20383
rect 52871 20349 52880 20383
rect 52828 20340 52880 20349
rect 53012 20383 53064 20392
rect 53012 20349 53021 20383
rect 53021 20349 53055 20383
rect 53055 20349 53064 20383
rect 53012 20340 53064 20349
rect 53840 20340 53892 20392
rect 54484 20383 54536 20392
rect 54484 20349 54493 20383
rect 54493 20349 54527 20383
rect 54527 20349 54536 20383
rect 54484 20340 54536 20349
rect 54760 20383 54812 20392
rect 54760 20349 54769 20383
rect 54769 20349 54803 20383
rect 54803 20349 54812 20383
rect 54760 20340 54812 20349
rect 55404 20340 55456 20392
rect 55496 20383 55548 20392
rect 55496 20349 55505 20383
rect 55505 20349 55539 20383
rect 55539 20349 55548 20383
rect 55496 20340 55548 20349
rect 53472 20315 53524 20324
rect 53472 20281 53481 20315
rect 53481 20281 53515 20315
rect 53515 20281 53524 20315
rect 53472 20272 53524 20281
rect 54944 20272 54996 20324
rect 50712 20204 50764 20256
rect 55772 20204 55824 20256
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 22616 20102 22668 20154
rect 22680 20102 22732 20154
rect 22744 20102 22796 20154
rect 22808 20102 22860 20154
rect 22872 20102 22924 20154
rect 37060 20102 37112 20154
rect 37124 20102 37176 20154
rect 37188 20102 37240 20154
rect 37252 20102 37304 20154
rect 37316 20102 37368 20154
rect 51504 20102 51556 20154
rect 51568 20102 51620 20154
rect 51632 20102 51684 20154
rect 51696 20102 51748 20154
rect 51760 20102 51812 20154
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 7656 20000 7708 20052
rect 8760 20000 8812 20052
rect 10140 20000 10192 20052
rect 12808 20000 12860 20052
rect 13636 20000 13688 20052
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 4252 19796 4304 19848
rect 4436 19771 4488 19780
rect 4436 19737 4470 19771
rect 4470 19737 4488 19771
rect 4436 19728 4488 19737
rect 12072 19932 12124 19984
rect 15752 20000 15804 20052
rect 18236 20000 18288 20052
rect 20628 20000 20680 20052
rect 21732 20043 21784 20052
rect 21732 20009 21741 20043
rect 21741 20009 21775 20043
rect 21775 20009 21784 20043
rect 21732 20000 21784 20009
rect 23572 20043 23624 20052
rect 23572 20009 23581 20043
rect 23581 20009 23615 20043
rect 23615 20009 23624 20043
rect 23572 20000 23624 20009
rect 25044 20000 25096 20052
rect 27712 20043 27764 20052
rect 27712 20009 27721 20043
rect 27721 20009 27755 20043
rect 27755 20009 27764 20043
rect 27712 20000 27764 20009
rect 28908 20000 28960 20052
rect 30840 20000 30892 20052
rect 7288 19728 7340 19780
rect 7656 19728 7708 19780
rect 9772 19796 9824 19848
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 12440 19864 12492 19916
rect 17132 19907 17184 19916
rect 17132 19873 17141 19907
rect 17141 19873 17175 19907
rect 17175 19873 17184 19907
rect 17132 19864 17184 19873
rect 10876 19796 10928 19805
rect 15936 19796 15988 19848
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 21456 19864 21508 19916
rect 20076 19796 20128 19848
rect 21548 19796 21600 19848
rect 23756 19864 23808 19916
rect 33232 20000 33284 20052
rect 34152 20000 34204 20052
rect 34612 20000 34664 20052
rect 38660 20000 38712 20052
rect 39028 20000 39080 20052
rect 43260 20000 43312 20052
rect 43996 20000 44048 20052
rect 47768 20000 47820 20052
rect 35716 19864 35768 19916
rect 43720 19975 43772 19984
rect 43720 19941 43729 19975
rect 43729 19941 43763 19975
rect 43763 19941 43772 19975
rect 43720 19932 43772 19941
rect 11520 19728 11572 19780
rect 12624 19728 12676 19780
rect 13360 19728 13412 19780
rect 15752 19728 15804 19780
rect 17592 19728 17644 19780
rect 9128 19660 9180 19712
rect 9864 19660 9916 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 14556 19660 14608 19712
rect 19892 19660 19944 19712
rect 20352 19660 20404 19712
rect 20720 19660 20772 19712
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 25228 19728 25280 19780
rect 28080 19796 28132 19848
rect 29644 19796 29696 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 26976 19728 27028 19780
rect 35256 19839 35308 19848
rect 35256 19805 35265 19839
rect 35265 19805 35299 19839
rect 35299 19805 35308 19839
rect 35256 19796 35308 19805
rect 35532 19796 35584 19848
rect 39580 19864 39632 19916
rect 40500 19864 40552 19916
rect 43352 19907 43404 19916
rect 43352 19873 43361 19907
rect 43361 19873 43395 19907
rect 43395 19873 43404 19907
rect 43352 19864 43404 19873
rect 43628 19864 43680 19916
rect 43812 19864 43864 19916
rect 47584 19932 47636 19984
rect 49056 20000 49108 20052
rect 49424 20000 49476 20052
rect 44640 19864 44692 19916
rect 47492 19907 47544 19916
rect 47492 19873 47501 19907
rect 47501 19873 47535 19907
rect 47535 19873 47544 19907
rect 47492 19864 47544 19873
rect 50712 19907 50764 19916
rect 50712 19873 50721 19907
rect 50721 19873 50755 19907
rect 50755 19873 50764 19907
rect 50712 19864 50764 19873
rect 51908 20000 51960 20052
rect 52828 20000 52880 20052
rect 55496 20000 55548 20052
rect 53380 19932 53432 19984
rect 54760 19932 54812 19984
rect 39672 19796 39724 19848
rect 33508 19728 33560 19780
rect 24768 19703 24820 19712
rect 24768 19669 24777 19703
rect 24777 19669 24811 19703
rect 24811 19669 24820 19703
rect 24768 19660 24820 19669
rect 25780 19660 25832 19712
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 34336 19703 34388 19712
rect 34336 19669 34345 19703
rect 34345 19669 34379 19703
rect 34379 19669 34388 19703
rect 34336 19660 34388 19669
rect 35348 19660 35400 19712
rect 37280 19728 37332 19780
rect 38752 19728 38804 19780
rect 39212 19660 39264 19712
rect 43076 19796 43128 19848
rect 44824 19796 44876 19848
rect 45008 19796 45060 19848
rect 45928 19796 45980 19848
rect 47400 19796 47452 19848
rect 48964 19796 49016 19848
rect 52920 19864 52972 19916
rect 56784 20043 56836 20052
rect 56784 20009 56793 20043
rect 56793 20009 56827 20043
rect 56827 20009 56836 20043
rect 56784 20000 56836 20009
rect 55404 19796 55456 19848
rect 42984 19660 43036 19712
rect 48504 19728 48556 19780
rect 55864 19728 55916 19780
rect 48320 19660 48372 19712
rect 50160 19703 50212 19712
rect 50160 19669 50169 19703
rect 50169 19669 50203 19703
rect 50203 19669 50212 19703
rect 50160 19660 50212 19669
rect 53380 19660 53432 19712
rect 54300 19703 54352 19712
rect 54300 19669 54309 19703
rect 54309 19669 54343 19703
rect 54343 19669 54352 19703
rect 54300 19660 54352 19669
rect 54944 19660 54996 19712
rect 15394 19558 15446 19610
rect 15458 19558 15510 19610
rect 15522 19558 15574 19610
rect 15586 19558 15638 19610
rect 15650 19558 15702 19610
rect 29838 19558 29890 19610
rect 29902 19558 29954 19610
rect 29966 19558 30018 19610
rect 30030 19558 30082 19610
rect 30094 19558 30146 19610
rect 44282 19558 44334 19610
rect 44346 19558 44398 19610
rect 44410 19558 44462 19610
rect 44474 19558 44526 19610
rect 44538 19558 44590 19610
rect 58726 19558 58778 19610
rect 58790 19558 58842 19610
rect 58854 19558 58906 19610
rect 58918 19558 58970 19610
rect 58982 19558 59034 19610
rect 7656 19499 7708 19508
rect 7656 19465 7665 19499
rect 7665 19465 7699 19499
rect 7699 19465 7708 19499
rect 7656 19456 7708 19465
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 10968 19456 11020 19508
rect 14556 19499 14608 19508
rect 14556 19465 14565 19499
rect 14565 19465 14599 19499
rect 14599 19465 14608 19499
rect 14556 19456 14608 19465
rect 15752 19499 15804 19508
rect 15752 19465 15761 19499
rect 15761 19465 15795 19499
rect 15795 19465 15804 19499
rect 15752 19456 15804 19465
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 22560 19456 22612 19508
rect 23664 19456 23716 19508
rect 25780 19456 25832 19508
rect 33508 19456 33560 19508
rect 33968 19456 34020 19508
rect 35256 19456 35308 19508
rect 37280 19499 37332 19508
rect 37280 19465 37289 19499
rect 37289 19465 37323 19499
rect 37323 19465 37332 19499
rect 37280 19456 37332 19465
rect 38752 19499 38804 19508
rect 38752 19465 38761 19499
rect 38761 19465 38795 19499
rect 38795 19465 38804 19499
rect 38752 19456 38804 19465
rect 39672 19499 39724 19508
rect 39672 19465 39681 19499
rect 39681 19465 39715 19499
rect 39715 19465 39724 19499
rect 39672 19456 39724 19465
rect 43352 19456 43404 19508
rect 48780 19456 48832 19508
rect 48964 19499 49016 19508
rect 48964 19465 48973 19499
rect 48973 19465 49007 19499
rect 49007 19465 49016 19499
rect 48964 19456 49016 19465
rect 50160 19456 50212 19508
rect 55404 19456 55456 19508
rect 55864 19499 55916 19508
rect 55864 19465 55873 19499
rect 55873 19465 55907 19499
rect 55907 19465 55916 19499
rect 55864 19456 55916 19465
rect 22284 19388 22336 19440
rect 22468 19388 22520 19440
rect 7012 19363 7064 19372
rect 7012 19329 7021 19363
rect 7021 19329 7055 19363
rect 7055 19329 7064 19363
rect 7012 19320 7064 19329
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 13728 19320 13780 19372
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 4620 19295 4672 19304
rect 4620 19261 4629 19295
rect 4629 19261 4663 19295
rect 4663 19261 4672 19295
rect 4620 19252 4672 19261
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 7748 19252 7800 19304
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 11336 19252 11388 19304
rect 9404 19184 9456 19236
rect 3516 19159 3568 19168
rect 3516 19125 3525 19159
rect 3525 19125 3559 19159
rect 3559 19125 3568 19159
rect 3516 19116 3568 19125
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 11520 19159 11572 19168
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 13544 19252 13596 19304
rect 14832 19320 14884 19372
rect 14188 19184 14240 19236
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 44640 19388 44692 19440
rect 15292 19252 15344 19304
rect 17132 19252 17184 19304
rect 17776 19252 17828 19304
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 19340 19252 19392 19261
rect 19708 19227 19760 19236
rect 19708 19193 19717 19227
rect 19717 19193 19751 19227
rect 19751 19193 19760 19227
rect 19708 19184 19760 19193
rect 22468 19252 22520 19304
rect 34980 19320 35032 19372
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 26148 19252 26200 19304
rect 27988 19295 28040 19304
rect 27988 19261 27997 19295
rect 27997 19261 28031 19295
rect 28031 19261 28040 19295
rect 27988 19252 28040 19261
rect 28540 19252 28592 19304
rect 31116 19295 31168 19304
rect 31116 19261 31125 19295
rect 31125 19261 31159 19295
rect 31159 19261 31168 19295
rect 31116 19252 31168 19261
rect 21180 19116 21232 19168
rect 22836 19116 22888 19168
rect 23388 19116 23440 19168
rect 33600 19295 33652 19304
rect 33600 19261 33609 19295
rect 33609 19261 33643 19295
rect 33643 19261 33652 19295
rect 33600 19252 33652 19261
rect 34336 19252 34388 19304
rect 40040 19320 40092 19372
rect 44088 19363 44140 19372
rect 44088 19329 44097 19363
rect 44097 19329 44131 19363
rect 44131 19329 44140 19363
rect 44088 19320 44140 19329
rect 44180 19320 44232 19372
rect 45284 19320 45336 19372
rect 38108 19252 38160 19304
rect 38568 19252 38620 19304
rect 38660 19295 38712 19304
rect 38660 19261 38669 19295
rect 38669 19261 38703 19295
rect 38703 19261 38712 19295
rect 38660 19252 38712 19261
rect 42248 19295 42300 19304
rect 42248 19261 42257 19295
rect 42257 19261 42291 19295
rect 42291 19261 42300 19295
rect 42248 19252 42300 19261
rect 42708 19252 42760 19304
rect 43260 19295 43312 19304
rect 43260 19261 43278 19295
rect 43278 19261 43312 19295
rect 43260 19252 43312 19261
rect 43628 19227 43680 19236
rect 43628 19193 43637 19227
rect 43637 19193 43671 19227
rect 43671 19193 43680 19227
rect 43628 19184 43680 19193
rect 46020 19295 46072 19304
rect 46020 19261 46029 19295
rect 46029 19261 46063 19295
rect 46063 19261 46072 19295
rect 46020 19252 46072 19261
rect 48320 19252 48372 19304
rect 48780 19252 48832 19304
rect 49332 19320 49384 19372
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 27436 19159 27488 19168
rect 27436 19125 27445 19159
rect 27445 19125 27479 19159
rect 27479 19125 27488 19159
rect 27436 19116 27488 19125
rect 28264 19159 28316 19168
rect 28264 19125 28273 19159
rect 28273 19125 28307 19159
rect 28307 19125 28316 19159
rect 28264 19116 28316 19125
rect 30564 19159 30616 19168
rect 30564 19125 30573 19159
rect 30573 19125 30607 19159
rect 30607 19125 30616 19159
rect 30564 19116 30616 19125
rect 31576 19159 31628 19168
rect 31576 19125 31585 19159
rect 31585 19125 31619 19159
rect 31619 19125 31628 19159
rect 31576 19116 31628 19125
rect 31944 19116 31996 19168
rect 32772 19116 32824 19168
rect 33140 19159 33192 19168
rect 33140 19125 33149 19159
rect 33149 19125 33183 19159
rect 33183 19125 33192 19159
rect 33140 19116 33192 19125
rect 34888 19116 34940 19168
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 38016 19159 38068 19168
rect 38016 19125 38025 19159
rect 38025 19125 38059 19159
rect 38059 19125 38068 19159
rect 38016 19116 38068 19125
rect 41604 19159 41656 19168
rect 41604 19125 41613 19159
rect 41613 19125 41647 19159
rect 41647 19125 41656 19159
rect 41604 19116 41656 19125
rect 43720 19116 43772 19168
rect 43812 19116 43864 19168
rect 44180 19116 44232 19168
rect 45744 19184 45796 19236
rect 49700 19184 49752 19236
rect 44916 19116 44968 19168
rect 47676 19116 47728 19168
rect 48228 19159 48280 19168
rect 48228 19125 48237 19159
rect 48237 19125 48271 19159
rect 48271 19125 48280 19159
rect 48228 19116 48280 19125
rect 48596 19159 48648 19168
rect 48596 19125 48605 19159
rect 48605 19125 48639 19159
rect 48639 19125 48648 19159
rect 48596 19116 48648 19125
rect 51264 19388 51316 19440
rect 56140 19252 56192 19304
rect 51356 19116 51408 19168
rect 52184 19159 52236 19168
rect 52184 19125 52193 19159
rect 52193 19125 52227 19159
rect 52227 19125 52236 19159
rect 52184 19116 52236 19125
rect 52552 19116 52604 19168
rect 52920 19159 52972 19168
rect 52920 19125 52929 19159
rect 52929 19125 52963 19159
rect 52963 19125 52972 19159
rect 52920 19116 52972 19125
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 22616 19014 22668 19066
rect 22680 19014 22732 19066
rect 22744 19014 22796 19066
rect 22808 19014 22860 19066
rect 22872 19014 22924 19066
rect 37060 19014 37112 19066
rect 37124 19014 37176 19066
rect 37188 19014 37240 19066
rect 37252 19014 37304 19066
rect 37316 19014 37368 19066
rect 51504 19014 51556 19066
rect 51568 19014 51620 19066
rect 51632 19014 51684 19066
rect 51696 19014 51748 19066
rect 51760 19014 51812 19066
rect 4620 18912 4672 18964
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 7104 18912 7156 18964
rect 8024 18912 8076 18964
rect 11244 18912 11296 18964
rect 4712 18844 4764 18896
rect 10324 18844 10376 18896
rect 4436 18776 4488 18828
rect 6460 18776 6512 18828
rect 10048 18819 10100 18828
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 11704 18912 11756 18964
rect 13544 18912 13596 18964
rect 6368 18708 6420 18760
rect 8576 18708 8628 18760
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 13912 18844 13964 18896
rect 12900 18776 12952 18828
rect 17960 18844 18012 18896
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 5816 18572 5868 18624
rect 6460 18572 6512 18624
rect 9128 18572 9180 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 10416 18615 10468 18624
rect 10416 18581 10425 18615
rect 10425 18581 10459 18615
rect 10459 18581 10468 18615
rect 10416 18572 10468 18581
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 12808 18572 12860 18624
rect 18236 18819 18288 18828
rect 18236 18785 18245 18819
rect 18245 18785 18279 18819
rect 18279 18785 18288 18819
rect 18236 18776 18288 18785
rect 19708 18776 19760 18828
rect 19984 18819 20036 18828
rect 19984 18785 19993 18819
rect 19993 18785 20027 18819
rect 20027 18785 20036 18819
rect 19984 18776 20036 18785
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 14924 18751 14976 18760
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 18696 18708 18748 18760
rect 19064 18751 19116 18760
rect 19064 18717 19073 18751
rect 19073 18717 19107 18751
rect 19107 18717 19116 18751
rect 19064 18708 19116 18717
rect 14004 18640 14056 18692
rect 20812 18708 20864 18760
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 14096 18572 14148 18624
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 15752 18572 15804 18624
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 18328 18572 18380 18624
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 18788 18572 18840 18624
rect 20260 18683 20312 18692
rect 20260 18649 20294 18683
rect 20294 18649 20312 18683
rect 20260 18640 20312 18649
rect 27988 18912 28040 18964
rect 31116 18912 31168 18964
rect 22100 18844 22152 18896
rect 21180 18776 21232 18828
rect 30932 18844 30984 18896
rect 31576 18844 31628 18896
rect 36912 18912 36964 18964
rect 39672 18912 39724 18964
rect 21916 18708 21968 18760
rect 22284 18708 22336 18760
rect 25228 18708 25280 18760
rect 26240 18708 26292 18760
rect 27252 18776 27304 18828
rect 28264 18708 28316 18760
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 28908 18708 28960 18760
rect 27896 18683 27948 18692
rect 27896 18649 27905 18683
rect 27905 18649 27939 18683
rect 27939 18649 27948 18683
rect 27896 18640 27948 18649
rect 28724 18640 28776 18692
rect 20352 18572 20404 18624
rect 20904 18572 20956 18624
rect 21732 18615 21784 18624
rect 21732 18581 21741 18615
rect 21741 18581 21775 18615
rect 21775 18581 21784 18615
rect 21732 18572 21784 18581
rect 21824 18615 21876 18624
rect 21824 18581 21833 18615
rect 21833 18581 21867 18615
rect 21867 18581 21876 18615
rect 21824 18572 21876 18581
rect 22192 18572 22244 18624
rect 23572 18615 23624 18624
rect 23572 18581 23581 18615
rect 23581 18581 23615 18615
rect 23615 18581 23624 18615
rect 23572 18572 23624 18581
rect 24768 18615 24820 18624
rect 24768 18581 24777 18615
rect 24777 18581 24811 18615
rect 24811 18581 24820 18615
rect 24768 18572 24820 18581
rect 25872 18572 25924 18624
rect 26240 18572 26292 18624
rect 27068 18615 27120 18624
rect 27068 18581 27077 18615
rect 27077 18581 27111 18615
rect 27111 18581 27120 18615
rect 27068 18572 27120 18581
rect 27252 18572 27304 18624
rect 28264 18615 28316 18624
rect 28264 18581 28273 18615
rect 28273 18581 28307 18615
rect 28307 18581 28316 18615
rect 28264 18572 28316 18581
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 33140 18776 33192 18828
rect 34888 18819 34940 18828
rect 34888 18785 34897 18819
rect 34897 18785 34931 18819
rect 34931 18785 34940 18819
rect 34888 18776 34940 18785
rect 35164 18776 35216 18828
rect 38016 18776 38068 18828
rect 41420 18912 41472 18964
rect 42248 18912 42300 18964
rect 43628 18912 43680 18964
rect 46020 18912 46072 18964
rect 54300 18912 54352 18964
rect 43076 18776 43128 18828
rect 43812 18776 43864 18828
rect 46756 18776 46808 18828
rect 31944 18708 31996 18760
rect 32036 18751 32088 18760
rect 32036 18717 32045 18751
rect 32045 18717 32079 18751
rect 32079 18717 32088 18751
rect 32036 18708 32088 18717
rect 31484 18640 31536 18692
rect 33600 18708 33652 18760
rect 31116 18572 31168 18624
rect 31576 18615 31628 18624
rect 31576 18581 31585 18615
rect 31585 18581 31619 18615
rect 31619 18581 31628 18615
rect 31576 18572 31628 18581
rect 34244 18751 34296 18760
rect 34244 18717 34253 18751
rect 34253 18717 34287 18751
rect 34287 18717 34296 18751
rect 34244 18708 34296 18717
rect 35900 18708 35952 18760
rect 36820 18751 36872 18760
rect 36820 18717 36829 18751
rect 36829 18717 36863 18751
rect 36863 18717 36872 18751
rect 36820 18708 36872 18717
rect 37740 18708 37792 18760
rect 43996 18751 44048 18760
rect 43996 18717 44005 18751
rect 44005 18717 44039 18751
rect 44039 18717 44048 18751
rect 43996 18708 44048 18717
rect 47584 18844 47636 18896
rect 48228 18844 48280 18896
rect 47492 18776 47544 18828
rect 47032 18751 47084 18760
rect 47032 18717 47041 18751
rect 47041 18717 47075 18751
rect 47075 18717 47084 18751
rect 47032 18708 47084 18717
rect 48596 18776 48648 18828
rect 58164 18844 58216 18896
rect 41144 18640 41196 18692
rect 41604 18640 41656 18692
rect 48136 18640 48188 18692
rect 49056 18751 49108 18760
rect 49056 18717 49065 18751
rect 49065 18717 49099 18751
rect 49099 18717 49108 18751
rect 49056 18708 49108 18717
rect 49332 18708 49384 18760
rect 50344 18751 50396 18760
rect 50344 18717 50353 18751
rect 50353 18717 50387 18751
rect 50387 18717 50396 18751
rect 50344 18708 50396 18717
rect 56324 18776 56376 18828
rect 53656 18751 53708 18760
rect 53656 18717 53665 18751
rect 53665 18717 53699 18751
rect 53699 18717 53708 18751
rect 53656 18708 53708 18717
rect 55772 18751 55824 18760
rect 55772 18717 55781 18751
rect 55781 18717 55815 18751
rect 55815 18717 55824 18751
rect 55772 18708 55824 18717
rect 56600 18708 56652 18760
rect 32956 18572 33008 18624
rect 33600 18615 33652 18624
rect 33600 18581 33609 18615
rect 33609 18581 33643 18615
rect 33643 18581 33652 18615
rect 33600 18572 33652 18581
rect 35532 18615 35584 18624
rect 35532 18581 35541 18615
rect 35541 18581 35575 18615
rect 35575 18581 35584 18615
rect 35532 18572 35584 18581
rect 37556 18572 37608 18624
rect 37832 18615 37884 18624
rect 37832 18581 37841 18615
rect 37841 18581 37875 18615
rect 37875 18581 37884 18615
rect 37832 18572 37884 18581
rect 39212 18615 39264 18624
rect 39212 18581 39221 18615
rect 39221 18581 39255 18615
rect 39255 18581 39264 18615
rect 39212 18572 39264 18581
rect 39580 18615 39632 18624
rect 39580 18581 39589 18615
rect 39589 18581 39623 18615
rect 39623 18581 39632 18615
rect 39580 18572 39632 18581
rect 42064 18572 42116 18624
rect 42984 18615 43036 18624
rect 42984 18581 42993 18615
rect 42993 18581 43027 18615
rect 43027 18581 43036 18615
rect 42984 18572 43036 18581
rect 46020 18615 46072 18624
rect 46020 18581 46029 18615
rect 46029 18581 46063 18615
rect 46063 18581 46072 18615
rect 46020 18572 46072 18581
rect 46204 18572 46256 18624
rect 46388 18615 46440 18624
rect 46388 18581 46397 18615
rect 46397 18581 46431 18615
rect 46431 18581 46440 18615
rect 46388 18572 46440 18581
rect 46664 18572 46716 18624
rect 48412 18572 48464 18624
rect 52184 18640 52236 18692
rect 53012 18640 53064 18692
rect 48872 18572 48924 18624
rect 48964 18615 49016 18624
rect 48964 18581 48973 18615
rect 48973 18581 49007 18615
rect 49007 18581 49016 18615
rect 48964 18572 49016 18581
rect 49148 18572 49200 18624
rect 50988 18615 51040 18624
rect 50988 18581 50997 18615
rect 50997 18581 51031 18615
rect 51031 18581 51040 18615
rect 50988 18572 51040 18581
rect 51908 18572 51960 18624
rect 52736 18615 52788 18624
rect 52736 18581 52745 18615
rect 52745 18581 52779 18615
rect 52779 18581 52788 18615
rect 52736 18572 52788 18581
rect 52828 18572 52880 18624
rect 54576 18572 54628 18624
rect 55588 18572 55640 18624
rect 55680 18615 55732 18624
rect 55680 18581 55689 18615
rect 55689 18581 55723 18615
rect 55723 18581 55732 18615
rect 55680 18572 55732 18581
rect 56232 18615 56284 18624
rect 56232 18581 56241 18615
rect 56241 18581 56275 18615
rect 56275 18581 56284 18615
rect 56232 18572 56284 18581
rect 56968 18615 57020 18624
rect 56968 18581 56977 18615
rect 56977 18581 57011 18615
rect 57011 18581 57020 18615
rect 56968 18572 57020 18581
rect 57244 18572 57296 18624
rect 15394 18470 15446 18522
rect 15458 18470 15510 18522
rect 15522 18470 15574 18522
rect 15586 18470 15638 18522
rect 15650 18470 15702 18522
rect 29838 18470 29890 18522
rect 29902 18470 29954 18522
rect 29966 18470 30018 18522
rect 30030 18470 30082 18522
rect 30094 18470 30146 18522
rect 44282 18470 44334 18522
rect 44346 18470 44398 18522
rect 44410 18470 44462 18522
rect 44474 18470 44526 18522
rect 44538 18470 44590 18522
rect 58726 18470 58778 18522
rect 58790 18470 58842 18522
rect 58854 18470 58906 18522
rect 58918 18470 58970 18522
rect 58982 18470 59034 18522
rect 5264 18300 5316 18352
rect 2136 18164 2188 18216
rect 3516 18232 3568 18284
rect 4252 18232 4304 18284
rect 6368 18275 6420 18284
rect 6368 18241 6377 18275
rect 6377 18241 6411 18275
rect 6411 18241 6420 18275
rect 6368 18232 6420 18241
rect 9220 18368 9272 18420
rect 11060 18368 11112 18420
rect 11704 18368 11756 18420
rect 11980 18411 12032 18420
rect 11980 18377 11989 18411
rect 11989 18377 12023 18411
rect 12023 18377 12032 18411
rect 11980 18368 12032 18377
rect 14372 18368 14424 18420
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 18420 18368 18472 18420
rect 18788 18411 18840 18420
rect 18788 18377 18797 18411
rect 18797 18377 18831 18411
rect 18831 18377 18840 18411
rect 18788 18368 18840 18377
rect 19064 18368 19116 18420
rect 8852 18300 8904 18352
rect 10692 18300 10744 18352
rect 15752 18343 15804 18352
rect 15752 18309 15770 18343
rect 15770 18309 15804 18343
rect 15752 18300 15804 18309
rect 18696 18343 18748 18352
rect 18696 18309 18705 18343
rect 18705 18309 18739 18343
rect 18739 18309 18748 18343
rect 20904 18368 20956 18420
rect 21824 18368 21876 18420
rect 23572 18368 23624 18420
rect 27068 18368 27120 18420
rect 28540 18411 28592 18420
rect 28540 18377 28549 18411
rect 28549 18377 28583 18411
rect 28583 18377 28592 18411
rect 28540 18368 28592 18377
rect 28816 18368 28868 18420
rect 29552 18368 29604 18420
rect 32404 18411 32456 18420
rect 32404 18377 32413 18411
rect 32413 18377 32447 18411
rect 32447 18377 32456 18411
rect 32404 18368 32456 18377
rect 33876 18368 33928 18420
rect 18696 18300 18748 18309
rect 5816 18139 5868 18148
rect 5816 18105 5825 18139
rect 5825 18105 5859 18139
rect 5859 18105 5868 18139
rect 7380 18207 7432 18216
rect 7380 18173 7414 18207
rect 7414 18173 7432 18207
rect 7380 18164 7432 18173
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 5816 18096 5868 18105
rect 7104 18096 7156 18148
rect 5448 18028 5500 18080
rect 7380 18028 7432 18080
rect 9772 18232 9824 18284
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 15936 18232 15988 18284
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 20352 18232 20404 18284
rect 21364 18232 21416 18284
rect 27436 18343 27488 18352
rect 27436 18309 27470 18343
rect 27470 18309 27488 18343
rect 27436 18300 27488 18309
rect 28724 18300 28776 18352
rect 30564 18300 30616 18352
rect 29736 18232 29788 18284
rect 33140 18275 33192 18284
rect 33140 18241 33149 18275
rect 33149 18241 33183 18275
rect 33183 18241 33192 18275
rect 33140 18232 33192 18241
rect 36820 18368 36872 18420
rect 37832 18368 37884 18420
rect 38660 18411 38712 18420
rect 38660 18377 38669 18411
rect 38669 18377 38703 18411
rect 38703 18377 38712 18411
rect 38660 18368 38712 18377
rect 39212 18368 39264 18420
rect 43996 18368 44048 18420
rect 35348 18300 35400 18352
rect 35532 18275 35584 18284
rect 41420 18300 41472 18352
rect 42616 18300 42668 18352
rect 35532 18241 35550 18275
rect 35550 18241 35584 18275
rect 35532 18232 35584 18241
rect 8668 18028 8720 18080
rect 12716 18164 12768 18216
rect 10232 18028 10284 18080
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 12532 18028 12584 18080
rect 13820 18139 13872 18148
rect 13820 18105 13829 18139
rect 13829 18105 13863 18139
rect 13863 18105 13872 18139
rect 13820 18096 13872 18105
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 18328 18164 18380 18216
rect 19892 18164 19944 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 22100 18164 22152 18216
rect 16212 18028 16264 18080
rect 20720 18096 20772 18148
rect 22376 18207 22428 18216
rect 22376 18173 22385 18207
rect 22385 18173 22419 18207
rect 22419 18173 22428 18207
rect 22376 18164 22428 18173
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 25596 18207 25648 18216
rect 25596 18173 25605 18207
rect 25605 18173 25639 18207
rect 25639 18173 25648 18207
rect 25596 18164 25648 18173
rect 25780 18207 25832 18216
rect 25780 18173 25798 18207
rect 25798 18173 25832 18207
rect 25780 18164 25832 18173
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 26148 18207 26200 18216
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 27068 18164 27120 18216
rect 29184 18207 29236 18216
rect 29184 18173 29193 18207
rect 29193 18173 29227 18207
rect 29227 18173 29236 18207
rect 29184 18164 29236 18173
rect 32772 18164 32824 18216
rect 33416 18207 33468 18216
rect 33416 18173 33425 18207
rect 33425 18173 33459 18207
rect 33459 18173 33468 18207
rect 33416 18164 33468 18173
rect 34244 18164 34296 18216
rect 33876 18096 33928 18148
rect 28908 18028 28960 18080
rect 31944 18028 31996 18080
rect 32128 18028 32180 18080
rect 33784 18028 33836 18080
rect 35992 18028 36044 18080
rect 37556 18028 37608 18080
rect 41144 18275 41196 18284
rect 41144 18241 41178 18275
rect 41178 18241 41196 18275
rect 41144 18232 41196 18241
rect 42248 18232 42300 18284
rect 42984 18300 43036 18352
rect 45008 18368 45060 18420
rect 46204 18411 46256 18420
rect 46204 18377 46213 18411
rect 46213 18377 46247 18411
rect 46247 18377 46256 18411
rect 46204 18368 46256 18377
rect 46388 18368 46440 18420
rect 46664 18411 46716 18420
rect 46664 18377 46673 18411
rect 46673 18377 46707 18411
rect 46707 18377 46716 18411
rect 46664 18368 46716 18377
rect 47032 18411 47084 18420
rect 47032 18377 47041 18411
rect 47041 18377 47075 18411
rect 47075 18377 47084 18411
rect 47032 18368 47084 18377
rect 47492 18368 47544 18420
rect 48964 18368 49016 18420
rect 50988 18368 51040 18420
rect 52552 18411 52604 18420
rect 52552 18377 52561 18411
rect 52561 18377 52595 18411
rect 52595 18377 52604 18411
rect 52552 18368 52604 18377
rect 52828 18368 52880 18420
rect 52920 18368 52972 18420
rect 53656 18368 53708 18420
rect 55680 18368 55732 18420
rect 47676 18300 47728 18352
rect 53012 18343 53064 18352
rect 53012 18309 53021 18343
rect 53021 18309 53055 18343
rect 53055 18309 53064 18343
rect 53012 18300 53064 18309
rect 56692 18368 56744 18420
rect 57244 18411 57296 18420
rect 38752 18164 38804 18216
rect 39580 18164 39632 18216
rect 42524 18207 42576 18216
rect 42524 18173 42533 18207
rect 42533 18173 42567 18207
rect 42567 18173 42576 18207
rect 42524 18164 42576 18173
rect 48320 18232 48372 18284
rect 52552 18232 52604 18284
rect 43260 18096 43312 18148
rect 48504 18207 48556 18216
rect 48504 18173 48513 18207
rect 48513 18173 48547 18207
rect 48547 18173 48556 18207
rect 48504 18164 48556 18173
rect 48780 18207 48832 18216
rect 48780 18173 48789 18207
rect 48789 18173 48823 18207
rect 48823 18173 48832 18207
rect 48780 18164 48832 18173
rect 46756 18096 46808 18148
rect 47124 18096 47176 18148
rect 49424 18207 49476 18216
rect 49424 18173 49433 18207
rect 49433 18173 49467 18207
rect 49467 18173 49476 18207
rect 49424 18164 49476 18173
rect 51172 18207 51224 18216
rect 51172 18173 51181 18207
rect 51181 18173 51215 18207
rect 51215 18173 51224 18207
rect 51172 18164 51224 18173
rect 52828 18207 52880 18216
rect 52828 18173 52837 18207
rect 52837 18173 52871 18207
rect 52871 18173 52880 18207
rect 52828 18164 52880 18173
rect 54576 18275 54628 18284
rect 54576 18241 54585 18275
rect 54585 18241 54619 18275
rect 54619 18241 54628 18275
rect 54576 18232 54628 18241
rect 56232 18300 56284 18352
rect 57244 18377 57253 18411
rect 57253 18377 57287 18411
rect 57287 18377 57296 18411
rect 57244 18368 57296 18377
rect 54852 18207 54904 18216
rect 54852 18173 54861 18207
rect 54861 18173 54895 18207
rect 54895 18173 54904 18207
rect 54852 18164 54904 18173
rect 39580 18071 39632 18080
rect 39580 18037 39589 18071
rect 39589 18037 39623 18071
rect 39623 18037 39632 18071
rect 39580 18028 39632 18037
rect 42524 18028 42576 18080
rect 45836 18028 45888 18080
rect 46572 18028 46624 18080
rect 50712 18028 50764 18080
rect 54392 18028 54444 18080
rect 57704 18164 57756 18216
rect 56140 18028 56192 18080
rect 57336 18028 57388 18080
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 22616 17926 22668 17978
rect 22680 17926 22732 17978
rect 22744 17926 22796 17978
rect 22808 17926 22860 17978
rect 22872 17926 22924 17978
rect 37060 17926 37112 17978
rect 37124 17926 37176 17978
rect 37188 17926 37240 17978
rect 37252 17926 37304 17978
rect 37316 17926 37368 17978
rect 51504 17926 51556 17978
rect 51568 17926 51620 17978
rect 51632 17926 51684 17978
rect 51696 17926 51748 17978
rect 51760 17926 51812 17978
rect 4160 17824 4212 17876
rect 6368 17824 6420 17876
rect 8668 17867 8720 17876
rect 8668 17833 8677 17867
rect 8677 17833 8711 17867
rect 8711 17833 8720 17867
rect 8668 17824 8720 17833
rect 9588 17824 9640 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 9772 17867 9824 17876
rect 9772 17833 9781 17867
rect 9781 17833 9815 17867
rect 9815 17833 9824 17867
rect 9772 17824 9824 17833
rect 12440 17824 12492 17876
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 14924 17824 14976 17876
rect 18052 17824 18104 17876
rect 20260 17824 20312 17876
rect 20720 17824 20772 17876
rect 23848 17824 23900 17876
rect 25596 17824 25648 17876
rect 25780 17867 25832 17876
rect 25780 17833 25789 17867
rect 25789 17833 25823 17867
rect 25823 17833 25832 17867
rect 25780 17824 25832 17833
rect 28908 17824 28960 17876
rect 34244 17824 34296 17876
rect 4160 17688 4212 17740
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 4436 17620 4488 17672
rect 5448 17688 5500 17740
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 9680 17688 9732 17740
rect 10232 17688 10284 17740
rect 14464 17688 14516 17740
rect 14740 17688 14792 17740
rect 16212 17731 16264 17740
rect 16212 17697 16221 17731
rect 16221 17697 16255 17731
rect 16255 17697 16264 17731
rect 16212 17688 16264 17697
rect 16948 17731 17000 17740
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 20536 17688 20588 17740
rect 7012 17663 7064 17672
rect 7012 17629 7030 17663
rect 7030 17629 7064 17663
rect 7012 17620 7064 17629
rect 9496 17620 9548 17672
rect 10416 17620 10468 17672
rect 12624 17620 12676 17672
rect 13268 17620 13320 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 20812 17620 20864 17672
rect 23480 17688 23532 17740
rect 35992 17756 36044 17808
rect 37924 17756 37976 17808
rect 27068 17731 27120 17740
rect 22100 17620 22152 17672
rect 27068 17697 27077 17731
rect 27077 17697 27111 17731
rect 27111 17697 27120 17731
rect 27068 17688 27120 17697
rect 29736 17688 29788 17740
rect 25780 17620 25832 17672
rect 28264 17620 28316 17672
rect 33784 17688 33836 17740
rect 34428 17731 34480 17740
rect 34428 17697 34437 17731
rect 34437 17697 34471 17731
rect 34471 17697 34480 17731
rect 34428 17688 34480 17697
rect 37740 17688 37792 17740
rect 38660 17824 38712 17876
rect 45008 17824 45060 17876
rect 46020 17824 46072 17876
rect 42616 17756 42668 17808
rect 37648 17663 37700 17672
rect 37648 17629 37657 17663
rect 37657 17629 37691 17663
rect 37691 17629 37700 17663
rect 37648 17620 37700 17629
rect 38476 17663 38528 17672
rect 38476 17629 38510 17663
rect 38510 17629 38528 17663
rect 38476 17620 38528 17629
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 9220 17527 9272 17536
rect 9220 17493 9229 17527
rect 9229 17493 9263 17527
rect 9263 17493 9272 17527
rect 9220 17484 9272 17493
rect 9680 17484 9732 17536
rect 12532 17552 12584 17604
rect 12992 17552 13044 17604
rect 13452 17552 13504 17604
rect 17408 17552 17460 17604
rect 22192 17552 22244 17604
rect 25044 17552 25096 17604
rect 21272 17484 21324 17536
rect 21732 17527 21784 17536
rect 21732 17493 21741 17527
rect 21741 17493 21775 17527
rect 21775 17493 21784 17527
rect 21732 17484 21784 17493
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 24860 17484 24912 17536
rect 26148 17552 26200 17604
rect 26884 17552 26936 17604
rect 31024 17552 31076 17604
rect 31944 17552 31996 17604
rect 32864 17552 32916 17604
rect 32956 17552 33008 17604
rect 25872 17527 25924 17536
rect 25872 17493 25881 17527
rect 25881 17493 25915 17527
rect 25915 17493 25924 17527
rect 25872 17484 25924 17493
rect 28724 17527 28776 17536
rect 28724 17493 28733 17527
rect 28733 17493 28767 17527
rect 28767 17493 28776 17527
rect 28724 17484 28776 17493
rect 29184 17484 29236 17536
rect 33416 17484 33468 17536
rect 34520 17484 34572 17536
rect 34704 17552 34756 17604
rect 36728 17595 36780 17604
rect 36728 17561 36737 17595
rect 36737 17561 36771 17595
rect 36771 17561 36780 17595
rect 36728 17552 36780 17561
rect 35440 17527 35492 17536
rect 35440 17493 35449 17527
rect 35449 17493 35483 17527
rect 35483 17493 35492 17527
rect 35440 17484 35492 17493
rect 48504 17824 48556 17876
rect 49424 17824 49476 17876
rect 50344 17824 50396 17876
rect 52736 17824 52788 17876
rect 54300 17824 54352 17876
rect 56600 17824 56652 17876
rect 56692 17824 56744 17876
rect 57704 17867 57756 17876
rect 57704 17833 57713 17867
rect 57713 17833 57747 17867
rect 57747 17833 57756 17867
rect 57704 17824 57756 17833
rect 45284 17663 45336 17672
rect 45284 17629 45318 17663
rect 45318 17629 45336 17663
rect 45284 17620 45336 17629
rect 47400 17620 47452 17672
rect 48596 17620 48648 17672
rect 47768 17552 47820 17604
rect 39304 17527 39356 17536
rect 39304 17493 39313 17527
rect 39313 17493 39347 17527
rect 39347 17493 39356 17527
rect 39304 17484 39356 17493
rect 42524 17484 42576 17536
rect 42708 17484 42760 17536
rect 43444 17484 43496 17536
rect 48780 17484 48832 17536
rect 50712 17731 50764 17740
rect 50712 17697 50721 17731
rect 50721 17697 50755 17731
rect 50755 17697 50764 17731
rect 50712 17688 50764 17697
rect 54852 17688 54904 17740
rect 51172 17663 51224 17672
rect 51172 17629 51181 17663
rect 51181 17629 51215 17663
rect 51215 17629 51224 17663
rect 51172 17620 51224 17629
rect 51908 17595 51960 17604
rect 51908 17561 51942 17595
rect 51942 17561 51960 17595
rect 51908 17552 51960 17561
rect 49332 17484 49384 17536
rect 49884 17484 49936 17536
rect 52000 17484 52052 17536
rect 54300 17484 54352 17536
rect 56140 17620 56192 17672
rect 56968 17620 57020 17672
rect 58348 17663 58400 17672
rect 58348 17629 58357 17663
rect 58357 17629 58391 17663
rect 58391 17629 58400 17663
rect 58348 17620 58400 17629
rect 55680 17527 55732 17536
rect 55680 17493 55689 17527
rect 55689 17493 55723 17527
rect 55723 17493 55732 17527
rect 55680 17484 55732 17493
rect 15394 17382 15446 17434
rect 15458 17382 15510 17434
rect 15522 17382 15574 17434
rect 15586 17382 15638 17434
rect 15650 17382 15702 17434
rect 29838 17382 29890 17434
rect 29902 17382 29954 17434
rect 29966 17382 30018 17434
rect 30030 17382 30082 17434
rect 30094 17382 30146 17434
rect 44282 17382 44334 17434
rect 44346 17382 44398 17434
rect 44410 17382 44462 17434
rect 44474 17382 44526 17434
rect 44538 17382 44590 17434
rect 58726 17382 58778 17434
rect 58790 17382 58842 17434
rect 58854 17382 58906 17434
rect 58918 17382 58970 17434
rect 58982 17382 59034 17434
rect 3516 17280 3568 17332
rect 7288 17280 7340 17332
rect 9404 17280 9456 17332
rect 12992 17323 13044 17332
rect 12992 17289 13001 17323
rect 13001 17289 13035 17323
rect 13035 17289 13044 17323
rect 12992 17280 13044 17289
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 19616 17280 19668 17332
rect 21732 17280 21784 17332
rect 22376 17280 22428 17332
rect 25044 17323 25096 17332
rect 25044 17289 25053 17323
rect 25053 17289 25087 17323
rect 25087 17289 25096 17323
rect 25044 17280 25096 17289
rect 25872 17280 25924 17332
rect 26608 17280 26660 17332
rect 28172 17280 28224 17332
rect 31024 17323 31076 17332
rect 31024 17289 31033 17323
rect 31033 17289 31067 17323
rect 31067 17289 31076 17323
rect 31024 17280 31076 17289
rect 32036 17280 32088 17332
rect 32864 17323 32916 17332
rect 32864 17289 32873 17323
rect 32873 17289 32907 17323
rect 32907 17289 32916 17323
rect 32864 17280 32916 17289
rect 37740 17280 37792 17332
rect 38844 17280 38896 17332
rect 39304 17280 39356 17332
rect 43720 17323 43772 17332
rect 43720 17289 43729 17323
rect 43729 17289 43763 17323
rect 43763 17289 43772 17323
rect 43720 17280 43772 17289
rect 47400 17280 47452 17332
rect 47768 17323 47820 17332
rect 47768 17289 47777 17323
rect 47777 17289 47811 17323
rect 47811 17289 47820 17323
rect 47768 17280 47820 17289
rect 48872 17280 48924 17332
rect 57336 17280 57388 17332
rect 58348 17280 58400 17332
rect 3976 17212 4028 17264
rect 9128 17212 9180 17264
rect 19892 17212 19944 17264
rect 8300 17144 8352 17196
rect 9772 17144 9824 17196
rect 13176 17144 13228 17196
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 25504 17144 25556 17196
rect 31576 17187 31628 17196
rect 31576 17153 31585 17187
rect 31585 17153 31619 17187
rect 31619 17153 31628 17187
rect 31576 17144 31628 17153
rect 33416 17144 33468 17196
rect 33600 17144 33652 17196
rect 39580 17212 39632 17264
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 2596 16983 2648 16992
rect 2596 16949 2605 16983
rect 2605 16949 2639 16983
rect 2639 16949 2648 16983
rect 2596 16940 2648 16949
rect 4620 17076 4672 17128
rect 5264 17076 5316 17128
rect 8668 17076 8720 17128
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 9220 17008 9272 17060
rect 9956 17008 10008 17060
rect 24768 17076 24820 17128
rect 25136 17076 25188 17128
rect 48412 17187 48464 17196
rect 48412 17153 48421 17187
rect 48421 17153 48455 17187
rect 48455 17153 48464 17187
rect 48412 17144 48464 17153
rect 49424 17144 49476 17196
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 6000 16940 6052 16992
rect 6276 16940 6328 16992
rect 7104 16940 7156 16992
rect 7932 16940 7984 16992
rect 12716 16940 12768 16992
rect 12992 16940 13044 16992
rect 17592 16940 17644 16992
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 19708 16940 19760 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 34520 16940 34572 16992
rect 35348 16940 35400 16992
rect 38844 16940 38896 16992
rect 42984 17119 43036 17128
rect 42984 17085 42993 17119
rect 42993 17085 43027 17119
rect 43027 17085 43036 17119
rect 42984 17076 43036 17085
rect 43444 17119 43496 17128
rect 43444 17085 43453 17119
rect 43453 17085 43487 17119
rect 43487 17085 43496 17119
rect 43444 17076 43496 17085
rect 43628 17119 43680 17128
rect 43628 17085 43637 17119
rect 43637 17085 43671 17119
rect 43671 17085 43680 17119
rect 43628 17076 43680 17085
rect 44272 17119 44324 17128
rect 44272 17085 44281 17119
rect 44281 17085 44315 17119
rect 44315 17085 44324 17119
rect 44272 17076 44324 17085
rect 45652 17076 45704 17128
rect 56876 17119 56928 17128
rect 56876 17085 56885 17119
rect 56885 17085 56919 17119
rect 56919 17085 56928 17119
rect 56876 17076 56928 17085
rect 43996 17008 44048 17060
rect 55680 17008 55732 17060
rect 57704 17076 57756 17128
rect 58256 17008 58308 17060
rect 39304 16983 39356 16992
rect 39304 16949 39313 16983
rect 39313 16949 39347 16983
rect 39347 16949 39356 16983
rect 39304 16940 39356 16949
rect 39856 16940 39908 16992
rect 41604 16983 41656 16992
rect 41604 16949 41613 16983
rect 41613 16949 41647 16983
rect 41647 16949 41656 16983
rect 41604 16940 41656 16949
rect 42340 16940 42392 16992
rect 42432 16983 42484 16992
rect 42432 16949 42441 16983
rect 42441 16949 42475 16983
rect 42475 16949 42484 16983
rect 42432 16940 42484 16949
rect 44088 16983 44140 16992
rect 44088 16949 44097 16983
rect 44097 16949 44131 16983
rect 44131 16949 44140 16983
rect 44088 16940 44140 16949
rect 44824 16983 44876 16992
rect 44824 16949 44833 16983
rect 44833 16949 44867 16983
rect 44867 16949 44876 16983
rect 44824 16940 44876 16949
rect 53196 16983 53248 16992
rect 53196 16949 53205 16983
rect 53205 16949 53239 16983
rect 53239 16949 53248 16983
rect 53196 16940 53248 16949
rect 56140 16983 56192 16992
rect 56140 16949 56149 16983
rect 56149 16949 56183 16983
rect 56183 16949 56192 16983
rect 56140 16940 56192 16949
rect 57888 16983 57940 16992
rect 57888 16949 57897 16983
rect 57897 16949 57931 16983
rect 57931 16949 57940 16983
rect 57888 16940 57940 16949
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 22616 16838 22668 16890
rect 22680 16838 22732 16890
rect 22744 16838 22796 16890
rect 22808 16838 22860 16890
rect 22872 16838 22924 16890
rect 37060 16838 37112 16890
rect 37124 16838 37176 16890
rect 37188 16838 37240 16890
rect 37252 16838 37304 16890
rect 37316 16838 37368 16890
rect 51504 16838 51556 16890
rect 51568 16838 51620 16890
rect 51632 16838 51684 16890
rect 51696 16838 51748 16890
rect 51760 16838 51812 16890
rect 6368 16736 6420 16788
rect 6276 16668 6328 16720
rect 2136 16532 2188 16584
rect 2964 16532 3016 16584
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 9404 16600 9456 16652
rect 23756 16736 23808 16788
rect 26608 16736 26660 16788
rect 31944 16736 31996 16788
rect 32864 16736 32916 16788
rect 34520 16736 34572 16788
rect 38292 16736 38344 16788
rect 39856 16736 39908 16788
rect 9680 16668 9732 16720
rect 12164 16668 12216 16720
rect 12900 16668 12952 16720
rect 17592 16668 17644 16720
rect 23388 16668 23440 16720
rect 32404 16668 32456 16720
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 25596 16643 25648 16652
rect 25596 16609 25605 16643
rect 25605 16609 25639 16643
rect 25639 16609 25648 16643
rect 25596 16600 25648 16609
rect 26240 16600 26292 16652
rect 4620 16464 4672 16516
rect 7288 16532 7340 16584
rect 7932 16532 7984 16584
rect 7472 16464 7524 16516
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 5448 16396 5500 16448
rect 8760 16532 8812 16584
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 13820 16575 13872 16584
rect 13820 16541 13829 16575
rect 13829 16541 13863 16575
rect 13863 16541 13872 16575
rect 13820 16532 13872 16541
rect 13912 16532 13964 16584
rect 15200 16532 15252 16584
rect 18052 16532 18104 16584
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 24308 16532 24360 16584
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 30840 16575 30892 16584
rect 30840 16541 30849 16575
rect 30849 16541 30883 16575
rect 30883 16541 30892 16575
rect 30840 16532 30892 16541
rect 35624 16600 35676 16652
rect 37832 16643 37884 16652
rect 37832 16609 37841 16643
rect 37841 16609 37875 16643
rect 37875 16609 37884 16643
rect 37832 16600 37884 16609
rect 38476 16600 38528 16652
rect 33508 16532 33560 16584
rect 35256 16575 35308 16584
rect 35256 16541 35265 16575
rect 35265 16541 35299 16575
rect 35299 16541 35308 16575
rect 35256 16532 35308 16541
rect 36820 16532 36872 16584
rect 37924 16575 37976 16584
rect 37924 16541 37933 16575
rect 37933 16541 37967 16575
rect 37967 16541 37976 16575
rect 37924 16532 37976 16541
rect 38844 16532 38896 16584
rect 42432 16736 42484 16788
rect 42340 16643 42392 16652
rect 42340 16609 42349 16643
rect 42349 16609 42383 16643
rect 42383 16609 42392 16643
rect 42340 16600 42392 16609
rect 45560 16736 45612 16788
rect 49700 16736 49752 16788
rect 44272 16711 44324 16720
rect 44272 16677 44281 16711
rect 44281 16677 44315 16711
rect 44315 16677 44324 16711
rect 44272 16668 44324 16677
rect 44640 16668 44692 16720
rect 50528 16668 50580 16720
rect 45100 16600 45152 16652
rect 48780 16600 48832 16652
rect 49424 16600 49476 16652
rect 54576 16600 54628 16652
rect 57060 16600 57112 16652
rect 42984 16532 43036 16584
rect 43996 16532 44048 16584
rect 44824 16532 44876 16584
rect 45652 16532 45704 16584
rect 47768 16575 47820 16584
rect 47768 16541 47777 16575
rect 47777 16541 47811 16575
rect 47811 16541 47820 16575
rect 47768 16532 47820 16541
rect 49148 16575 49200 16584
rect 49148 16541 49157 16575
rect 49157 16541 49191 16575
rect 49191 16541 49200 16575
rect 49148 16532 49200 16541
rect 49976 16532 50028 16584
rect 53840 16575 53892 16584
rect 53840 16541 53849 16575
rect 53849 16541 53883 16575
rect 53883 16541 53892 16575
rect 53840 16532 53892 16541
rect 57888 16532 57940 16584
rect 34244 16507 34296 16516
rect 34244 16473 34253 16507
rect 34253 16473 34287 16507
rect 34287 16473 34296 16507
rect 34244 16464 34296 16473
rect 8116 16396 8168 16448
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13268 16439 13320 16448
rect 13268 16405 13277 16439
rect 13277 16405 13311 16439
rect 13311 16405 13320 16439
rect 13268 16396 13320 16405
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 16856 16396 16908 16448
rect 17776 16439 17828 16448
rect 17776 16405 17785 16439
rect 17785 16405 17819 16439
rect 17819 16405 17828 16439
rect 17776 16396 17828 16405
rect 20720 16396 20772 16448
rect 24216 16439 24268 16448
rect 24216 16405 24225 16439
rect 24225 16405 24259 16439
rect 24259 16405 24268 16439
rect 24216 16396 24268 16405
rect 24400 16439 24452 16448
rect 24400 16405 24409 16439
rect 24409 16405 24443 16439
rect 24443 16405 24452 16439
rect 24400 16396 24452 16405
rect 25596 16396 25648 16448
rect 30288 16439 30340 16448
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 31208 16439 31260 16448
rect 31208 16405 31217 16439
rect 31217 16405 31251 16439
rect 31251 16405 31260 16439
rect 31208 16396 31260 16405
rect 34704 16439 34756 16448
rect 34704 16405 34713 16439
rect 34713 16405 34747 16439
rect 34747 16405 34756 16439
rect 34704 16396 34756 16405
rect 35440 16439 35492 16448
rect 35440 16405 35449 16439
rect 35449 16405 35483 16439
rect 35483 16405 35492 16439
rect 35440 16396 35492 16405
rect 36452 16439 36504 16448
rect 36452 16405 36461 16439
rect 36461 16405 36495 16439
rect 36495 16405 36504 16439
rect 36452 16396 36504 16405
rect 36912 16396 36964 16448
rect 38568 16439 38620 16448
rect 38568 16405 38577 16439
rect 38577 16405 38611 16439
rect 38611 16405 38620 16439
rect 38568 16396 38620 16405
rect 41236 16464 41288 16516
rect 41788 16439 41840 16448
rect 41788 16405 41797 16439
rect 41797 16405 41831 16439
rect 41831 16405 41840 16439
rect 41788 16396 41840 16405
rect 42248 16396 42300 16448
rect 43352 16464 43404 16516
rect 44180 16396 44232 16448
rect 45744 16464 45796 16516
rect 55772 16464 55824 16516
rect 45376 16396 45428 16448
rect 48228 16396 48280 16448
rect 48596 16439 48648 16448
rect 48596 16405 48605 16439
rect 48605 16405 48639 16439
rect 48639 16405 48648 16439
rect 48596 16396 48648 16405
rect 50160 16439 50212 16448
rect 50160 16405 50169 16439
rect 50169 16405 50203 16439
rect 50203 16405 50212 16439
rect 50160 16396 50212 16405
rect 53104 16396 53156 16448
rect 56784 16396 56836 16448
rect 57428 16439 57480 16448
rect 57428 16405 57437 16439
rect 57437 16405 57471 16439
rect 57471 16405 57480 16439
rect 57428 16396 57480 16405
rect 15394 16294 15446 16346
rect 15458 16294 15510 16346
rect 15522 16294 15574 16346
rect 15586 16294 15638 16346
rect 15650 16294 15702 16346
rect 29838 16294 29890 16346
rect 29902 16294 29954 16346
rect 29966 16294 30018 16346
rect 30030 16294 30082 16346
rect 30094 16294 30146 16346
rect 44282 16294 44334 16346
rect 44346 16294 44398 16346
rect 44410 16294 44462 16346
rect 44474 16294 44526 16346
rect 44538 16294 44590 16346
rect 58726 16294 58778 16346
rect 58790 16294 58842 16346
rect 58854 16294 58906 16346
rect 58918 16294 58970 16346
rect 58982 16294 59034 16346
rect 3240 16192 3292 16244
rect 3792 16192 3844 16244
rect 3976 16235 4028 16244
rect 3976 16201 3985 16235
rect 3985 16201 4019 16235
rect 4019 16201 4028 16235
rect 3976 16192 4028 16201
rect 6276 16192 6328 16244
rect 2596 16124 2648 16176
rect 7472 16192 7524 16244
rect 2136 16056 2188 16108
rect 7288 16056 7340 16108
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 11704 16192 11756 16244
rect 13268 16192 13320 16244
rect 13912 16192 13964 16244
rect 14832 16192 14884 16244
rect 17776 16192 17828 16244
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 20628 16192 20680 16244
rect 20812 16192 20864 16244
rect 24216 16192 24268 16244
rect 24860 16235 24912 16244
rect 24860 16201 24869 16235
rect 24869 16201 24903 16235
rect 24903 16201 24912 16235
rect 24860 16192 24912 16201
rect 26332 16192 26384 16244
rect 30840 16192 30892 16244
rect 34520 16192 34572 16244
rect 35256 16192 35308 16244
rect 35440 16192 35492 16244
rect 36452 16192 36504 16244
rect 37832 16192 37884 16244
rect 38568 16192 38620 16244
rect 41236 16235 41288 16244
rect 41236 16201 41245 16235
rect 41245 16201 41279 16235
rect 41279 16201 41288 16235
rect 41236 16192 41288 16201
rect 41788 16192 41840 16244
rect 43628 16192 43680 16244
rect 47768 16192 47820 16244
rect 48596 16192 48648 16244
rect 10784 16056 10836 16108
rect 11612 16056 11664 16108
rect 11888 16056 11940 16108
rect 19892 16056 19944 16108
rect 21088 16056 21140 16108
rect 34244 16124 34296 16176
rect 4344 15920 4396 15972
rect 6736 16031 6788 16040
rect 6736 15997 6745 16031
rect 6745 15997 6779 16031
rect 6779 15997 6788 16031
rect 6736 15988 6788 15997
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 11796 15988 11848 16040
rect 12164 16031 12216 16040
rect 12164 15997 12173 16031
rect 12173 15997 12207 16031
rect 12207 15997 12216 16031
rect 12164 15988 12216 15997
rect 12716 15988 12768 16040
rect 14648 15988 14700 16040
rect 16488 15988 16540 16040
rect 20168 15988 20220 16040
rect 24676 16056 24728 16108
rect 25780 16056 25832 16108
rect 30840 16099 30892 16108
rect 30840 16065 30849 16099
rect 30849 16065 30883 16099
rect 30883 16065 30892 16099
rect 30840 16056 30892 16065
rect 35348 16099 35400 16108
rect 35348 16065 35357 16099
rect 35357 16065 35391 16099
rect 35391 16065 35400 16099
rect 35348 16056 35400 16065
rect 38844 16056 38896 16108
rect 43352 16099 43404 16108
rect 43352 16065 43361 16099
rect 43361 16065 43395 16099
rect 43395 16065 43404 16099
rect 43352 16056 43404 16065
rect 44640 16056 44692 16108
rect 19064 15920 19116 15972
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11520 15852 11572 15904
rect 12900 15852 12952 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 18328 15895 18380 15904
rect 18328 15861 18337 15895
rect 18337 15861 18371 15895
rect 18371 15861 18380 15895
rect 18328 15852 18380 15861
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 22008 15920 22060 15972
rect 23756 15988 23808 16040
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 25504 15988 25556 15997
rect 26608 15988 26660 16040
rect 27528 16031 27580 16040
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 28356 16031 28408 16040
rect 28356 15997 28365 16031
rect 28365 15997 28399 16031
rect 28399 15997 28408 16031
rect 28356 15988 28408 15997
rect 31024 16031 31076 16040
rect 31024 15997 31033 16031
rect 31033 15997 31067 16031
rect 31067 15997 31076 16031
rect 31024 15988 31076 15997
rect 31852 16031 31904 16040
rect 31852 15997 31861 16031
rect 31861 15997 31895 16031
rect 31895 15997 31904 16031
rect 31852 15988 31904 15997
rect 24308 15920 24360 15972
rect 41328 15988 41380 16040
rect 42892 15988 42944 16040
rect 43076 16031 43128 16040
rect 43076 15997 43085 16031
rect 43085 15997 43119 16031
rect 43119 15997 43128 16031
rect 43076 15988 43128 15997
rect 43260 16031 43312 16040
rect 43260 15997 43278 16031
rect 43278 15997 43312 16031
rect 43260 15988 43312 15997
rect 43536 15988 43588 16040
rect 44732 15988 44784 16040
rect 22100 15852 22152 15904
rect 23388 15852 23440 15904
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 24952 15895 25004 15904
rect 24952 15861 24961 15895
rect 24961 15861 24995 15895
rect 24995 15861 25004 15895
rect 24952 15852 25004 15861
rect 26608 15852 26660 15904
rect 27804 15895 27856 15904
rect 27804 15861 27813 15895
rect 27813 15861 27847 15895
rect 27847 15861 27856 15895
rect 27804 15852 27856 15861
rect 32864 15852 32916 15904
rect 37648 15852 37700 15904
rect 42616 15920 42668 15972
rect 47584 16056 47636 16108
rect 48044 16056 48096 16108
rect 52000 16192 52052 16244
rect 53196 16192 53248 16244
rect 53840 16192 53892 16244
rect 55772 16235 55824 16244
rect 55772 16201 55781 16235
rect 55781 16201 55815 16235
rect 55815 16201 55824 16235
rect 55772 16192 55824 16201
rect 57428 16192 57480 16244
rect 57704 16235 57756 16244
rect 57704 16201 57713 16235
rect 57713 16201 57747 16235
rect 57747 16201 57756 16235
rect 57704 16192 57756 16201
rect 50160 16124 50212 16176
rect 47124 15988 47176 16040
rect 38752 15895 38804 15904
rect 38752 15861 38761 15895
rect 38761 15861 38795 15895
rect 38795 15861 38804 15895
rect 38752 15852 38804 15861
rect 41052 15895 41104 15904
rect 41052 15861 41061 15895
rect 41061 15861 41095 15895
rect 41095 15861 41104 15895
rect 41052 15852 41104 15861
rect 42064 15852 42116 15904
rect 43536 15852 43588 15904
rect 57152 16056 57204 16108
rect 49056 16031 49108 16040
rect 49056 15997 49065 16031
rect 49065 15997 49099 16031
rect 49099 15997 49108 16031
rect 49056 15988 49108 15997
rect 53748 16031 53800 16040
rect 53748 15997 53757 16031
rect 53757 15997 53791 16031
rect 53791 15997 53800 16031
rect 53748 15988 53800 15997
rect 54668 16031 54720 16040
rect 54668 15997 54677 16031
rect 54677 15997 54711 16031
rect 54711 15997 54720 16031
rect 54668 15988 54720 15997
rect 56048 15920 56100 15972
rect 44364 15895 44416 15904
rect 44364 15861 44373 15895
rect 44373 15861 44407 15895
rect 44407 15861 44416 15895
rect 44364 15852 44416 15861
rect 45100 15852 45152 15904
rect 46848 15852 46900 15904
rect 47124 15852 47176 15904
rect 48412 15895 48464 15904
rect 48412 15861 48421 15895
rect 48421 15861 48455 15895
rect 48455 15861 48464 15895
rect 48412 15852 48464 15861
rect 49056 15852 49108 15904
rect 49516 15852 49568 15904
rect 50620 15895 50672 15904
rect 50620 15861 50629 15895
rect 50629 15861 50663 15895
rect 50663 15861 50672 15895
rect 50620 15852 50672 15861
rect 50712 15895 50764 15904
rect 50712 15861 50721 15895
rect 50721 15861 50755 15895
rect 50755 15861 50764 15895
rect 50712 15852 50764 15861
rect 52552 15895 52604 15904
rect 52552 15861 52561 15895
rect 52561 15861 52595 15895
rect 52595 15861 52604 15895
rect 52552 15852 52604 15861
rect 54116 15895 54168 15904
rect 54116 15861 54125 15895
rect 54125 15861 54159 15895
rect 54159 15861 54168 15895
rect 54116 15852 54168 15861
rect 54208 15852 54260 15904
rect 56140 15895 56192 15904
rect 56140 15861 56149 15895
rect 56149 15861 56183 15895
rect 56183 15861 56192 15895
rect 56140 15852 56192 15861
rect 57888 15895 57940 15904
rect 57888 15861 57897 15895
rect 57897 15861 57931 15895
rect 57931 15861 57940 15895
rect 57888 15852 57940 15861
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 22616 15750 22668 15802
rect 22680 15750 22732 15802
rect 22744 15750 22796 15802
rect 22808 15750 22860 15802
rect 22872 15750 22924 15802
rect 37060 15750 37112 15802
rect 37124 15750 37176 15802
rect 37188 15750 37240 15802
rect 37252 15750 37304 15802
rect 37316 15750 37368 15802
rect 51504 15750 51556 15802
rect 51568 15750 51620 15802
rect 51632 15750 51684 15802
rect 51696 15750 51748 15802
rect 51760 15750 51812 15802
rect 6736 15648 6788 15700
rect 8944 15648 8996 15700
rect 9864 15648 9916 15700
rect 11520 15691 11572 15700
rect 11520 15657 11529 15691
rect 11529 15657 11563 15691
rect 11563 15657 11572 15691
rect 11520 15648 11572 15657
rect 8852 15580 8904 15632
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 4344 15487 4396 15496
rect 4344 15453 4353 15487
rect 4353 15453 4387 15487
rect 4387 15453 4396 15487
rect 4344 15444 4396 15453
rect 6184 15444 6236 15496
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 12900 15512 12952 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13176 15512 13228 15564
rect 13636 15512 13688 15564
rect 15200 15648 15252 15700
rect 15568 15648 15620 15700
rect 18052 15691 18104 15700
rect 18052 15657 18061 15691
rect 18061 15657 18095 15691
rect 18095 15657 18104 15691
rect 18052 15648 18104 15657
rect 18328 15648 18380 15700
rect 21364 15648 21416 15700
rect 24308 15648 24360 15700
rect 25044 15648 25096 15700
rect 25504 15648 25556 15700
rect 13820 15512 13872 15564
rect 19064 15580 19116 15632
rect 20628 15580 20680 15632
rect 9864 15444 9916 15496
rect 10232 15444 10284 15496
rect 10692 15444 10744 15496
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 18880 15512 18932 15564
rect 20168 15555 20220 15564
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 22100 15512 22152 15564
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 6460 15376 6512 15428
rect 11796 15376 11848 15428
rect 2688 15351 2740 15360
rect 2688 15317 2697 15351
rect 2697 15317 2731 15351
rect 2731 15317 2740 15351
rect 2688 15308 2740 15317
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 5264 15351 5316 15360
rect 5264 15317 5273 15351
rect 5273 15317 5307 15351
rect 5307 15317 5316 15351
rect 5264 15308 5316 15317
rect 5724 15308 5776 15360
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 7932 15308 7984 15360
rect 9588 15308 9640 15360
rect 11980 15351 12032 15360
rect 11980 15317 11989 15351
rect 11989 15317 12023 15351
rect 12023 15317 12032 15351
rect 11980 15308 12032 15317
rect 13360 15308 13412 15360
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 16488 15444 16540 15496
rect 16856 15487 16908 15496
rect 16856 15453 16890 15487
rect 16890 15453 16908 15487
rect 16856 15444 16908 15453
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 15752 15308 15804 15317
rect 18420 15351 18472 15360
rect 18420 15317 18429 15351
rect 18429 15317 18463 15351
rect 18463 15317 18472 15351
rect 18420 15308 18472 15317
rect 19616 15308 19668 15360
rect 19800 15308 19852 15360
rect 21456 15444 21508 15496
rect 23480 15444 23532 15496
rect 25964 15512 26016 15564
rect 26332 15555 26384 15564
rect 26332 15521 26341 15555
rect 26341 15521 26375 15555
rect 26375 15521 26384 15555
rect 26332 15512 26384 15521
rect 26884 15623 26936 15632
rect 26884 15589 26893 15623
rect 26893 15589 26927 15623
rect 26927 15589 26936 15623
rect 26884 15580 26936 15589
rect 28356 15648 28408 15700
rect 31760 15580 31812 15632
rect 31852 15580 31904 15632
rect 32956 15555 33008 15564
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 27528 15487 27580 15496
rect 27528 15453 27537 15487
rect 27537 15453 27571 15487
rect 27571 15453 27580 15487
rect 27528 15444 27580 15453
rect 24952 15376 25004 15428
rect 20996 15308 21048 15360
rect 26608 15308 26660 15360
rect 26700 15308 26752 15360
rect 29184 15376 29236 15428
rect 30564 15444 30616 15496
rect 31208 15444 31260 15496
rect 32956 15521 32965 15555
rect 32965 15521 32999 15555
rect 32999 15521 33008 15555
rect 32956 15512 33008 15521
rect 36820 15691 36872 15700
rect 36820 15657 36829 15691
rect 36829 15657 36863 15691
rect 36863 15657 36872 15691
rect 36820 15648 36872 15657
rect 37924 15648 37976 15700
rect 38752 15648 38804 15700
rect 38844 15648 38896 15700
rect 33508 15623 33560 15632
rect 33508 15589 33517 15623
rect 33517 15589 33551 15623
rect 33551 15589 33560 15623
rect 33508 15580 33560 15589
rect 34520 15512 34572 15564
rect 35164 15512 35216 15564
rect 32220 15444 32272 15496
rect 33140 15487 33192 15496
rect 33140 15453 33158 15487
rect 33158 15453 33192 15487
rect 33140 15444 33192 15453
rect 34336 15444 34388 15496
rect 38660 15580 38712 15632
rect 36912 15512 36964 15564
rect 31300 15376 31352 15428
rect 29736 15308 29788 15360
rect 30840 15308 30892 15360
rect 31944 15308 31996 15360
rect 32036 15351 32088 15360
rect 32036 15317 32045 15351
rect 32045 15317 32079 15351
rect 32079 15317 32088 15351
rect 32036 15308 32088 15317
rect 34796 15376 34848 15428
rect 37464 15512 37516 15564
rect 42616 15648 42668 15700
rect 43444 15648 43496 15700
rect 42156 15512 42208 15564
rect 43260 15580 43312 15632
rect 43536 15555 43588 15564
rect 43536 15521 43545 15555
rect 43545 15521 43579 15555
rect 43579 15521 43588 15555
rect 43536 15512 43588 15521
rect 44364 15648 44416 15700
rect 49148 15648 49200 15700
rect 49608 15648 49660 15700
rect 49976 15691 50028 15700
rect 49976 15657 49985 15691
rect 49985 15657 50019 15691
rect 50019 15657 50028 15691
rect 49976 15648 50028 15657
rect 54208 15691 54260 15700
rect 54208 15657 54217 15691
rect 54217 15657 54251 15691
rect 54251 15657 54260 15691
rect 54208 15648 54260 15657
rect 54668 15648 54720 15700
rect 42248 15487 42300 15496
rect 42248 15453 42257 15487
rect 42257 15453 42291 15487
rect 42291 15453 42300 15487
rect 42248 15444 42300 15453
rect 45376 15444 45428 15496
rect 45560 15444 45612 15496
rect 46296 15444 46348 15496
rect 46848 15444 46900 15496
rect 48228 15444 48280 15496
rect 49700 15444 49752 15496
rect 50712 15444 50764 15496
rect 41236 15376 41288 15428
rect 43076 15376 43128 15428
rect 45744 15376 45796 15428
rect 46756 15376 46808 15428
rect 48044 15376 48096 15428
rect 34888 15308 34940 15360
rect 34980 15351 35032 15360
rect 34980 15317 34989 15351
rect 34989 15317 35023 15351
rect 35023 15317 35032 15351
rect 34980 15308 35032 15317
rect 35072 15351 35124 15360
rect 35072 15317 35081 15351
rect 35081 15317 35115 15351
rect 35115 15317 35124 15351
rect 35072 15308 35124 15317
rect 35532 15351 35584 15360
rect 35532 15317 35541 15351
rect 35541 15317 35575 15351
rect 35575 15317 35584 15351
rect 35532 15308 35584 15317
rect 36544 15308 36596 15360
rect 37556 15308 37608 15360
rect 38660 15308 38712 15360
rect 41788 15351 41840 15360
rect 41788 15317 41797 15351
rect 41797 15317 41831 15351
rect 41831 15317 41840 15351
rect 41788 15308 41840 15317
rect 44640 15308 44692 15360
rect 46204 15308 46256 15360
rect 49056 15308 49108 15360
rect 50436 15308 50488 15360
rect 54852 15555 54904 15564
rect 54852 15521 54861 15555
rect 54861 15521 54895 15555
rect 54895 15521 54904 15555
rect 54852 15512 54904 15521
rect 57244 15648 57296 15700
rect 57704 15648 57756 15700
rect 57888 15648 57940 15700
rect 56784 15580 56836 15632
rect 55772 15512 55824 15564
rect 56048 15512 56100 15564
rect 56508 15555 56560 15564
rect 56508 15521 56517 15555
rect 56517 15521 56551 15555
rect 56551 15521 56560 15555
rect 56508 15512 56560 15521
rect 56600 15512 56652 15564
rect 57152 15555 57204 15564
rect 57152 15521 57161 15555
rect 57161 15521 57195 15555
rect 57195 15521 57204 15555
rect 57152 15512 57204 15521
rect 57244 15512 57296 15564
rect 53104 15419 53156 15428
rect 53104 15385 53138 15419
rect 53138 15385 53156 15419
rect 53104 15376 53156 15385
rect 53196 15376 53248 15428
rect 53748 15376 53800 15428
rect 56232 15487 56284 15496
rect 56232 15453 56241 15487
rect 56241 15453 56275 15487
rect 56275 15453 56284 15487
rect 56232 15444 56284 15453
rect 54484 15308 54536 15360
rect 54760 15351 54812 15360
rect 54760 15317 54769 15351
rect 54769 15317 54803 15351
rect 54803 15317 54812 15351
rect 54760 15308 54812 15317
rect 56324 15308 56376 15360
rect 56784 15308 56836 15360
rect 57980 15351 58032 15360
rect 57980 15317 57989 15351
rect 57989 15317 58023 15351
rect 58023 15317 58032 15351
rect 57980 15308 58032 15317
rect 15394 15206 15446 15258
rect 15458 15206 15510 15258
rect 15522 15206 15574 15258
rect 15586 15206 15638 15258
rect 15650 15206 15702 15258
rect 29838 15206 29890 15258
rect 29902 15206 29954 15258
rect 29966 15206 30018 15258
rect 30030 15206 30082 15258
rect 30094 15206 30146 15258
rect 44282 15206 44334 15258
rect 44346 15206 44398 15258
rect 44410 15206 44462 15258
rect 44474 15206 44526 15258
rect 44538 15206 44590 15258
rect 58726 15206 58778 15258
rect 58790 15206 58842 15258
rect 58854 15206 58906 15258
rect 58918 15206 58970 15258
rect 58982 15206 59034 15258
rect 3240 15104 3292 15156
rect 3792 15104 3844 15156
rect 3976 15104 4028 15156
rect 6092 15104 6144 15156
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 6368 15104 6420 15156
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 7748 15104 7800 15156
rect 10048 15104 10100 15156
rect 11336 15104 11388 15156
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 11980 15104 12032 15156
rect 12716 15104 12768 15156
rect 13820 15104 13872 15156
rect 10876 15036 10928 15088
rect 11060 15036 11112 15088
rect 12256 15036 12308 15088
rect 14740 15036 14792 15088
rect 17684 15104 17736 15156
rect 18696 15104 18748 15156
rect 18788 15104 18840 15156
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 4160 14900 4212 14952
rect 4712 14900 4764 14952
rect 5356 14832 5408 14884
rect 5724 14900 5776 14952
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13084 14968 13136 15020
rect 13728 14968 13780 15020
rect 18880 14968 18932 15020
rect 21088 15104 21140 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 23756 15104 23808 15156
rect 24584 15104 24636 15156
rect 25504 15104 25556 15156
rect 25780 15104 25832 15156
rect 20720 15036 20772 15088
rect 24400 15036 24452 15088
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 22468 14968 22520 15020
rect 6552 14900 6604 14952
rect 8576 14943 8628 14952
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 9864 14900 9916 14952
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 3516 14764 3568 14816
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 7104 14807 7156 14816
rect 7104 14773 7113 14807
rect 7113 14773 7147 14807
rect 7147 14773 7156 14807
rect 7104 14764 7156 14773
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 11704 14900 11756 14952
rect 12256 14900 12308 14952
rect 12348 14832 12400 14884
rect 15752 14900 15804 14952
rect 17132 14832 17184 14884
rect 18420 14900 18472 14952
rect 19156 14900 19208 14952
rect 19800 14900 19852 14952
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 23940 14764 23992 14816
rect 25596 15011 25648 15020
rect 25596 14977 25630 15011
rect 25630 14977 25648 15011
rect 25596 14968 25648 14977
rect 26056 14968 26108 15020
rect 26700 15147 26752 15156
rect 26700 15113 26709 15147
rect 26709 15113 26743 15147
rect 26743 15113 26752 15147
rect 26700 15104 26752 15113
rect 27804 15104 27856 15156
rect 29184 15147 29236 15156
rect 29184 15113 29193 15147
rect 29193 15113 29227 15147
rect 29227 15113 29236 15147
rect 29184 15104 29236 15113
rect 31300 15147 31352 15156
rect 31300 15113 31309 15147
rect 31309 15113 31343 15147
rect 31343 15113 31352 15147
rect 31300 15104 31352 15113
rect 31944 15104 31996 15156
rect 34704 15104 34756 15156
rect 34980 15104 35032 15156
rect 36728 15104 36780 15156
rect 38016 15104 38068 15156
rect 41236 15147 41288 15156
rect 41236 15113 41245 15147
rect 41245 15113 41279 15147
rect 41279 15113 41288 15147
rect 41236 15104 41288 15113
rect 43536 15104 43588 15156
rect 30288 15036 30340 15088
rect 35532 15036 35584 15088
rect 27896 14968 27948 15020
rect 32036 14968 32088 15020
rect 26700 14764 26752 14816
rect 29736 14900 29788 14952
rect 31760 14900 31812 14952
rect 33048 14968 33100 15020
rect 37464 15011 37516 15020
rect 32864 14900 32916 14952
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 31852 14832 31904 14884
rect 35072 14900 35124 14952
rect 35624 14900 35676 14952
rect 34888 14832 34940 14884
rect 34336 14807 34388 14816
rect 34336 14773 34345 14807
rect 34345 14773 34379 14807
rect 34379 14773 34388 14807
rect 38200 14900 38252 14952
rect 39764 14875 39816 14884
rect 39764 14841 39773 14875
rect 39773 14841 39807 14875
rect 39807 14841 39816 14875
rect 41788 15011 41840 15020
rect 41788 14977 41797 15011
rect 41797 14977 41831 15011
rect 41831 14977 41840 15011
rect 41788 14968 41840 14977
rect 45560 15104 45612 15156
rect 46756 15147 46808 15156
rect 46756 15113 46765 15147
rect 46765 15113 46799 15147
rect 46799 15113 46808 15147
rect 46756 15104 46808 15113
rect 48412 15104 48464 15156
rect 52644 15104 52696 15156
rect 53196 15104 53248 15156
rect 54760 15104 54812 15156
rect 57152 15104 57204 15156
rect 44640 14900 44692 14952
rect 48044 14943 48096 14952
rect 48044 14909 48053 14943
rect 48053 14909 48087 14943
rect 48087 14909 48096 14943
rect 48044 14900 48096 14909
rect 48688 15079 48740 15088
rect 48688 15045 48697 15079
rect 48697 15045 48731 15079
rect 48731 15045 48740 15079
rect 48688 15036 48740 15045
rect 50896 15036 50948 15088
rect 49424 15011 49476 15020
rect 49424 14977 49433 15011
rect 49433 14977 49467 15011
rect 49467 14977 49476 15011
rect 49424 14968 49476 14977
rect 49516 14968 49568 15020
rect 49700 15011 49752 15020
rect 49700 14977 49709 15011
rect 49709 14977 49743 15011
rect 49743 14977 49752 15011
rect 49700 14968 49752 14977
rect 50620 15011 50672 15020
rect 50620 14977 50629 15011
rect 50629 14977 50663 15011
rect 50663 14977 50672 15011
rect 50620 14968 50672 14977
rect 52000 14968 52052 15020
rect 54116 15036 54168 15088
rect 49976 14943 50028 14952
rect 39764 14832 39816 14841
rect 34336 14764 34388 14773
rect 36544 14764 36596 14816
rect 39304 14807 39356 14816
rect 39304 14773 39313 14807
rect 39313 14773 39347 14807
rect 39347 14773 39356 14807
rect 39304 14764 39356 14773
rect 42156 14807 42208 14816
rect 42156 14773 42165 14807
rect 42165 14773 42199 14807
rect 42199 14773 42208 14807
rect 42156 14764 42208 14773
rect 44732 14764 44784 14816
rect 46572 14807 46624 14816
rect 46572 14773 46581 14807
rect 46581 14773 46615 14807
rect 46615 14773 46624 14807
rect 49976 14909 49985 14943
rect 49985 14909 50019 14943
rect 50019 14909 50028 14943
rect 49976 14900 50028 14909
rect 46572 14764 46624 14773
rect 50804 14764 50856 14816
rect 56232 14968 56284 15020
rect 57980 14968 58032 15020
rect 52092 14764 52144 14816
rect 55220 14764 55272 14816
rect 56140 14764 56192 14816
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 22616 14662 22668 14714
rect 22680 14662 22732 14714
rect 22744 14662 22796 14714
rect 22808 14662 22860 14714
rect 22872 14662 22924 14714
rect 37060 14662 37112 14714
rect 37124 14662 37176 14714
rect 37188 14662 37240 14714
rect 37252 14662 37304 14714
rect 37316 14662 37368 14714
rect 51504 14662 51556 14714
rect 51568 14662 51620 14714
rect 51632 14662 51684 14714
rect 51696 14662 51748 14714
rect 51760 14662 51812 14714
rect 4160 14560 4212 14612
rect 6552 14560 6604 14612
rect 8668 14560 8720 14612
rect 9588 14560 9640 14612
rect 12348 14560 12400 14612
rect 13176 14560 13228 14612
rect 14188 14560 14240 14612
rect 19984 14560 20036 14612
rect 6184 14492 6236 14544
rect 12256 14492 12308 14544
rect 4344 14424 4396 14476
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 6644 14424 6696 14476
rect 9864 14424 9916 14476
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2688 14356 2740 14408
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 8024 14356 8076 14408
rect 10600 14399 10652 14408
rect 10600 14365 10609 14399
rect 10609 14365 10643 14399
rect 10643 14365 10652 14399
rect 10600 14356 10652 14365
rect 12992 14356 13044 14408
rect 13544 14356 13596 14408
rect 17224 14356 17276 14408
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 22376 14560 22428 14612
rect 32312 14560 32364 14612
rect 32404 14560 32456 14612
rect 38200 14603 38252 14612
rect 38200 14569 38209 14603
rect 38209 14569 38243 14603
rect 38243 14569 38252 14603
rect 38200 14560 38252 14569
rect 39764 14560 39816 14612
rect 52000 14560 52052 14612
rect 54300 14560 54352 14612
rect 54852 14560 54904 14612
rect 49424 14492 49476 14544
rect 50528 14535 50580 14544
rect 50528 14501 50537 14535
rect 50537 14501 50571 14535
rect 50571 14501 50580 14535
rect 50528 14492 50580 14501
rect 2504 14220 2556 14272
rect 6276 14220 6328 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 20720 14356 20772 14408
rect 22468 14356 22520 14408
rect 25412 14399 25464 14408
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 26792 14356 26844 14408
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 34336 14399 34388 14408
rect 34336 14365 34345 14399
rect 34345 14365 34379 14399
rect 34379 14365 34388 14399
rect 34336 14356 34388 14365
rect 34980 14356 35032 14408
rect 38568 14356 38620 14408
rect 40408 14399 40460 14408
rect 40408 14365 40417 14399
rect 40417 14365 40451 14399
rect 40451 14365 40460 14399
rect 40408 14356 40460 14365
rect 43076 14399 43128 14408
rect 43076 14365 43085 14399
rect 43085 14365 43119 14399
rect 43119 14365 43128 14399
rect 43076 14356 43128 14365
rect 44916 14356 44968 14408
rect 49148 14399 49200 14408
rect 49148 14365 49157 14399
rect 49157 14365 49191 14399
rect 49191 14365 49200 14399
rect 49148 14356 49200 14365
rect 52092 14467 52144 14476
rect 52092 14433 52101 14467
rect 52101 14433 52135 14467
rect 52135 14433 52144 14467
rect 52092 14424 52144 14433
rect 24032 14288 24084 14340
rect 30196 14288 30248 14340
rect 31116 14288 31168 14340
rect 37832 14288 37884 14340
rect 47952 14288 48004 14340
rect 50896 14288 50948 14340
rect 53656 14399 53708 14408
rect 53656 14365 53665 14399
rect 53665 14365 53699 14399
rect 53699 14365 53708 14399
rect 53656 14356 53708 14365
rect 57888 14288 57940 14340
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9864 14220 9916 14272
rect 15292 14220 15344 14272
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 17592 14220 17644 14272
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 18420 14220 18472 14272
rect 20996 14220 21048 14272
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25596 14263 25648 14272
rect 25596 14229 25605 14263
rect 25605 14229 25639 14263
rect 25639 14229 25648 14263
rect 25596 14220 25648 14229
rect 26056 14220 26108 14272
rect 29736 14220 29788 14272
rect 30288 14263 30340 14272
rect 30288 14229 30297 14263
rect 30297 14229 30331 14263
rect 30331 14229 30340 14263
rect 30288 14220 30340 14229
rect 32220 14263 32272 14272
rect 32220 14229 32229 14263
rect 32229 14229 32263 14263
rect 32263 14229 32272 14263
rect 32220 14220 32272 14229
rect 32864 14263 32916 14272
rect 32864 14229 32873 14263
rect 32873 14229 32907 14263
rect 32907 14229 32916 14263
rect 32864 14220 32916 14229
rect 33784 14263 33836 14272
rect 33784 14229 33793 14263
rect 33793 14229 33827 14263
rect 33827 14229 33836 14263
rect 33784 14220 33836 14229
rect 34704 14263 34756 14272
rect 34704 14229 34713 14263
rect 34713 14229 34747 14263
rect 34747 14229 34756 14263
rect 34704 14220 34756 14229
rect 37464 14263 37516 14272
rect 37464 14229 37473 14263
rect 37473 14229 37507 14263
rect 37507 14229 37516 14263
rect 37464 14220 37516 14229
rect 42524 14263 42576 14272
rect 42524 14229 42533 14263
rect 42533 14229 42567 14263
rect 42567 14229 42576 14263
rect 42524 14220 42576 14229
rect 43812 14220 43864 14272
rect 44640 14220 44692 14272
rect 47032 14220 47084 14272
rect 50528 14220 50580 14272
rect 53012 14220 53064 14272
rect 56784 14263 56836 14272
rect 56784 14229 56793 14263
rect 56793 14229 56827 14263
rect 56827 14229 56836 14263
rect 56784 14220 56836 14229
rect 57336 14263 57388 14272
rect 57336 14229 57345 14263
rect 57345 14229 57379 14263
rect 57379 14229 57388 14263
rect 57336 14220 57388 14229
rect 15394 14118 15446 14170
rect 15458 14118 15510 14170
rect 15522 14118 15574 14170
rect 15586 14118 15638 14170
rect 15650 14118 15702 14170
rect 29838 14118 29890 14170
rect 29902 14118 29954 14170
rect 29966 14118 30018 14170
rect 30030 14118 30082 14170
rect 30094 14118 30146 14170
rect 44282 14118 44334 14170
rect 44346 14118 44398 14170
rect 44410 14118 44462 14170
rect 44474 14118 44526 14170
rect 44538 14118 44590 14170
rect 58726 14118 58778 14170
rect 58790 14118 58842 14170
rect 58854 14118 58906 14170
rect 58918 14118 58970 14170
rect 58982 14118 59034 14170
rect 2872 14016 2924 14068
rect 3792 14016 3844 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 5816 14016 5868 14068
rect 6644 14016 6696 14068
rect 8944 14016 8996 14068
rect 9128 14016 9180 14068
rect 10600 14016 10652 14068
rect 11888 14016 11940 14068
rect 12532 14059 12584 14068
rect 12532 14025 12541 14059
rect 12541 14025 12575 14059
rect 12575 14025 12584 14059
rect 12532 14016 12584 14025
rect 12716 14016 12768 14068
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 13728 14016 13780 14068
rect 2504 13948 2556 14000
rect 2044 13880 2096 13932
rect 2228 13880 2280 13932
rect 3976 13923 4028 13932
rect 3976 13889 3985 13923
rect 3985 13889 4019 13923
rect 4019 13889 4028 13923
rect 3976 13880 4028 13889
rect 5264 13948 5316 14000
rect 8576 13948 8628 14000
rect 6736 13880 6788 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 4712 13812 4764 13864
rect 3516 13787 3568 13796
rect 3516 13753 3525 13787
rect 3525 13753 3559 13787
rect 3559 13753 3568 13787
rect 3516 13744 3568 13753
rect 9496 13948 9548 14000
rect 14924 13880 14976 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 10784 13812 10836 13864
rect 11060 13812 11112 13864
rect 11152 13812 11204 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 14372 13855 14424 13864
rect 14372 13821 14381 13855
rect 14381 13821 14415 13855
rect 14415 13821 14424 13855
rect 14372 13812 14424 13821
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 17224 14016 17276 14068
rect 17776 14016 17828 14068
rect 18420 14016 18472 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20628 14016 20680 14068
rect 22284 14016 22336 14068
rect 24860 14016 24912 14068
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19248 13812 19300 13864
rect 19432 13812 19484 13864
rect 24032 13880 24084 13932
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 25596 14016 25648 14068
rect 26608 14016 26660 14068
rect 28356 14016 28408 14068
rect 30196 14016 30248 14068
rect 30840 14016 30892 14068
rect 30932 14059 30984 14068
rect 30932 14025 30941 14059
rect 30941 14025 30975 14059
rect 30975 14025 30984 14059
rect 30932 14016 30984 14025
rect 33968 14016 34020 14068
rect 18236 13744 18288 13796
rect 22376 13855 22428 13864
rect 22376 13821 22385 13855
rect 22385 13821 22419 13855
rect 22419 13821 22428 13855
rect 22376 13812 22428 13821
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 25780 13880 25832 13889
rect 26792 13880 26844 13932
rect 25228 13744 25280 13796
rect 27528 13812 27580 13864
rect 32864 13880 32916 13932
rect 27804 13812 27856 13864
rect 31116 13855 31168 13864
rect 31116 13821 31125 13855
rect 31125 13821 31159 13855
rect 31159 13821 31168 13855
rect 31116 13812 31168 13821
rect 31208 13812 31260 13864
rect 32312 13812 32364 13864
rect 32680 13855 32732 13864
rect 32680 13821 32689 13855
rect 32689 13821 32723 13855
rect 32723 13821 32732 13855
rect 32680 13812 32732 13821
rect 33784 13880 33836 13932
rect 34152 13880 34204 13932
rect 37464 14016 37516 14068
rect 39304 14016 39356 14068
rect 40408 14016 40460 14068
rect 47952 14059 48004 14068
rect 47952 14025 47961 14059
rect 47961 14025 47995 14059
rect 47995 14025 48004 14059
rect 47952 14016 48004 14025
rect 41604 13948 41656 14000
rect 34244 13744 34296 13796
rect 37740 13923 37792 13932
rect 37740 13889 37749 13923
rect 37749 13889 37783 13923
rect 37783 13889 37792 13923
rect 37740 13880 37792 13889
rect 40500 13923 40552 13932
rect 34796 13812 34848 13864
rect 35348 13812 35400 13864
rect 37832 13855 37884 13864
rect 37832 13821 37841 13855
rect 37841 13821 37875 13855
rect 37875 13821 37884 13855
rect 37832 13812 37884 13821
rect 38844 13855 38896 13864
rect 38844 13821 38853 13855
rect 38853 13821 38887 13855
rect 38887 13821 38896 13855
rect 40500 13889 40509 13923
rect 40509 13889 40543 13923
rect 40543 13889 40552 13923
rect 40500 13880 40552 13889
rect 50620 14016 50672 14068
rect 50896 13948 50948 14000
rect 38844 13812 38896 13821
rect 39580 13855 39632 13864
rect 39580 13821 39589 13855
rect 39589 13821 39623 13855
rect 39623 13821 39632 13855
rect 39580 13812 39632 13821
rect 42616 13812 42668 13864
rect 44272 13812 44324 13864
rect 45284 13812 45336 13864
rect 46572 13812 46624 13864
rect 47400 13855 47452 13864
rect 47400 13821 47409 13855
rect 47409 13821 47443 13855
rect 47443 13821 47452 13855
rect 47400 13812 47452 13821
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 11888 13676 11940 13728
rect 14464 13676 14516 13728
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 18144 13676 18196 13728
rect 22100 13676 22152 13728
rect 28172 13719 28224 13728
rect 28172 13685 28181 13719
rect 28181 13685 28215 13719
rect 28215 13685 28224 13719
rect 28172 13676 28224 13685
rect 29276 13719 29328 13728
rect 29276 13685 29285 13719
rect 29285 13685 29319 13719
rect 29319 13685 29328 13719
rect 29276 13676 29328 13685
rect 31392 13676 31444 13728
rect 32128 13719 32180 13728
rect 32128 13685 32137 13719
rect 32137 13685 32171 13719
rect 32171 13685 32180 13719
rect 32128 13676 32180 13685
rect 32956 13676 33008 13728
rect 35256 13719 35308 13728
rect 35256 13685 35265 13719
rect 35265 13685 35299 13719
rect 35299 13685 35308 13719
rect 35256 13676 35308 13685
rect 36452 13719 36504 13728
rect 36452 13685 36461 13719
rect 36461 13685 36495 13719
rect 36495 13685 36504 13719
rect 36452 13676 36504 13685
rect 38108 13744 38160 13796
rect 38292 13676 38344 13728
rect 39120 13676 39172 13728
rect 40224 13719 40276 13728
rect 40224 13685 40233 13719
rect 40233 13685 40267 13719
rect 40267 13685 40276 13719
rect 40224 13676 40276 13685
rect 42248 13719 42300 13728
rect 42248 13685 42257 13719
rect 42257 13685 42291 13719
rect 42291 13685 42300 13719
rect 42248 13676 42300 13685
rect 43168 13676 43220 13728
rect 44916 13676 44968 13728
rect 46756 13719 46808 13728
rect 46756 13685 46765 13719
rect 46765 13685 46799 13719
rect 46799 13685 46808 13719
rect 46756 13676 46808 13685
rect 47032 13676 47084 13728
rect 47952 13812 48004 13864
rect 52644 14016 52696 14068
rect 51264 13812 51316 13864
rect 53656 14016 53708 14068
rect 57336 14016 57388 14068
rect 57888 14059 57940 14068
rect 57888 14025 57897 14059
rect 57897 14025 57931 14059
rect 57931 14025 57940 14059
rect 57888 14016 57940 14025
rect 53656 13855 53708 13864
rect 53656 13821 53665 13855
rect 53665 13821 53699 13855
rect 53699 13821 53708 13855
rect 53656 13812 53708 13821
rect 54944 13812 54996 13864
rect 55312 13855 55364 13864
rect 55312 13821 55321 13855
rect 55321 13821 55355 13855
rect 55355 13821 55364 13855
rect 55312 13812 55364 13821
rect 57704 13787 57756 13796
rect 57704 13753 57713 13787
rect 57713 13753 57747 13787
rect 57747 13753 57756 13787
rect 57704 13744 57756 13753
rect 48412 13719 48464 13728
rect 48412 13685 48421 13719
rect 48421 13685 48455 13719
rect 48455 13685 48464 13719
rect 48412 13676 48464 13685
rect 51172 13676 51224 13728
rect 54760 13719 54812 13728
rect 54760 13685 54769 13719
rect 54769 13685 54803 13719
rect 54803 13685 54812 13719
rect 54760 13676 54812 13685
rect 56140 13719 56192 13728
rect 56140 13685 56149 13719
rect 56149 13685 56183 13719
rect 56183 13685 56192 13719
rect 56140 13676 56192 13685
rect 56324 13676 56376 13728
rect 57612 13676 57664 13728
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 22616 13574 22668 13626
rect 22680 13574 22732 13626
rect 22744 13574 22796 13626
rect 22808 13574 22860 13626
rect 22872 13574 22924 13626
rect 37060 13574 37112 13626
rect 37124 13574 37176 13626
rect 37188 13574 37240 13626
rect 37252 13574 37304 13626
rect 37316 13574 37368 13626
rect 51504 13574 51556 13626
rect 51568 13574 51620 13626
rect 51632 13574 51684 13626
rect 51696 13574 51748 13626
rect 51760 13574 51812 13626
rect 12072 13472 12124 13524
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 11888 13336 11940 13388
rect 12164 13336 12216 13388
rect 15200 13472 15252 13524
rect 15476 13472 15528 13524
rect 15108 13404 15160 13456
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 11336 13268 11388 13320
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 13544 13379 13596 13388
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 14464 13336 14516 13388
rect 15752 13336 15804 13388
rect 18604 13472 18656 13524
rect 18696 13472 18748 13524
rect 19340 13472 19392 13524
rect 19432 13472 19484 13524
rect 22376 13472 22428 13524
rect 26056 13472 26108 13524
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 17960 13336 18012 13388
rect 18236 13336 18288 13388
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 22284 13404 22336 13456
rect 27528 13472 27580 13524
rect 27804 13515 27856 13524
rect 27804 13481 27813 13515
rect 27813 13481 27847 13515
rect 27847 13481 27856 13515
rect 27804 13472 27856 13481
rect 32680 13472 32732 13524
rect 19524 13336 19576 13345
rect 21180 13336 21232 13388
rect 10416 13200 10468 13252
rect 14096 13268 14148 13320
rect 14740 13268 14792 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 18144 13268 18196 13320
rect 19616 13268 19668 13320
rect 20168 13268 20220 13320
rect 20996 13311 21048 13320
rect 20996 13277 21005 13311
rect 21005 13277 21039 13311
rect 21039 13277 21048 13311
rect 20996 13268 21048 13277
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 18420 13200 18472 13252
rect 24124 13268 24176 13320
rect 25780 13336 25832 13388
rect 26976 13404 27028 13456
rect 26332 13336 26384 13388
rect 31392 13379 31444 13388
rect 31392 13345 31401 13379
rect 31401 13345 31435 13379
rect 31435 13345 31444 13379
rect 31392 13336 31444 13345
rect 32128 13336 32180 13388
rect 26608 13268 26660 13320
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 27804 13268 27856 13320
rect 29276 13268 29328 13320
rect 29736 13268 29788 13320
rect 30932 13268 30984 13320
rect 31484 13268 31536 13320
rect 32956 13336 33008 13388
rect 34980 13472 35032 13524
rect 35348 13472 35400 13524
rect 38292 13472 38344 13524
rect 38752 13472 38804 13524
rect 40500 13472 40552 13524
rect 33508 13404 33560 13456
rect 33600 13404 33652 13456
rect 34428 13404 34480 13456
rect 35808 13447 35860 13456
rect 35808 13413 35817 13447
rect 35817 13413 35851 13447
rect 35851 13413 35860 13447
rect 35808 13404 35860 13413
rect 34244 13336 34296 13388
rect 34612 13268 34664 13320
rect 34796 13268 34848 13320
rect 35164 13268 35216 13320
rect 35808 13268 35860 13320
rect 38108 13404 38160 13456
rect 38476 13379 38528 13388
rect 38476 13345 38485 13379
rect 38485 13345 38519 13379
rect 38519 13345 38528 13379
rect 38476 13336 38528 13345
rect 39580 13336 39632 13388
rect 40040 13379 40092 13388
rect 40040 13345 40049 13379
rect 40049 13345 40083 13379
rect 40083 13345 40092 13379
rect 40040 13336 40092 13345
rect 42524 13336 42576 13388
rect 43168 13336 43220 13388
rect 44272 13515 44324 13524
rect 44272 13481 44281 13515
rect 44281 13481 44315 13515
rect 44315 13481 44324 13515
rect 44272 13472 44324 13481
rect 49148 13472 49200 13524
rect 49516 13472 49568 13524
rect 51264 13472 51316 13524
rect 43812 13379 43864 13388
rect 43812 13345 43821 13379
rect 43821 13345 43855 13379
rect 43855 13345 43864 13379
rect 43812 13336 43864 13345
rect 46296 13336 46348 13388
rect 29092 13200 29144 13252
rect 31300 13200 31352 13252
rect 32128 13200 32180 13252
rect 34152 13200 34204 13252
rect 36820 13200 36872 13252
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 11060 13132 11112 13184
rect 11244 13132 11296 13184
rect 13268 13132 13320 13184
rect 14464 13175 14516 13184
rect 14464 13141 14473 13175
rect 14473 13141 14507 13175
rect 14507 13141 14516 13175
rect 14464 13132 14516 13141
rect 14832 13175 14884 13184
rect 14832 13141 14841 13175
rect 14841 13141 14875 13175
rect 14875 13141 14884 13175
rect 14832 13132 14884 13141
rect 16120 13132 16172 13184
rect 19340 13132 19392 13184
rect 19616 13175 19668 13184
rect 19616 13141 19625 13175
rect 19625 13141 19659 13175
rect 19659 13141 19668 13175
rect 19616 13132 19668 13141
rect 23572 13175 23624 13184
rect 23572 13141 23581 13175
rect 23581 13141 23615 13175
rect 23615 13141 23624 13175
rect 23572 13132 23624 13141
rect 23664 13132 23716 13184
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 25780 13132 25832 13184
rect 26240 13132 26292 13184
rect 31116 13132 31168 13184
rect 32036 13175 32088 13184
rect 32036 13141 32045 13175
rect 32045 13141 32079 13175
rect 32079 13141 32088 13175
rect 32036 13132 32088 13141
rect 35072 13175 35124 13184
rect 35072 13141 35081 13175
rect 35081 13141 35115 13175
rect 35115 13141 35124 13175
rect 35072 13132 35124 13141
rect 35164 13175 35216 13184
rect 35164 13141 35173 13175
rect 35173 13141 35207 13175
rect 35207 13141 35216 13175
rect 35164 13132 35216 13141
rect 38752 13311 38804 13320
rect 38752 13277 38761 13311
rect 38761 13277 38795 13311
rect 38795 13277 38804 13311
rect 38752 13268 38804 13277
rect 38844 13311 38896 13320
rect 38844 13277 38878 13311
rect 38878 13277 38896 13311
rect 38844 13268 38896 13277
rect 39028 13311 39080 13320
rect 39028 13277 39037 13311
rect 39037 13277 39071 13311
rect 39071 13277 39080 13311
rect 39028 13268 39080 13277
rect 40224 13311 40276 13320
rect 40224 13277 40233 13311
rect 40233 13277 40267 13311
rect 40267 13277 40276 13311
rect 40224 13268 40276 13277
rect 40316 13268 40368 13320
rect 45560 13268 45612 13320
rect 45744 13311 45796 13320
rect 45744 13277 45753 13311
rect 45753 13277 45787 13311
rect 45787 13277 45796 13311
rect 45744 13268 45796 13277
rect 50344 13379 50396 13388
rect 50344 13345 50353 13379
rect 50353 13345 50387 13379
rect 50387 13345 50396 13379
rect 50344 13336 50396 13345
rect 51540 13336 51592 13388
rect 48596 13268 48648 13320
rect 38200 13132 38252 13184
rect 38568 13132 38620 13184
rect 38844 13132 38896 13184
rect 38936 13132 38988 13184
rect 39672 13175 39724 13184
rect 39672 13141 39681 13175
rect 39681 13141 39715 13175
rect 39715 13141 39724 13175
rect 39672 13132 39724 13141
rect 41604 13200 41656 13252
rect 40592 13175 40644 13184
rect 40592 13141 40601 13175
rect 40601 13141 40635 13175
rect 40635 13141 40644 13175
rect 40592 13132 40644 13141
rect 43076 13200 43128 13252
rect 46756 13200 46808 13252
rect 48412 13200 48464 13252
rect 42340 13175 42392 13184
rect 42340 13141 42349 13175
rect 42349 13141 42383 13175
rect 42383 13141 42392 13175
rect 42340 13132 42392 13141
rect 43812 13132 43864 13184
rect 44824 13175 44876 13184
rect 44824 13141 44833 13175
rect 44833 13141 44867 13175
rect 44867 13141 44876 13175
rect 44824 13132 44876 13141
rect 45192 13175 45244 13184
rect 45192 13141 45201 13175
rect 45201 13141 45235 13175
rect 45235 13141 45244 13175
rect 45192 13132 45244 13141
rect 49700 13268 49752 13320
rect 51172 13268 51224 13320
rect 52368 13404 52420 13456
rect 55312 13404 55364 13456
rect 54760 13336 54812 13388
rect 54944 13336 54996 13388
rect 56508 13379 56560 13388
rect 56508 13345 56517 13379
rect 56517 13345 56551 13379
rect 56551 13345 56560 13379
rect 56508 13336 56560 13345
rect 56600 13336 56652 13388
rect 57704 13336 57756 13388
rect 52276 13268 52328 13320
rect 49240 13200 49292 13252
rect 53012 13311 53064 13320
rect 53012 13277 53046 13311
rect 53046 13277 53064 13311
rect 53012 13268 53064 13277
rect 54116 13268 54168 13320
rect 55956 13311 56008 13320
rect 55956 13277 55965 13311
rect 55965 13277 55999 13311
rect 55999 13277 56008 13311
rect 55956 13268 56008 13277
rect 57152 13311 57204 13320
rect 57152 13277 57161 13311
rect 57161 13277 57195 13311
rect 57195 13277 57204 13311
rect 57152 13268 57204 13277
rect 57612 13311 57664 13320
rect 57612 13277 57621 13311
rect 57621 13277 57655 13311
rect 57655 13277 57664 13311
rect 57612 13268 57664 13277
rect 49332 13175 49384 13184
rect 49332 13141 49341 13175
rect 49341 13141 49375 13175
rect 49375 13141 49384 13175
rect 49332 13132 49384 13141
rect 50528 13175 50580 13184
rect 50528 13141 50537 13175
rect 50537 13141 50571 13175
rect 50571 13141 50580 13175
rect 50528 13132 50580 13141
rect 50804 13132 50856 13184
rect 52460 13175 52512 13184
rect 52460 13141 52469 13175
rect 52469 13141 52503 13175
rect 52503 13141 52512 13175
rect 52460 13132 52512 13141
rect 54944 13175 54996 13184
rect 54944 13141 54953 13175
rect 54953 13141 54987 13175
rect 54987 13141 54996 13175
rect 54944 13132 54996 13141
rect 55128 13132 55180 13184
rect 57520 13132 57572 13184
rect 15394 13030 15446 13082
rect 15458 13030 15510 13082
rect 15522 13030 15574 13082
rect 15586 13030 15638 13082
rect 15650 13030 15702 13082
rect 29838 13030 29890 13082
rect 29902 13030 29954 13082
rect 29966 13030 30018 13082
rect 30030 13030 30082 13082
rect 30094 13030 30146 13082
rect 44282 13030 44334 13082
rect 44346 13030 44398 13082
rect 44410 13030 44462 13082
rect 44474 13030 44526 13082
rect 44538 13030 44590 13082
rect 58726 13030 58778 13082
rect 58790 13030 58842 13082
rect 58854 13030 58906 13082
rect 58918 13030 58970 13082
rect 58982 13030 59034 13082
rect 2044 12928 2096 12980
rect 6460 12928 6512 12980
rect 11152 12928 11204 12980
rect 11336 12928 11388 12980
rect 1860 12835 1912 12844
rect 1860 12801 1894 12835
rect 1894 12801 1912 12835
rect 1860 12792 1912 12801
rect 4160 12792 4212 12844
rect 4436 12792 4488 12844
rect 8024 12860 8076 12912
rect 9864 12835 9916 12844
rect 9864 12801 9898 12835
rect 9898 12801 9916 12835
rect 9864 12792 9916 12801
rect 11244 12792 11296 12844
rect 12164 12860 12216 12912
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 11612 12724 11664 12776
rect 13452 12928 13504 12980
rect 13636 12928 13688 12980
rect 14832 12928 14884 12980
rect 18328 12928 18380 12980
rect 19064 12928 19116 12980
rect 19340 12928 19392 12980
rect 20168 12928 20220 12980
rect 20628 12928 20680 12980
rect 23572 12928 23624 12980
rect 24768 12928 24820 12980
rect 25872 12928 25924 12980
rect 26608 12928 26660 12980
rect 27620 12928 27672 12980
rect 28172 12928 28224 12980
rect 29092 12928 29144 12980
rect 29736 12928 29788 12980
rect 14372 12860 14424 12912
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 13084 12792 13136 12844
rect 16948 12903 17000 12912
rect 16948 12869 16982 12903
rect 16982 12869 17000 12903
rect 16948 12860 17000 12869
rect 18420 12860 18472 12912
rect 20260 12903 20312 12912
rect 20260 12869 20269 12903
rect 20269 12869 20303 12903
rect 20303 12869 20312 12903
rect 20260 12860 20312 12869
rect 16304 12792 16356 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 19064 12792 19116 12844
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 19800 12792 19852 12844
rect 15752 12656 15804 12708
rect 11244 12588 11296 12597
rect 14096 12588 14148 12640
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 16304 12588 16356 12640
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 20628 12724 20680 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 19892 12656 19944 12708
rect 22192 12656 22244 12708
rect 25780 12724 25832 12776
rect 27896 12835 27948 12844
rect 27896 12801 27905 12835
rect 27905 12801 27939 12835
rect 27939 12801 27948 12835
rect 27896 12792 27948 12801
rect 29644 12792 29696 12844
rect 31668 12928 31720 12980
rect 32312 12971 32364 12980
rect 32312 12937 32321 12971
rect 32321 12937 32355 12971
rect 32355 12937 32364 12971
rect 32312 12928 32364 12937
rect 34336 12928 34388 12980
rect 35256 12928 35308 12980
rect 38568 12928 38620 12980
rect 39580 12928 39632 12980
rect 41604 12971 41656 12980
rect 41604 12937 41613 12971
rect 41613 12937 41647 12971
rect 41647 12937 41656 12971
rect 41604 12928 41656 12937
rect 42340 12928 42392 12980
rect 43076 12928 43128 12980
rect 43996 12928 44048 12980
rect 30288 12860 30340 12912
rect 31300 12903 31352 12912
rect 31300 12869 31309 12903
rect 31309 12869 31343 12903
rect 31343 12869 31352 12903
rect 31300 12860 31352 12869
rect 32036 12860 32088 12912
rect 34704 12860 34756 12912
rect 36452 12860 36504 12912
rect 37556 12860 37608 12912
rect 37740 12860 37792 12912
rect 37832 12860 37884 12912
rect 38016 12860 38068 12912
rect 39028 12860 39080 12912
rect 27344 12724 27396 12776
rect 27068 12656 27120 12708
rect 16396 12588 16448 12597
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21180 12588 21232 12597
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 23204 12588 23256 12597
rect 25872 12588 25924 12640
rect 27436 12631 27488 12640
rect 27436 12597 27445 12631
rect 27445 12597 27479 12631
rect 27479 12597 27488 12631
rect 31484 12724 31536 12776
rect 34336 12792 34388 12844
rect 34520 12724 34572 12776
rect 35072 12792 35124 12844
rect 35808 12792 35860 12844
rect 39580 12792 39632 12844
rect 43904 12835 43956 12844
rect 43904 12801 43922 12835
rect 43922 12801 43956 12835
rect 43904 12792 43956 12801
rect 43996 12835 44048 12844
rect 43996 12801 44005 12835
rect 44005 12801 44039 12835
rect 44039 12801 44048 12835
rect 43996 12792 44048 12801
rect 45744 12928 45796 12980
rect 47400 12928 47452 12980
rect 47952 12971 48004 12980
rect 47952 12937 47961 12971
rect 47961 12937 47995 12971
rect 47995 12937 48004 12971
rect 47952 12928 48004 12937
rect 48596 12971 48648 12980
rect 48596 12937 48605 12971
rect 48605 12937 48639 12971
rect 48639 12937 48648 12971
rect 48596 12928 48648 12937
rect 49332 12928 49384 12980
rect 50528 12928 50580 12980
rect 51080 12928 51132 12980
rect 51540 12928 51592 12980
rect 52276 12928 52328 12980
rect 54944 12928 54996 12980
rect 55220 12928 55272 12980
rect 56508 12928 56560 12980
rect 56784 12928 56836 12980
rect 57152 12928 57204 12980
rect 46296 12792 46348 12844
rect 46848 12792 46900 12844
rect 49424 12835 49476 12844
rect 49424 12801 49433 12835
rect 49433 12801 49467 12835
rect 49467 12801 49476 12835
rect 49424 12792 49476 12801
rect 49516 12792 49568 12844
rect 49700 12835 49752 12844
rect 49700 12801 49709 12835
rect 49709 12801 49743 12835
rect 49743 12801 49752 12835
rect 49700 12792 49752 12801
rect 50620 12835 50672 12844
rect 50620 12801 50629 12835
rect 50629 12801 50663 12835
rect 50663 12801 50672 12835
rect 50620 12792 50672 12801
rect 55128 12860 55180 12912
rect 55956 12792 56008 12844
rect 56140 12835 56192 12844
rect 56140 12801 56149 12835
rect 56149 12801 56183 12835
rect 56183 12801 56192 12835
rect 56140 12792 56192 12801
rect 57244 12792 57296 12844
rect 35532 12724 35584 12776
rect 37740 12767 37792 12776
rect 37740 12733 37749 12767
rect 37749 12733 37783 12767
rect 37783 12733 37792 12767
rect 37740 12724 37792 12733
rect 31208 12699 31260 12708
rect 31208 12665 31217 12699
rect 31217 12665 31251 12699
rect 31251 12665 31260 12699
rect 31208 12656 31260 12665
rect 36728 12656 36780 12708
rect 27436 12588 27488 12597
rect 28724 12588 28776 12640
rect 32404 12588 32456 12640
rect 34612 12588 34664 12640
rect 37464 12588 37516 12640
rect 37648 12588 37700 12640
rect 38476 12588 38528 12640
rect 40316 12724 40368 12776
rect 40592 12724 40644 12776
rect 41236 12724 41288 12776
rect 42616 12767 42668 12776
rect 42616 12733 42625 12767
rect 42625 12733 42659 12767
rect 42659 12733 42668 12767
rect 42616 12724 42668 12733
rect 44824 12724 44876 12776
rect 44916 12767 44968 12776
rect 44916 12733 44925 12767
rect 44925 12733 44959 12767
rect 44959 12733 44968 12767
rect 44916 12724 44968 12733
rect 47032 12767 47084 12776
rect 47032 12733 47041 12767
rect 47041 12733 47075 12767
rect 47075 12733 47084 12767
rect 47032 12724 47084 12733
rect 47400 12724 47452 12776
rect 49240 12724 49292 12776
rect 49976 12767 50028 12776
rect 42248 12656 42300 12708
rect 44732 12588 44784 12640
rect 45468 12588 45520 12640
rect 47216 12588 47268 12640
rect 48504 12588 48556 12640
rect 49976 12733 49985 12767
rect 49985 12733 50019 12767
rect 50019 12733 50028 12767
rect 49976 12724 50028 12733
rect 50436 12767 50488 12776
rect 50436 12733 50445 12767
rect 50445 12733 50479 12767
rect 50479 12733 50488 12767
rect 50436 12724 50488 12733
rect 51356 12724 51408 12776
rect 52460 12724 52512 12776
rect 55312 12656 55364 12708
rect 52184 12588 52236 12640
rect 55220 12631 55272 12640
rect 55220 12597 55229 12631
rect 55229 12597 55263 12631
rect 55263 12597 55272 12631
rect 55220 12588 55272 12597
rect 57612 12588 57664 12640
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 22616 12486 22668 12538
rect 22680 12486 22732 12538
rect 22744 12486 22796 12538
rect 22808 12486 22860 12538
rect 22872 12486 22924 12538
rect 37060 12486 37112 12538
rect 37124 12486 37176 12538
rect 37188 12486 37240 12538
rect 37252 12486 37304 12538
rect 37316 12486 37368 12538
rect 51504 12486 51556 12538
rect 51568 12486 51620 12538
rect 51632 12486 51684 12538
rect 51696 12486 51748 12538
rect 51760 12486 51812 12538
rect 1860 12384 1912 12436
rect 3700 12384 3752 12436
rect 5540 12384 5592 12436
rect 6000 12384 6052 12436
rect 10416 12427 10468 12436
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 14372 12384 14424 12436
rect 4160 12180 4212 12232
rect 5172 12248 5224 12300
rect 10784 12316 10836 12368
rect 12532 12316 12584 12368
rect 14740 12359 14792 12368
rect 14740 12325 14749 12359
rect 14749 12325 14783 12359
rect 14783 12325 14792 12359
rect 14740 12316 14792 12325
rect 6276 12248 6328 12300
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 5632 12180 5684 12232
rect 6092 12180 6144 12232
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 3332 12044 3384 12096
rect 3608 12044 3660 12096
rect 4252 12044 4304 12096
rect 4528 12044 4580 12096
rect 7104 12044 7156 12096
rect 7564 12044 7616 12096
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 8760 12044 8812 12096
rect 9496 12044 9548 12096
rect 11152 12044 11204 12096
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 12808 12155 12860 12164
rect 12808 12121 12817 12155
rect 12817 12121 12851 12155
rect 12851 12121 12860 12155
rect 14096 12291 14148 12300
rect 14096 12257 14105 12291
rect 14105 12257 14139 12291
rect 14139 12257 14148 12291
rect 14096 12248 14148 12257
rect 19524 12384 19576 12436
rect 20812 12384 20864 12436
rect 27252 12384 27304 12436
rect 27344 12384 27396 12436
rect 31668 12427 31720 12436
rect 31668 12393 31677 12427
rect 31677 12393 31711 12427
rect 31711 12393 31720 12427
rect 31668 12384 31720 12393
rect 34520 12384 34572 12436
rect 35164 12384 35216 12436
rect 36820 12427 36872 12436
rect 36820 12393 36829 12427
rect 36829 12393 36863 12427
rect 36863 12393 36872 12427
rect 36820 12384 36872 12393
rect 37740 12384 37792 12436
rect 38108 12384 38160 12436
rect 12808 12112 12860 12121
rect 16028 12112 16080 12164
rect 16856 12180 16908 12232
rect 24860 12316 24912 12368
rect 22008 12248 22060 12300
rect 37556 12316 37608 12368
rect 38936 12316 38988 12368
rect 27804 12248 27856 12300
rect 34704 12291 34756 12300
rect 34704 12257 34713 12291
rect 34713 12257 34747 12291
rect 34747 12257 34756 12291
rect 34704 12248 34756 12257
rect 37464 12291 37516 12300
rect 37464 12257 37473 12291
rect 37473 12257 37507 12291
rect 37507 12257 37516 12291
rect 37464 12248 37516 12257
rect 38292 12291 38344 12300
rect 38292 12257 38301 12291
rect 38301 12257 38335 12291
rect 38335 12257 38344 12291
rect 38292 12248 38344 12257
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 26976 12180 27028 12232
rect 27068 12180 27120 12232
rect 18696 12112 18748 12164
rect 19984 12112 20036 12164
rect 22100 12112 22152 12164
rect 24492 12112 24544 12164
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 19340 12044 19392 12096
rect 21824 12087 21876 12096
rect 21824 12053 21833 12087
rect 21833 12053 21867 12087
rect 21867 12053 21876 12087
rect 21824 12044 21876 12053
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 24308 12044 24360 12096
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 25872 12087 25924 12096
rect 25872 12053 25881 12087
rect 25881 12053 25915 12087
rect 25915 12053 25924 12087
rect 25872 12044 25924 12053
rect 26516 12155 26568 12164
rect 26516 12121 26550 12155
rect 26550 12121 26568 12155
rect 26516 12112 26568 12121
rect 26608 12112 26660 12164
rect 29552 12155 29604 12164
rect 29552 12121 29561 12155
rect 29561 12121 29595 12155
rect 29595 12121 29604 12155
rect 29552 12112 29604 12121
rect 31024 12180 31076 12232
rect 36176 12180 36228 12232
rect 36268 12223 36320 12232
rect 36268 12189 36277 12223
rect 36277 12189 36311 12223
rect 36311 12189 36320 12223
rect 36268 12180 36320 12189
rect 36728 12180 36780 12232
rect 42156 12384 42208 12436
rect 46848 12427 46900 12436
rect 46848 12393 46857 12427
rect 46857 12393 46891 12427
rect 46891 12393 46900 12427
rect 46848 12384 46900 12393
rect 47032 12384 47084 12436
rect 48504 12427 48556 12436
rect 48504 12393 48513 12427
rect 48513 12393 48547 12427
rect 48547 12393 48556 12427
rect 48504 12384 48556 12393
rect 48596 12384 48648 12436
rect 43904 12316 43956 12368
rect 42524 12248 42576 12300
rect 42708 12248 42760 12300
rect 43996 12248 44048 12300
rect 50436 12316 50488 12368
rect 52460 12384 52512 12436
rect 54116 12427 54168 12436
rect 54116 12393 54125 12427
rect 54125 12393 54159 12427
rect 54159 12393 54168 12427
rect 54116 12384 54168 12393
rect 54300 12384 54352 12436
rect 57244 12427 57296 12436
rect 57244 12393 57253 12427
rect 57253 12393 57287 12427
rect 57287 12393 57296 12427
rect 57244 12384 57296 12393
rect 41236 12223 41288 12232
rect 33324 12112 33376 12164
rect 38108 12112 38160 12164
rect 40316 12112 40368 12164
rect 41236 12189 41245 12223
rect 41245 12189 41279 12223
rect 41279 12189 41288 12223
rect 41236 12180 41288 12189
rect 45468 12248 45520 12300
rect 47216 12248 47268 12300
rect 51540 12291 51592 12300
rect 51540 12257 51549 12291
rect 51549 12257 51583 12291
rect 51583 12257 51592 12291
rect 51540 12248 51592 12257
rect 52184 12291 52236 12300
rect 52184 12257 52193 12291
rect 52193 12257 52227 12291
rect 52227 12257 52236 12291
rect 52184 12248 52236 12257
rect 54484 12248 54536 12300
rect 30656 12044 30708 12096
rect 32036 12087 32088 12096
rect 32036 12053 32045 12087
rect 32045 12053 32079 12087
rect 32079 12053 32088 12087
rect 32036 12044 32088 12053
rect 35716 12087 35768 12096
rect 35716 12053 35725 12087
rect 35725 12053 35759 12087
rect 35759 12053 35768 12087
rect 35716 12044 35768 12053
rect 36452 12044 36504 12096
rect 36636 12087 36688 12096
rect 36636 12053 36645 12087
rect 36645 12053 36679 12087
rect 36679 12053 36688 12087
rect 36636 12044 36688 12053
rect 40224 12044 40276 12096
rect 42432 12112 42484 12164
rect 44640 12112 44692 12164
rect 45192 12180 45244 12232
rect 45560 12180 45612 12232
rect 47400 12223 47452 12232
rect 47400 12189 47409 12223
rect 47409 12189 47443 12223
rect 47443 12189 47452 12223
rect 47400 12180 47452 12189
rect 42708 12087 42760 12096
rect 42708 12053 42717 12087
rect 42717 12053 42751 12087
rect 42751 12053 42760 12087
rect 42708 12044 42760 12053
rect 42892 12044 42944 12096
rect 43812 12044 43864 12096
rect 48780 12087 48832 12096
rect 48780 12053 48789 12087
rect 48789 12053 48823 12087
rect 48823 12053 48832 12087
rect 48780 12044 48832 12053
rect 49424 12044 49476 12096
rect 57612 12180 57664 12232
rect 56232 12087 56284 12096
rect 56232 12053 56241 12087
rect 56241 12053 56275 12087
rect 56275 12053 56284 12087
rect 56232 12044 56284 12053
rect 56784 12087 56836 12096
rect 56784 12053 56793 12087
rect 56793 12053 56827 12087
rect 56827 12053 56836 12087
rect 56784 12044 56836 12053
rect 57612 12044 57664 12096
rect 15394 11942 15446 11994
rect 15458 11942 15510 11994
rect 15522 11942 15574 11994
rect 15586 11942 15638 11994
rect 15650 11942 15702 11994
rect 29838 11942 29890 11994
rect 29902 11942 29954 11994
rect 29966 11942 30018 11994
rect 30030 11942 30082 11994
rect 30094 11942 30146 11994
rect 44282 11942 44334 11994
rect 44346 11942 44398 11994
rect 44410 11942 44462 11994
rect 44474 11942 44526 11994
rect 44538 11942 44590 11994
rect 58726 11942 58778 11994
rect 58790 11942 58842 11994
rect 58854 11942 58906 11994
rect 58918 11942 58970 11994
rect 58982 11942 59034 11994
rect 4252 11840 4304 11892
rect 4528 11883 4580 11892
rect 4528 11849 4537 11883
rect 4537 11849 4571 11883
rect 4571 11849 4580 11883
rect 4528 11840 4580 11849
rect 4804 11772 4856 11824
rect 3976 11636 4028 11688
rect 4528 11704 4580 11756
rect 6092 11883 6144 11892
rect 6092 11849 6101 11883
rect 6101 11849 6135 11883
rect 6135 11849 6144 11883
rect 6092 11840 6144 11849
rect 7748 11840 7800 11892
rect 9680 11840 9732 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 19984 11883 20036 11892
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 5632 11704 5684 11756
rect 13544 11772 13596 11824
rect 16396 11772 16448 11824
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 9404 11704 9456 11756
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 16764 11704 16816 11756
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 21824 11840 21876 11892
rect 20260 11772 20312 11824
rect 18328 11704 18380 11756
rect 19432 11704 19484 11756
rect 4344 11500 4396 11552
rect 4896 11500 4948 11552
rect 5540 11500 5592 11552
rect 6276 11500 6328 11552
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8024 11500 8076 11552
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 9956 11636 10008 11688
rect 14556 11636 14608 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 8944 11500 8996 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 14372 11500 14424 11552
rect 15108 11500 15160 11552
rect 16580 11500 16632 11552
rect 20628 11568 20680 11620
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 22284 11840 22336 11892
rect 23480 11840 23532 11892
rect 24032 11883 24084 11892
rect 24032 11849 24041 11883
rect 24041 11849 24075 11883
rect 24075 11849 24084 11883
rect 24032 11840 24084 11849
rect 24400 11840 24452 11892
rect 25780 11840 25832 11892
rect 26516 11840 26568 11892
rect 31116 11883 31168 11892
rect 31116 11849 31125 11883
rect 31125 11849 31159 11883
rect 31159 11849 31168 11883
rect 31116 11840 31168 11849
rect 32772 11883 32824 11892
rect 32772 11849 32781 11883
rect 32781 11849 32815 11883
rect 32815 11849 32824 11883
rect 32772 11840 32824 11849
rect 33508 11840 33560 11892
rect 36268 11840 36320 11892
rect 24308 11704 24360 11756
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 36728 11772 36780 11824
rect 22468 11679 22520 11688
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 22284 11568 22336 11620
rect 23572 11636 23624 11688
rect 24584 11679 24636 11688
rect 24584 11645 24593 11679
rect 24593 11645 24627 11679
rect 24627 11645 24636 11679
rect 24584 11636 24636 11645
rect 24952 11636 25004 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 20260 11543 20312 11552
rect 20260 11509 20269 11543
rect 20269 11509 20303 11543
rect 20303 11509 20312 11543
rect 20260 11500 20312 11509
rect 21272 11500 21324 11552
rect 35348 11704 35400 11756
rect 29092 11636 29144 11688
rect 30564 11636 30616 11688
rect 30932 11636 30984 11688
rect 33140 11679 33192 11688
rect 33140 11645 33149 11679
rect 33149 11645 33183 11679
rect 33183 11645 33192 11679
rect 33140 11636 33192 11645
rect 34428 11679 34480 11688
rect 34428 11645 34437 11679
rect 34437 11645 34471 11679
rect 34471 11645 34480 11679
rect 34428 11636 34480 11645
rect 36544 11636 36596 11688
rect 23204 11500 23256 11552
rect 23664 11500 23716 11552
rect 31024 11568 31076 11620
rect 32404 11611 32456 11620
rect 32404 11577 32413 11611
rect 32413 11577 32447 11611
rect 32447 11577 32456 11611
rect 37648 11840 37700 11892
rect 38016 11840 38068 11892
rect 39120 11883 39172 11892
rect 39120 11849 39129 11883
rect 39129 11849 39163 11883
rect 39163 11849 39172 11883
rect 39120 11840 39172 11849
rect 39580 11840 39632 11892
rect 39672 11883 39724 11892
rect 39672 11849 39681 11883
rect 39681 11849 39715 11883
rect 39715 11849 39724 11883
rect 39672 11840 39724 11849
rect 42432 11883 42484 11892
rect 42432 11849 42441 11883
rect 42441 11849 42475 11883
rect 42475 11849 42484 11883
rect 42432 11840 42484 11849
rect 42708 11840 42760 11892
rect 43996 11840 44048 11892
rect 46940 11883 46992 11892
rect 46940 11849 46949 11883
rect 46949 11849 46983 11883
rect 46983 11849 46992 11883
rect 46940 11840 46992 11849
rect 51540 11840 51592 11892
rect 54576 11883 54628 11892
rect 54576 11849 54585 11883
rect 54585 11849 54619 11883
rect 54619 11849 54628 11883
rect 54576 11840 54628 11849
rect 55128 11840 55180 11892
rect 37464 11636 37516 11688
rect 37648 11636 37700 11688
rect 38292 11636 38344 11688
rect 42524 11772 42576 11824
rect 44180 11772 44232 11824
rect 49976 11704 50028 11756
rect 55220 11704 55272 11756
rect 32404 11568 32456 11577
rect 26148 11543 26200 11552
rect 26148 11509 26157 11543
rect 26157 11509 26191 11543
rect 26191 11509 26200 11543
rect 26148 11500 26200 11509
rect 26608 11500 26660 11552
rect 29000 11500 29052 11552
rect 29460 11500 29512 11552
rect 33784 11543 33836 11552
rect 33784 11509 33793 11543
rect 33793 11509 33827 11543
rect 33827 11509 33836 11543
rect 33784 11500 33836 11509
rect 33876 11543 33928 11552
rect 33876 11509 33885 11543
rect 33885 11509 33919 11543
rect 33919 11509 33928 11543
rect 33876 11500 33928 11509
rect 37556 11568 37608 11620
rect 45100 11679 45152 11688
rect 45100 11645 45109 11679
rect 45109 11645 45143 11679
rect 45143 11645 45152 11679
rect 45100 11636 45152 11645
rect 45652 11679 45704 11688
rect 45652 11645 45661 11679
rect 45661 11645 45695 11679
rect 45695 11645 45704 11679
rect 45652 11636 45704 11645
rect 48412 11679 48464 11688
rect 48412 11645 48421 11679
rect 48421 11645 48455 11679
rect 48455 11645 48464 11679
rect 48412 11636 48464 11645
rect 49608 11636 49660 11688
rect 50804 11636 50856 11688
rect 57152 11679 57204 11688
rect 57152 11645 57161 11679
rect 57161 11645 57195 11679
rect 57195 11645 57204 11679
rect 57152 11636 57204 11645
rect 43628 11568 43680 11620
rect 43720 11568 43772 11620
rect 44640 11568 44692 11620
rect 41512 11500 41564 11552
rect 43260 11500 43312 11552
rect 47124 11500 47176 11552
rect 47768 11543 47820 11552
rect 47768 11509 47777 11543
rect 47777 11509 47811 11543
rect 47811 11509 47820 11543
rect 47768 11500 47820 11509
rect 50712 11543 50764 11552
rect 50712 11509 50721 11543
rect 50721 11509 50755 11543
rect 50755 11509 50764 11543
rect 50712 11500 50764 11509
rect 51264 11500 51316 11552
rect 56600 11543 56652 11552
rect 56600 11509 56609 11543
rect 56609 11509 56643 11543
rect 56643 11509 56652 11543
rect 56600 11500 56652 11509
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 22616 11398 22668 11450
rect 22680 11398 22732 11450
rect 22744 11398 22796 11450
rect 22808 11398 22860 11450
rect 22872 11398 22924 11450
rect 37060 11398 37112 11450
rect 37124 11398 37176 11450
rect 37188 11398 37240 11450
rect 37252 11398 37304 11450
rect 37316 11398 37368 11450
rect 51504 11398 51556 11450
rect 51568 11398 51620 11450
rect 51632 11398 51684 11450
rect 51696 11398 51748 11450
rect 51760 11398 51812 11450
rect 3608 11339 3660 11348
rect 3608 11305 3617 11339
rect 3617 11305 3651 11339
rect 3651 11305 3660 11339
rect 3608 11296 3660 11305
rect 4160 11339 4212 11348
rect 4160 11305 4169 11339
rect 4169 11305 4203 11339
rect 4203 11305 4212 11339
rect 4160 11296 4212 11305
rect 4344 11296 4396 11348
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 9312 11296 9364 11348
rect 9864 11296 9916 11348
rect 11888 11296 11940 11348
rect 12808 11296 12860 11348
rect 13452 11296 13504 11348
rect 17316 11296 17368 11348
rect 19524 11296 19576 11348
rect 20352 11296 20404 11348
rect 8760 11160 8812 11212
rect 10048 11228 10100 11280
rect 10784 11228 10836 11280
rect 14096 11228 14148 11280
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 3884 11092 3936 11144
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4436 11092 4488 11144
rect 3240 11067 3292 11076
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 3976 11024 4028 11076
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 4988 11092 5040 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9680 11092 9732 11144
rect 4804 11024 4856 11076
rect 4252 10956 4304 11008
rect 4712 10956 4764 11008
rect 5632 10956 5684 11008
rect 9220 11024 9272 11076
rect 9864 11024 9916 11076
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 13912 11092 13964 11144
rect 16488 11160 16540 11212
rect 16580 11160 16632 11212
rect 16672 11092 16724 11144
rect 19616 11160 19668 11212
rect 22100 11296 22152 11348
rect 24492 11296 24544 11348
rect 24768 11296 24820 11348
rect 22468 11228 22520 11280
rect 18972 11135 19024 11144
rect 18972 11101 18981 11135
rect 18981 11101 19015 11135
rect 19015 11101 19024 11135
rect 18972 11092 19024 11101
rect 23572 11160 23624 11212
rect 23940 11160 23992 11212
rect 26608 11203 26660 11212
rect 26608 11169 26617 11203
rect 26617 11169 26651 11203
rect 26651 11169 26660 11203
rect 26608 11160 26660 11169
rect 29460 11296 29512 11348
rect 30932 11339 30984 11348
rect 30932 11305 30941 11339
rect 30941 11305 30975 11339
rect 30975 11305 30984 11339
rect 30932 11296 30984 11305
rect 33324 11296 33376 11348
rect 37372 11296 37424 11348
rect 38108 11296 38160 11348
rect 38476 11296 38528 11348
rect 29000 11228 29052 11280
rect 21272 11092 21324 11144
rect 23204 11092 23256 11144
rect 28540 11135 28592 11144
rect 28540 11101 28549 11135
rect 28549 11101 28583 11135
rect 28583 11101 28592 11135
rect 28540 11092 28592 11101
rect 14188 11024 14240 11076
rect 14372 11067 14424 11076
rect 14372 11033 14395 11067
rect 14395 11033 14424 11067
rect 14372 11024 14424 11033
rect 15292 11024 15344 11076
rect 18052 11067 18104 11076
rect 18052 11033 18070 11067
rect 18070 11033 18104 11067
rect 18052 11024 18104 11033
rect 20260 11024 20312 11076
rect 8852 10956 8904 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 9404 10956 9456 11008
rect 11520 10956 11572 11008
rect 11888 10956 11940 11008
rect 17224 10956 17276 11008
rect 17592 10956 17644 11008
rect 20720 10956 20772 11008
rect 22468 11024 22520 11076
rect 21548 10956 21600 11008
rect 23664 11024 23716 11076
rect 26148 11024 26200 11076
rect 31116 11092 31168 11144
rect 32404 11135 32456 11144
rect 32404 11101 32413 11135
rect 32413 11101 32447 11135
rect 32447 11101 32456 11135
rect 32404 11092 32456 11101
rect 36728 11228 36780 11280
rect 34520 11160 34572 11212
rect 36176 11160 36228 11212
rect 36912 11203 36964 11212
rect 36912 11169 36921 11203
rect 36921 11169 36955 11203
rect 36955 11169 36964 11203
rect 36912 11160 36964 11169
rect 37556 11271 37608 11280
rect 37556 11237 37565 11271
rect 37565 11237 37599 11271
rect 37599 11237 37608 11271
rect 37556 11228 37608 11237
rect 40776 11296 40828 11348
rect 44180 11296 44232 11348
rect 37372 11092 37424 11144
rect 37464 11092 37516 11144
rect 26700 10999 26752 11008
rect 26700 10965 26709 10999
rect 26709 10965 26743 10999
rect 26743 10965 26752 10999
rect 26700 10956 26752 10965
rect 27620 10956 27672 11008
rect 27896 10999 27948 11008
rect 27896 10965 27905 10999
rect 27905 10965 27939 10999
rect 27939 10965 27948 10999
rect 27896 10956 27948 10965
rect 28816 10956 28868 11008
rect 29368 10999 29420 11008
rect 29368 10965 29377 10999
rect 29377 10965 29411 10999
rect 29411 10965 29420 10999
rect 29368 10956 29420 10965
rect 29736 10956 29788 11008
rect 30564 11024 30616 11076
rect 32036 11024 32088 11076
rect 34152 11067 34204 11076
rect 34152 11033 34161 11067
rect 34161 11033 34195 11067
rect 34195 11033 34204 11067
rect 34152 11024 34204 11033
rect 34888 11024 34940 11076
rect 35808 11024 35860 11076
rect 34612 10956 34664 11008
rect 36360 10999 36412 11008
rect 36360 10965 36369 10999
rect 36369 10965 36403 10999
rect 36403 10965 36412 10999
rect 36360 10956 36412 10965
rect 36820 10999 36872 11008
rect 36820 10965 36829 10999
rect 36829 10965 36863 10999
rect 36863 10965 36872 10999
rect 36820 10956 36872 10965
rect 38016 11160 38068 11212
rect 38384 11203 38436 11212
rect 38384 11169 38402 11203
rect 38402 11169 38436 11203
rect 38384 11160 38436 11169
rect 39212 11203 39264 11212
rect 39212 11169 39221 11203
rect 39221 11169 39255 11203
rect 39255 11169 39264 11203
rect 43260 11228 43312 11280
rect 43628 11228 43680 11280
rect 39212 11160 39264 11169
rect 38476 11135 38528 11144
rect 38476 11101 38485 11135
rect 38485 11101 38519 11135
rect 38519 11101 38528 11135
rect 38476 11092 38528 11101
rect 39856 11092 39908 11144
rect 45100 11296 45152 11348
rect 50712 11296 50764 11348
rect 45836 11160 45888 11212
rect 48320 11228 48372 11280
rect 46940 11160 46992 11212
rect 50344 11203 50396 11212
rect 50344 11169 50353 11203
rect 50353 11169 50387 11203
rect 50387 11169 50396 11203
rect 50344 11160 50396 11169
rect 51172 11228 51224 11280
rect 51264 11160 51316 11212
rect 55404 11228 55456 11280
rect 44916 11092 44968 11144
rect 47492 11067 47544 11076
rect 47492 11033 47501 11067
rect 47501 11033 47535 11067
rect 47535 11033 47544 11067
rect 47492 11024 47544 11033
rect 48504 11135 48556 11144
rect 48504 11101 48513 11135
rect 48513 11101 48547 11135
rect 48547 11101 48556 11135
rect 48504 11092 48556 11101
rect 51356 11135 51408 11144
rect 51356 11101 51365 11135
rect 51365 11101 51399 11135
rect 51399 11101 51408 11135
rect 51356 11092 51408 11101
rect 53012 11135 53064 11144
rect 53012 11101 53021 11135
rect 53021 11101 53055 11135
rect 53055 11101 53064 11135
rect 53012 11092 53064 11101
rect 38476 10956 38528 11008
rect 38752 10956 38804 11008
rect 42524 10999 42576 11008
rect 42524 10965 42533 10999
rect 42533 10965 42567 10999
rect 42567 10965 42576 10999
rect 42524 10956 42576 10965
rect 42892 10956 42944 11008
rect 45744 10999 45796 11008
rect 45744 10965 45753 10999
rect 45753 10965 45787 10999
rect 45787 10965 45796 10999
rect 45744 10956 45796 10965
rect 46020 10956 46072 11008
rect 47952 10999 48004 11008
rect 47952 10965 47961 10999
rect 47961 10965 47995 10999
rect 47995 10965 48004 10999
rect 47952 10956 48004 10965
rect 48228 10956 48280 11008
rect 48780 10956 48832 11008
rect 49516 11024 49568 11076
rect 50436 11024 50488 11076
rect 49148 10956 49200 11008
rect 52276 10956 52328 11008
rect 52644 10956 52696 11008
rect 55036 11135 55088 11144
rect 55036 11101 55045 11135
rect 55045 11101 55079 11135
rect 55079 11101 55088 11135
rect 55036 11092 55088 11101
rect 56600 11135 56652 11144
rect 56600 11101 56634 11135
rect 56634 11101 56652 11135
rect 56600 11092 56652 11101
rect 56600 10956 56652 11008
rect 57796 11067 57848 11076
rect 57796 11033 57805 11067
rect 57805 11033 57839 11067
rect 57839 11033 57848 11067
rect 57796 11024 57848 11033
rect 15394 10854 15446 10906
rect 15458 10854 15510 10906
rect 15522 10854 15574 10906
rect 15586 10854 15638 10906
rect 15650 10854 15702 10906
rect 29838 10854 29890 10906
rect 29902 10854 29954 10906
rect 29966 10854 30018 10906
rect 30030 10854 30082 10906
rect 30094 10854 30146 10906
rect 44282 10854 44334 10906
rect 44346 10854 44398 10906
rect 44410 10854 44462 10906
rect 44474 10854 44526 10906
rect 44538 10854 44590 10906
rect 58726 10854 58778 10906
rect 58790 10854 58842 10906
rect 58854 10854 58906 10906
rect 58918 10854 58970 10906
rect 58982 10854 59034 10906
rect 4804 10752 4856 10804
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 3148 10616 3200 10668
rect 3884 10616 3936 10668
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6092 10548 6144 10600
rect 8576 10548 8628 10600
rect 11428 10752 11480 10804
rect 11520 10752 11572 10804
rect 11796 10752 11848 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 15292 10752 15344 10804
rect 9680 10684 9732 10736
rect 11244 10684 11296 10736
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9496 10616 9548 10668
rect 10048 10616 10100 10668
rect 8760 10548 8812 10600
rect 3332 10480 3384 10532
rect 4252 10480 4304 10532
rect 4436 10480 4488 10532
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 13912 10684 13964 10736
rect 14740 10684 14792 10736
rect 17132 10752 17184 10804
rect 17592 10752 17644 10804
rect 18972 10752 19024 10804
rect 20812 10752 20864 10804
rect 22100 10752 22152 10804
rect 22376 10752 22428 10804
rect 17040 10684 17092 10736
rect 13360 10659 13412 10668
rect 13360 10625 13394 10659
rect 13394 10625 13412 10659
rect 13360 10616 13412 10625
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 16764 10616 16816 10668
rect 17776 10616 17828 10668
rect 19984 10659 20036 10668
rect 19984 10625 19993 10659
rect 19993 10625 20027 10659
rect 20027 10625 20036 10659
rect 19984 10616 20036 10625
rect 6828 10412 6880 10464
rect 8024 10412 8076 10464
rect 8944 10412 8996 10464
rect 10876 10412 10928 10464
rect 14096 10548 14148 10600
rect 12992 10523 13044 10532
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 15844 10480 15896 10532
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 25504 10752 25556 10804
rect 26700 10752 26752 10804
rect 29736 10752 29788 10804
rect 30656 10752 30708 10804
rect 25228 10684 25280 10736
rect 27436 10684 27488 10736
rect 27896 10684 27948 10736
rect 20444 10616 20496 10668
rect 23664 10659 23716 10668
rect 23664 10625 23673 10659
rect 23673 10625 23707 10659
rect 23707 10625 23716 10659
rect 23664 10616 23716 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24768 10616 24820 10668
rect 24952 10616 25004 10668
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 24124 10548 24176 10600
rect 24492 10548 24544 10600
rect 25412 10548 25464 10600
rect 25688 10548 25740 10600
rect 26516 10616 26568 10668
rect 29368 10659 29420 10668
rect 29368 10625 29377 10659
rect 29377 10625 29411 10659
rect 29411 10625 29420 10659
rect 29368 10616 29420 10625
rect 30932 10659 30984 10668
rect 30932 10625 30950 10659
rect 30950 10625 30984 10659
rect 30932 10616 30984 10625
rect 31024 10659 31076 10668
rect 31024 10625 31033 10659
rect 31033 10625 31067 10659
rect 31067 10625 31076 10659
rect 31024 10616 31076 10625
rect 27620 10548 27672 10600
rect 30564 10548 30616 10600
rect 31300 10591 31352 10600
rect 31300 10557 31309 10591
rect 31309 10557 31343 10591
rect 31343 10557 31352 10591
rect 32772 10616 32824 10668
rect 33416 10616 33468 10668
rect 33784 10684 33836 10736
rect 35716 10684 35768 10736
rect 36912 10727 36964 10736
rect 36912 10693 36921 10727
rect 36921 10693 36955 10727
rect 36955 10693 36964 10727
rect 36912 10684 36964 10693
rect 40776 10752 40828 10804
rect 41236 10752 41288 10804
rect 33876 10616 33928 10668
rect 31300 10548 31352 10557
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16028 10412 16080 10464
rect 18328 10412 18380 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 19248 10412 19300 10464
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 23756 10412 23808 10464
rect 25412 10412 25464 10464
rect 29000 10412 29052 10464
rect 29276 10455 29328 10464
rect 29276 10421 29285 10455
rect 29285 10421 29319 10455
rect 29319 10421 29328 10455
rect 29276 10412 29328 10421
rect 31208 10412 31260 10464
rect 31944 10412 31996 10464
rect 33692 10548 33744 10600
rect 34520 10616 34572 10668
rect 37372 10616 37424 10668
rect 37648 10616 37700 10668
rect 45652 10752 45704 10804
rect 47768 10752 47820 10804
rect 47952 10752 48004 10804
rect 48504 10752 48556 10804
rect 50804 10795 50856 10804
rect 43720 10684 43772 10736
rect 42432 10659 42484 10668
rect 42432 10625 42441 10659
rect 42441 10625 42475 10659
rect 42475 10625 42484 10659
rect 42432 10616 42484 10625
rect 42524 10616 42576 10668
rect 45744 10684 45796 10736
rect 44456 10616 44508 10668
rect 34612 10548 34664 10600
rect 34428 10480 34480 10532
rect 33140 10412 33192 10464
rect 39212 10548 39264 10600
rect 44916 10548 44968 10600
rect 45836 10548 45888 10600
rect 46020 10591 46072 10600
rect 46020 10557 46029 10591
rect 46029 10557 46063 10591
rect 46063 10557 46072 10591
rect 46020 10548 46072 10557
rect 47308 10548 47360 10600
rect 48228 10616 48280 10668
rect 49516 10659 49568 10668
rect 49516 10625 49525 10659
rect 49525 10625 49559 10659
rect 49559 10625 49568 10659
rect 49516 10616 49568 10625
rect 49792 10659 49844 10668
rect 49792 10625 49801 10659
rect 49801 10625 49835 10659
rect 49835 10625 49844 10659
rect 49792 10616 49844 10625
rect 49148 10548 49200 10600
rect 49608 10548 49660 10600
rect 49976 10548 50028 10600
rect 50804 10761 50813 10795
rect 50813 10761 50847 10795
rect 50847 10761 50856 10795
rect 50804 10752 50856 10761
rect 56416 10752 56468 10804
rect 52644 10684 52696 10736
rect 52460 10616 52512 10668
rect 53012 10616 53064 10668
rect 53196 10659 53248 10668
rect 53196 10625 53230 10659
rect 53230 10625 53248 10659
rect 53196 10616 53248 10625
rect 55128 10659 55180 10668
rect 55128 10625 55137 10659
rect 55137 10625 55171 10659
rect 55171 10625 55180 10659
rect 55128 10616 55180 10625
rect 55404 10659 55456 10668
rect 55404 10625 55413 10659
rect 55413 10625 55447 10659
rect 55447 10625 55456 10659
rect 55404 10616 55456 10625
rect 56600 10616 56652 10668
rect 56968 10616 57020 10668
rect 37556 10480 37608 10532
rect 37740 10412 37792 10464
rect 43904 10412 43956 10464
rect 45836 10412 45888 10464
rect 48412 10480 48464 10532
rect 48136 10412 48188 10464
rect 54576 10548 54628 10600
rect 50160 10412 50212 10464
rect 50528 10412 50580 10464
rect 54484 10455 54536 10464
rect 54484 10421 54493 10455
rect 54493 10421 54527 10455
rect 54527 10421 54536 10455
rect 54484 10412 54536 10421
rect 55220 10412 55272 10464
rect 56692 10591 56744 10600
rect 56692 10557 56701 10591
rect 56701 10557 56735 10591
rect 56735 10557 56744 10591
rect 56692 10548 56744 10557
rect 56324 10412 56376 10464
rect 56600 10412 56652 10464
rect 56784 10412 56836 10464
rect 57888 10455 57940 10464
rect 57888 10421 57897 10455
rect 57897 10421 57931 10455
rect 57931 10421 57940 10455
rect 57888 10412 57940 10421
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 22616 10310 22668 10362
rect 22680 10310 22732 10362
rect 22744 10310 22796 10362
rect 22808 10310 22860 10362
rect 22872 10310 22924 10362
rect 37060 10310 37112 10362
rect 37124 10310 37176 10362
rect 37188 10310 37240 10362
rect 37252 10310 37304 10362
rect 37316 10310 37368 10362
rect 51504 10310 51556 10362
rect 51568 10310 51620 10362
rect 51632 10310 51684 10362
rect 51696 10310 51748 10362
rect 51760 10310 51812 10362
rect 2872 10208 2924 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 5816 10208 5868 10260
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 9128 10208 9180 10260
rect 9404 10208 9456 10260
rect 10048 10208 10100 10260
rect 13360 10208 13412 10260
rect 14924 10208 14976 10260
rect 15384 10208 15436 10260
rect 15844 10208 15896 10260
rect 16304 10208 16356 10260
rect 9036 10140 9088 10192
rect 2780 10004 2832 10056
rect 3056 9936 3108 9988
rect 6552 10072 6604 10124
rect 6828 10047 6880 10056
rect 6828 10013 6836 10047
rect 6836 10013 6870 10047
rect 6870 10013 6880 10047
rect 6828 10004 6880 10013
rect 9404 10072 9456 10124
rect 7932 10004 7984 10056
rect 7656 9936 7708 9988
rect 6276 9868 6328 9920
rect 8576 10004 8628 10056
rect 8944 10047 8996 10056
rect 8668 9979 8720 9988
rect 8668 9945 8677 9979
rect 8677 9945 8711 9979
rect 8711 9945 8720 9979
rect 8668 9936 8720 9945
rect 8300 9868 8352 9920
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9128 10047 9180 10056
rect 9128 10013 9157 10047
rect 9157 10013 9180 10047
rect 9128 10004 9180 10013
rect 14740 10115 14792 10124
rect 14740 10081 14749 10115
rect 14749 10081 14783 10115
rect 14783 10081 14792 10115
rect 14740 10072 14792 10081
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 16488 10115 16540 10124
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 16672 10072 16724 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 17592 10072 17644 10124
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 20904 10208 20956 10260
rect 23020 10208 23072 10260
rect 25136 10208 25188 10260
rect 28540 10251 28592 10260
rect 28540 10217 28549 10251
rect 28549 10217 28583 10251
rect 28583 10217 28592 10251
rect 28540 10208 28592 10217
rect 29276 10208 29328 10260
rect 20720 10140 20772 10192
rect 21456 10140 21508 10192
rect 22100 10072 22152 10124
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 8852 9936 8904 9988
rect 10048 9936 10100 9988
rect 13820 9936 13872 9988
rect 15292 9936 15344 9988
rect 17776 9936 17828 9988
rect 21456 10004 21508 10056
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 25228 10140 25280 10192
rect 26884 10140 26936 10192
rect 27988 10140 28040 10192
rect 24860 10072 24912 10124
rect 27068 10004 27120 10056
rect 29092 10115 29144 10124
rect 29092 10081 29101 10115
rect 29101 10081 29135 10115
rect 29135 10081 29144 10115
rect 29092 10072 29144 10081
rect 30932 10072 30984 10124
rect 31760 10072 31812 10124
rect 24308 9936 24360 9988
rect 25688 9936 25740 9988
rect 9680 9868 9732 9920
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 17040 9868 17092 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 33416 10004 33468 10056
rect 33508 10004 33560 10056
rect 35808 10251 35860 10260
rect 35808 10217 35817 10251
rect 35817 10217 35851 10251
rect 35851 10217 35860 10251
rect 35808 10208 35860 10217
rect 36820 10208 36872 10260
rect 37464 10251 37516 10260
rect 37464 10217 37473 10251
rect 37473 10217 37507 10251
rect 37507 10217 37516 10251
rect 37464 10208 37516 10217
rect 37648 10183 37700 10192
rect 37648 10149 37657 10183
rect 37657 10149 37691 10183
rect 37691 10149 37700 10183
rect 37648 10140 37700 10149
rect 36360 10115 36412 10124
rect 36360 10081 36369 10115
rect 36369 10081 36403 10115
rect 36403 10081 36412 10115
rect 36360 10072 36412 10081
rect 36728 10072 36780 10124
rect 39856 10183 39908 10192
rect 39856 10149 39865 10183
rect 39865 10149 39899 10183
rect 39899 10149 39908 10183
rect 39856 10140 39908 10149
rect 38844 10072 38896 10124
rect 41236 10115 41288 10124
rect 41236 10081 41245 10115
rect 41245 10081 41279 10115
rect 41279 10081 41288 10115
rect 41236 10072 41288 10081
rect 38752 10047 38804 10056
rect 38752 10013 38761 10047
rect 38761 10013 38795 10047
rect 38795 10013 38804 10047
rect 38752 10004 38804 10013
rect 44456 10208 44508 10260
rect 46204 10251 46256 10260
rect 43444 10072 43496 10124
rect 43904 10115 43956 10124
rect 43904 10081 43913 10115
rect 43913 10081 43947 10115
rect 43947 10081 43956 10115
rect 43904 10072 43956 10081
rect 44180 10115 44232 10124
rect 44180 10081 44189 10115
rect 44189 10081 44223 10115
rect 44223 10081 44232 10115
rect 44180 10072 44232 10081
rect 45652 10072 45704 10124
rect 43628 10047 43680 10056
rect 43628 10013 43637 10047
rect 43637 10013 43671 10047
rect 43671 10013 43680 10047
rect 43628 10004 43680 10013
rect 44640 10047 44692 10056
rect 44640 10013 44649 10047
rect 44649 10013 44683 10047
rect 44683 10013 44692 10047
rect 44640 10004 44692 10013
rect 46204 10217 46213 10251
rect 46213 10217 46247 10251
rect 46247 10217 46256 10251
rect 46204 10208 46256 10217
rect 49608 10208 49660 10260
rect 49976 10208 50028 10260
rect 51356 10208 51408 10260
rect 53840 10208 53892 10260
rect 55036 10208 55088 10260
rect 56692 10208 56744 10260
rect 57888 10208 57940 10260
rect 48412 10140 48464 10192
rect 52276 10140 52328 10192
rect 21364 9868 21416 9920
rect 23572 9868 23624 9920
rect 23756 9911 23808 9920
rect 23756 9877 23765 9911
rect 23765 9877 23799 9911
rect 23799 9877 23808 9911
rect 23756 9868 23808 9877
rect 24400 9868 24452 9920
rect 27712 9868 27764 9920
rect 28080 9868 28132 9920
rect 28816 9868 28868 9920
rect 29092 9868 29144 9920
rect 30564 9868 30616 9920
rect 31852 9911 31904 9920
rect 31852 9877 31861 9911
rect 31861 9877 31895 9911
rect 31895 9877 31904 9911
rect 31852 9868 31904 9877
rect 31944 9911 31996 9920
rect 31944 9877 31953 9911
rect 31953 9877 31987 9911
rect 31987 9877 31996 9911
rect 31944 9868 31996 9877
rect 33232 9868 33284 9920
rect 41144 9936 41196 9988
rect 41604 9979 41656 9988
rect 41604 9945 41638 9979
rect 41638 9945 41656 9979
rect 41604 9936 41656 9945
rect 44824 9936 44876 9988
rect 45836 9936 45888 9988
rect 48320 10004 48372 10056
rect 49884 10004 49936 10056
rect 52460 10072 52512 10124
rect 38936 9868 38988 9920
rect 39304 9868 39356 9920
rect 45468 9868 45520 9920
rect 49424 9979 49476 9988
rect 49424 9945 49433 9979
rect 49433 9945 49467 9979
rect 49467 9945 49476 9979
rect 49424 9936 49476 9945
rect 51816 9936 51868 9988
rect 49976 9911 50028 9920
rect 49976 9877 49985 9911
rect 49985 9877 50019 9911
rect 50019 9877 50028 9911
rect 49976 9868 50028 9877
rect 50528 9868 50580 9920
rect 52644 9868 52696 9920
rect 54392 10072 54444 10124
rect 55404 10072 55456 10124
rect 57704 10004 57756 10056
rect 54024 9936 54076 9988
rect 54116 9868 54168 9920
rect 56324 9868 56376 9920
rect 15394 9766 15446 9818
rect 15458 9766 15510 9818
rect 15522 9766 15574 9818
rect 15586 9766 15638 9818
rect 15650 9766 15702 9818
rect 29838 9766 29890 9818
rect 29902 9766 29954 9818
rect 29966 9766 30018 9818
rect 30030 9766 30082 9818
rect 30094 9766 30146 9818
rect 44282 9766 44334 9818
rect 44346 9766 44398 9818
rect 44410 9766 44462 9818
rect 44474 9766 44526 9818
rect 44538 9766 44590 9818
rect 58726 9766 58778 9818
rect 58790 9766 58842 9818
rect 58854 9766 58906 9818
rect 58918 9766 58970 9818
rect 58982 9766 59034 9818
rect 3056 9707 3108 9716
rect 3056 9673 3065 9707
rect 3065 9673 3099 9707
rect 3099 9673 3108 9707
rect 3056 9664 3108 9673
rect 2228 9596 2280 9648
rect 3240 9596 3292 9648
rect 3884 9528 3936 9580
rect 4068 9596 4120 9648
rect 6736 9639 6788 9648
rect 6736 9605 6745 9639
rect 6745 9605 6779 9639
rect 6779 9605 6788 9639
rect 6736 9596 6788 9605
rect 7656 9596 7708 9648
rect 8668 9664 8720 9716
rect 9128 9664 9180 9716
rect 12808 9664 12860 9716
rect 19616 9707 19668 9716
rect 19616 9673 19625 9707
rect 19625 9673 19659 9707
rect 19659 9673 19668 9707
rect 19616 9664 19668 9673
rect 22100 9664 22152 9716
rect 33508 9664 33560 9716
rect 33692 9664 33744 9716
rect 41144 9707 41196 9716
rect 41144 9673 41153 9707
rect 41153 9673 41187 9707
rect 41187 9673 41196 9707
rect 41144 9664 41196 9673
rect 41604 9707 41656 9716
rect 41604 9673 41613 9707
rect 41613 9673 41647 9707
rect 41647 9673 41656 9707
rect 41604 9664 41656 9673
rect 42432 9664 42484 9716
rect 43536 9664 43588 9716
rect 45468 9707 45520 9716
rect 45468 9673 45477 9707
rect 45477 9673 45511 9707
rect 45511 9673 45520 9707
rect 45468 9664 45520 9673
rect 8300 9596 8352 9648
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5448 9528 5500 9580
rect 5632 9528 5684 9580
rect 7104 9528 7156 9580
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 9496 9596 9548 9648
rect 15384 9596 15436 9648
rect 16212 9596 16264 9648
rect 18052 9596 18104 9648
rect 5540 9460 5592 9512
rect 7748 9460 7800 9512
rect 6184 9392 6236 9444
rect 4528 9324 4580 9376
rect 6828 9324 6880 9376
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9220 9460 9272 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11888 9460 11940 9512
rect 12072 9460 12124 9512
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 12992 9528 13044 9580
rect 16028 9528 16080 9580
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 16672 9460 16724 9512
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 21364 9596 21416 9648
rect 28080 9596 28132 9648
rect 28816 9596 28868 9648
rect 23480 9571 23532 9580
rect 23480 9537 23489 9571
rect 23489 9537 23523 9571
rect 23523 9537 23532 9571
rect 23480 9528 23532 9537
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 21916 9503 21968 9512
rect 11060 9392 11112 9444
rect 19248 9392 19300 9444
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 12348 9324 12400 9376
rect 13636 9324 13688 9376
rect 15936 9324 15988 9376
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 16304 9324 16356 9376
rect 17040 9324 17092 9376
rect 18604 9324 18656 9376
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 22100 9503 22152 9512
rect 22100 9469 22109 9503
rect 22109 9469 22143 9503
rect 22143 9469 22152 9503
rect 22100 9460 22152 9469
rect 22284 9460 22336 9512
rect 23940 9460 23992 9512
rect 24124 9460 24176 9512
rect 24400 9460 24452 9512
rect 22468 9324 22520 9376
rect 24676 9324 24728 9376
rect 26056 9571 26108 9580
rect 26056 9537 26074 9571
rect 26074 9537 26108 9571
rect 26056 9528 26108 9537
rect 30840 9596 30892 9648
rect 31300 9639 31352 9648
rect 31300 9605 31309 9639
rect 31309 9605 31343 9639
rect 31343 9605 31352 9639
rect 31300 9596 31352 9605
rect 32496 9639 32548 9648
rect 32496 9605 32505 9639
rect 32505 9605 32539 9639
rect 32539 9605 32548 9639
rect 32496 9596 32548 9605
rect 35900 9596 35952 9648
rect 30748 9571 30800 9580
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 27712 9460 27764 9512
rect 28540 9460 28592 9512
rect 31852 9528 31904 9580
rect 33232 9528 33284 9580
rect 34152 9528 34204 9580
rect 39304 9639 39356 9648
rect 39304 9605 39313 9639
rect 39313 9605 39347 9639
rect 39347 9605 39356 9639
rect 39304 9596 39356 9605
rect 39764 9596 39816 9648
rect 43628 9596 43680 9648
rect 36636 9528 36688 9580
rect 38200 9528 38252 9580
rect 38752 9528 38804 9580
rect 38844 9571 38896 9580
rect 38844 9537 38853 9571
rect 38853 9537 38887 9571
rect 38887 9537 38896 9571
rect 38844 9528 38896 9537
rect 39856 9528 39908 9580
rect 42800 9571 42852 9580
rect 42800 9537 42809 9571
rect 42809 9537 42843 9571
rect 42843 9537 42852 9571
rect 42800 9528 42852 9537
rect 42892 9571 42944 9580
rect 42892 9537 42901 9571
rect 42901 9537 42935 9571
rect 42935 9537 42944 9571
rect 42892 9528 42944 9537
rect 36084 9460 36136 9512
rect 37740 9460 37792 9512
rect 26608 9324 26660 9376
rect 27620 9324 27672 9376
rect 29460 9324 29512 9376
rect 31852 9367 31904 9376
rect 31852 9333 31861 9367
rect 31861 9333 31895 9367
rect 31895 9333 31904 9367
rect 31852 9324 31904 9333
rect 32404 9324 32456 9376
rect 34244 9324 34296 9376
rect 35900 9367 35952 9376
rect 35900 9333 35909 9367
rect 35909 9333 35943 9367
rect 35943 9333 35952 9367
rect 35900 9324 35952 9333
rect 37464 9324 37516 9376
rect 38660 9435 38712 9444
rect 38660 9401 38669 9435
rect 38669 9401 38703 9435
rect 38703 9401 38712 9435
rect 38660 9392 38712 9401
rect 38200 9367 38252 9376
rect 38200 9333 38209 9367
rect 38209 9333 38243 9367
rect 38243 9333 38252 9367
rect 38200 9324 38252 9333
rect 38292 9324 38344 9376
rect 39120 9324 39172 9376
rect 42340 9324 42392 9376
rect 43352 9528 43404 9580
rect 44180 9596 44232 9648
rect 44364 9639 44416 9648
rect 44364 9605 44373 9639
rect 44373 9605 44407 9639
rect 44407 9605 44416 9639
rect 44364 9596 44416 9605
rect 44732 9596 44784 9648
rect 48780 9664 48832 9716
rect 49056 9707 49108 9716
rect 49056 9673 49065 9707
rect 49065 9673 49099 9707
rect 49099 9673 49108 9707
rect 49056 9664 49108 9673
rect 49976 9664 50028 9716
rect 51816 9707 51868 9716
rect 51816 9673 51825 9707
rect 51825 9673 51859 9707
rect 51859 9673 51868 9707
rect 51816 9664 51868 9673
rect 53196 9664 53248 9716
rect 47492 9596 47544 9648
rect 44824 9528 44876 9580
rect 46756 9528 46808 9580
rect 48412 9571 48464 9580
rect 48412 9537 48421 9571
rect 48421 9537 48455 9571
rect 48455 9537 48464 9571
rect 48412 9528 48464 9537
rect 51172 9571 51224 9580
rect 51172 9537 51181 9571
rect 51181 9537 51215 9571
rect 51215 9537 51224 9571
rect 51172 9528 51224 9537
rect 53840 9571 53892 9580
rect 53840 9537 53849 9571
rect 53849 9537 53883 9571
rect 53883 9537 53892 9571
rect 53840 9528 53892 9537
rect 54024 9571 54076 9580
rect 54024 9537 54033 9571
rect 54033 9537 54067 9571
rect 54067 9537 54076 9571
rect 54024 9528 54076 9537
rect 54576 9571 54628 9580
rect 54576 9537 54585 9571
rect 54585 9537 54619 9571
rect 54619 9537 54628 9571
rect 54576 9528 54628 9537
rect 44180 9460 44232 9512
rect 45008 9460 45060 9512
rect 46940 9503 46992 9512
rect 46940 9469 46949 9503
rect 46949 9469 46983 9503
rect 46983 9469 46992 9503
rect 46940 9460 46992 9469
rect 56232 9596 56284 9648
rect 56692 9596 56744 9648
rect 57796 9596 57848 9648
rect 58256 9639 58308 9648
rect 58256 9605 58265 9639
rect 58265 9605 58299 9639
rect 58299 9605 58308 9639
rect 58256 9596 58308 9605
rect 57520 9571 57572 9580
rect 55864 9503 55916 9512
rect 55864 9469 55873 9503
rect 55873 9469 55907 9503
rect 55907 9469 55916 9503
rect 55864 9460 55916 9469
rect 47768 9392 47820 9444
rect 45100 9324 45152 9376
rect 45836 9324 45888 9376
rect 46204 9324 46256 9376
rect 47124 9324 47176 9376
rect 48688 9367 48740 9376
rect 48688 9333 48697 9367
rect 48697 9333 48731 9367
rect 48731 9333 48740 9367
rect 48688 9324 48740 9333
rect 49792 9324 49844 9376
rect 51172 9392 51224 9444
rect 52276 9392 52328 9444
rect 57520 9537 57529 9571
rect 57529 9537 57563 9571
rect 57563 9537 57572 9571
rect 57520 9528 57572 9537
rect 58440 9571 58492 9580
rect 58440 9537 58449 9571
rect 58449 9537 58483 9571
rect 58483 9537 58492 9571
rect 58440 9528 58492 9537
rect 56784 9460 56836 9512
rect 56968 9503 57020 9512
rect 56968 9469 56977 9503
rect 56977 9469 57011 9503
rect 57011 9469 57020 9503
rect 56968 9460 57020 9469
rect 57060 9503 57112 9512
rect 57060 9469 57069 9503
rect 57069 9469 57103 9503
rect 57103 9469 57112 9503
rect 57060 9460 57112 9469
rect 53012 9367 53064 9376
rect 53012 9333 53021 9367
rect 53021 9333 53055 9367
rect 53055 9333 53064 9367
rect 53012 9324 53064 9333
rect 53472 9324 53524 9376
rect 56324 9324 56376 9376
rect 57152 9324 57204 9376
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 22616 9222 22668 9274
rect 22680 9222 22732 9274
rect 22744 9222 22796 9274
rect 22808 9222 22860 9274
rect 22872 9222 22924 9274
rect 37060 9222 37112 9274
rect 37124 9222 37176 9274
rect 37188 9222 37240 9274
rect 37252 9222 37304 9274
rect 37316 9222 37368 9274
rect 51504 9222 51556 9274
rect 51568 9222 51620 9274
rect 51632 9222 51684 9274
rect 51696 9222 51748 9274
rect 51760 9222 51812 9274
rect 4344 9120 4396 9172
rect 4988 9120 5040 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 8668 9120 8720 9172
rect 9128 9120 9180 9172
rect 12348 9120 12400 9172
rect 14740 9120 14792 9172
rect 14832 9120 14884 9172
rect 6276 8984 6328 9036
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 7748 8984 7800 9036
rect 15936 9120 15988 9172
rect 19616 9120 19668 9172
rect 22100 9120 22152 9172
rect 23756 9120 23808 9172
rect 30840 9120 30892 9172
rect 30932 9120 30984 9172
rect 31392 9120 31444 9172
rect 36452 9120 36504 9172
rect 37648 9120 37700 9172
rect 23940 9052 23992 9104
rect 24676 9052 24728 9104
rect 29000 9052 29052 9104
rect 25688 9027 25740 9036
rect 3332 8916 3384 8968
rect 5540 8916 5592 8968
rect 2412 8848 2464 8900
rect 5356 8848 5408 8900
rect 8852 8848 8904 8900
rect 9220 8848 9272 8900
rect 9772 8916 9824 8968
rect 11060 8916 11112 8968
rect 11888 8916 11940 8968
rect 12256 8959 12308 8968
rect 12256 8925 12290 8959
rect 12290 8925 12308 8959
rect 9588 8891 9640 8900
rect 9588 8857 9597 8891
rect 9597 8857 9631 8891
rect 9631 8857 9640 8891
rect 9588 8848 9640 8857
rect 12256 8916 12308 8925
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 12348 8848 12400 8900
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 16672 8916 16724 8968
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 6092 8780 6144 8832
rect 9496 8780 9548 8832
rect 13452 8780 13504 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 14648 8780 14700 8832
rect 16948 8780 17000 8832
rect 17960 8848 18012 8900
rect 18696 8780 18748 8832
rect 20444 8916 20496 8968
rect 24032 8916 24084 8968
rect 25688 8993 25697 9027
rect 25697 8993 25731 9027
rect 25731 8993 25740 9027
rect 25688 8984 25740 8993
rect 25872 9027 25924 9036
rect 25872 8993 25881 9027
rect 25881 8993 25915 9027
rect 25915 8993 25924 9027
rect 25872 8984 25924 8993
rect 26608 9027 26660 9036
rect 26608 8993 26617 9027
rect 26617 8993 26651 9027
rect 26651 8993 26660 9027
rect 26608 8984 26660 8993
rect 27712 8959 27764 8968
rect 27712 8925 27746 8959
rect 27746 8925 27764 8959
rect 21824 8848 21876 8900
rect 23204 8848 23256 8900
rect 24860 8848 24912 8900
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 27712 8916 27764 8925
rect 31208 9027 31260 9036
rect 31208 8993 31217 9027
rect 31217 8993 31251 9027
rect 31251 8993 31260 9027
rect 31208 8984 31260 8993
rect 31760 8959 31812 8968
rect 31760 8925 31769 8959
rect 31769 8925 31803 8959
rect 31803 8925 31812 8959
rect 31760 8916 31812 8925
rect 27620 8848 27672 8900
rect 30196 8848 30248 8900
rect 42800 9163 42852 9172
rect 42800 9129 42809 9163
rect 42809 9129 42843 9163
rect 42843 9129 42852 9163
rect 42800 9120 42852 9129
rect 43352 9120 43404 9172
rect 44364 9120 44416 9172
rect 45376 9120 45428 9172
rect 46940 9120 46992 9172
rect 51080 9120 51132 9172
rect 39120 9052 39172 9104
rect 46664 9052 46716 9104
rect 49608 9052 49660 9104
rect 51264 9052 51316 9104
rect 43444 9027 43496 9036
rect 43444 8993 43453 9027
rect 43453 8993 43487 9027
rect 43487 8993 43496 9027
rect 43444 8984 43496 8993
rect 44824 8984 44876 9036
rect 46756 8984 46808 9036
rect 47124 9027 47176 9036
rect 47124 8993 47133 9027
rect 47133 8993 47167 9027
rect 47167 8993 47176 9027
rect 47124 8984 47176 8993
rect 32864 8959 32916 8968
rect 32864 8925 32873 8959
rect 32873 8925 32907 8959
rect 32907 8925 32916 8959
rect 32864 8916 32916 8925
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 30748 8780 30800 8832
rect 31300 8823 31352 8832
rect 31300 8789 31309 8823
rect 31309 8789 31343 8823
rect 31343 8789 31352 8823
rect 31300 8780 31352 8789
rect 31668 8823 31720 8832
rect 31668 8789 31677 8823
rect 31677 8789 31711 8823
rect 31711 8789 31720 8823
rect 31668 8780 31720 8789
rect 33784 8823 33836 8832
rect 33784 8789 33793 8823
rect 33793 8789 33827 8823
rect 33827 8789 33836 8823
rect 33784 8780 33836 8789
rect 34244 8780 34296 8832
rect 36728 8959 36780 8968
rect 36728 8925 36737 8959
rect 36737 8925 36771 8959
rect 36771 8925 36780 8959
rect 36728 8916 36780 8925
rect 38936 8959 38988 8968
rect 38936 8925 38945 8959
rect 38945 8925 38979 8959
rect 38979 8925 38988 8959
rect 38936 8916 38988 8925
rect 40408 8959 40460 8968
rect 40408 8925 40417 8959
rect 40417 8925 40451 8959
rect 40451 8925 40460 8959
rect 40408 8916 40460 8925
rect 48688 8984 48740 9036
rect 40316 8848 40368 8900
rect 48044 8959 48096 8968
rect 48044 8925 48053 8959
rect 48053 8925 48087 8959
rect 48087 8925 48096 8959
rect 48044 8916 48096 8925
rect 49332 8916 49384 8968
rect 49792 8984 49844 9036
rect 52276 8984 52328 9036
rect 55864 9120 55916 9172
rect 56692 9120 56744 9172
rect 53932 9052 53984 9104
rect 56784 9052 56836 9104
rect 51080 8916 51132 8968
rect 53012 8916 53064 8968
rect 54392 9027 54444 9036
rect 54392 8993 54401 9027
rect 54401 8993 54435 9027
rect 54435 8993 54444 9027
rect 54392 8984 54444 8993
rect 57244 8984 57296 9036
rect 57520 9027 57572 9036
rect 57520 8993 57529 9027
rect 57529 8993 57563 9027
rect 57563 8993 57572 9027
rect 57520 8984 57572 8993
rect 54024 8916 54076 8968
rect 54668 8916 54720 8968
rect 44732 8848 44784 8900
rect 48228 8848 48280 8900
rect 50344 8848 50396 8900
rect 51172 8848 51224 8900
rect 51356 8848 51408 8900
rect 57796 8848 57848 8900
rect 36084 8823 36136 8832
rect 36084 8789 36093 8823
rect 36093 8789 36127 8823
rect 36127 8789 36136 8823
rect 36084 8780 36136 8789
rect 36912 8780 36964 8832
rect 39672 8823 39724 8832
rect 39672 8789 39681 8823
rect 39681 8789 39715 8823
rect 39715 8789 39724 8823
rect 39672 8780 39724 8789
rect 40500 8780 40552 8832
rect 42340 8823 42392 8832
rect 42340 8789 42349 8823
rect 42349 8789 42383 8823
rect 42383 8789 42392 8823
rect 42340 8780 42392 8789
rect 45008 8780 45060 8832
rect 45376 8780 45428 8832
rect 45836 8780 45888 8832
rect 47768 8780 47820 8832
rect 48688 8823 48740 8832
rect 48688 8789 48697 8823
rect 48697 8789 48731 8823
rect 48731 8789 48740 8823
rect 48688 8780 48740 8789
rect 49148 8823 49200 8832
rect 49148 8789 49157 8823
rect 49157 8789 49191 8823
rect 49191 8789 49200 8823
rect 49148 8780 49200 8789
rect 50896 8823 50948 8832
rect 50896 8789 50905 8823
rect 50905 8789 50939 8823
rect 50939 8789 50948 8823
rect 50896 8780 50948 8789
rect 52920 8823 52972 8832
rect 52920 8789 52929 8823
rect 52929 8789 52963 8823
rect 52963 8789 52972 8823
rect 52920 8780 52972 8789
rect 53748 8780 53800 8832
rect 56876 8823 56928 8832
rect 56876 8789 56885 8823
rect 56885 8789 56919 8823
rect 56919 8789 56928 8823
rect 56876 8780 56928 8789
rect 57888 8780 57940 8832
rect 58072 8823 58124 8832
rect 58072 8789 58081 8823
rect 58081 8789 58115 8823
rect 58115 8789 58124 8823
rect 58072 8780 58124 8789
rect 15394 8678 15446 8730
rect 15458 8678 15510 8730
rect 15522 8678 15574 8730
rect 15586 8678 15638 8730
rect 15650 8678 15702 8730
rect 29838 8678 29890 8730
rect 29902 8678 29954 8730
rect 29966 8678 30018 8730
rect 30030 8678 30082 8730
rect 30094 8678 30146 8730
rect 44282 8678 44334 8730
rect 44346 8678 44398 8730
rect 44410 8678 44462 8730
rect 44474 8678 44526 8730
rect 44538 8678 44590 8730
rect 58726 8678 58778 8730
rect 58790 8678 58842 8730
rect 58854 8678 58906 8730
rect 58918 8678 58970 8730
rect 58982 8678 59034 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 3884 8576 3936 8628
rect 3792 8508 3844 8560
rect 3332 8440 3384 8492
rect 5540 8551 5592 8560
rect 5540 8517 5549 8551
rect 5549 8517 5583 8551
rect 5583 8517 5592 8551
rect 5540 8508 5592 8517
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 2228 8372 2280 8424
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 4528 8304 4580 8356
rect 5356 8304 5408 8356
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6092 8440 6144 8492
rect 9588 8576 9640 8628
rect 12992 8576 13044 8628
rect 16580 8576 16632 8628
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 21824 8619 21876 8628
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 22468 8576 22520 8628
rect 23204 8619 23256 8628
rect 23204 8585 23213 8619
rect 23213 8585 23247 8619
rect 23247 8585 23256 8619
rect 23204 8576 23256 8585
rect 25228 8576 25280 8628
rect 26056 8576 26108 8628
rect 31300 8576 31352 8628
rect 9496 8508 9548 8560
rect 14832 8508 14884 8560
rect 8668 8440 8720 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 10140 8440 10192 8492
rect 11888 8483 11940 8492
rect 11888 8449 11904 8483
rect 11904 8449 11938 8483
rect 11938 8449 11940 8483
rect 11888 8440 11940 8449
rect 12164 8483 12216 8492
rect 12164 8449 12198 8483
rect 12198 8449 12216 8483
rect 12164 8440 12216 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13452 8440 13504 8492
rect 14924 8483 14976 8492
rect 14924 8449 14958 8483
rect 14958 8449 14976 8483
rect 14924 8440 14976 8449
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 8576 8304 8628 8356
rect 9404 8304 9456 8356
rect 11428 8304 11480 8356
rect 13544 8304 13596 8356
rect 13820 8304 13872 8356
rect 16856 8304 16908 8356
rect 21180 8440 21232 8492
rect 19156 8372 19208 8424
rect 23572 8440 23624 8492
rect 23480 8372 23532 8424
rect 23664 8372 23716 8424
rect 28448 8440 28500 8492
rect 30564 8483 30616 8492
rect 30564 8449 30573 8483
rect 30573 8449 30607 8483
rect 30607 8449 30616 8483
rect 30564 8440 30616 8449
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 33416 8576 33468 8628
rect 35900 8576 35952 8628
rect 36728 8576 36780 8628
rect 38936 8576 38988 8628
rect 39672 8576 39724 8628
rect 39764 8619 39816 8628
rect 39764 8585 39773 8619
rect 39773 8585 39807 8619
rect 39807 8585 39816 8619
rect 39764 8576 39816 8585
rect 44640 8576 44692 8628
rect 46204 8576 46256 8628
rect 48044 8576 48096 8628
rect 48228 8576 48280 8628
rect 50896 8576 50948 8628
rect 40500 8551 40552 8560
rect 33416 8440 33468 8492
rect 34244 8483 34296 8492
rect 34244 8449 34253 8483
rect 34253 8449 34287 8483
rect 34287 8449 34296 8483
rect 34244 8440 34296 8449
rect 34520 8483 34572 8492
rect 34520 8449 34554 8483
rect 34554 8449 34572 8483
rect 34520 8440 34572 8449
rect 35992 8440 36044 8492
rect 36452 8440 36504 8492
rect 38384 8483 38436 8492
rect 38384 8449 38402 8483
rect 38402 8449 38436 8483
rect 38384 8440 38436 8449
rect 25872 8372 25924 8424
rect 27620 8372 27672 8424
rect 19248 8304 19300 8356
rect 26700 8347 26752 8356
rect 26700 8313 26709 8347
rect 26709 8313 26743 8347
rect 26743 8313 26752 8347
rect 26700 8304 26752 8313
rect 29368 8372 29420 8424
rect 31852 8372 31904 8424
rect 32404 8372 32456 8424
rect 40500 8517 40509 8551
rect 40509 8517 40543 8551
rect 40543 8517 40552 8551
rect 40500 8508 40552 8517
rect 45376 8508 45428 8560
rect 50160 8508 50212 8560
rect 29460 8304 29512 8356
rect 31392 8304 31444 8356
rect 32128 8304 32180 8356
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 12992 8236 13044 8288
rect 17316 8279 17368 8288
rect 17316 8245 17325 8279
rect 17325 8245 17359 8279
rect 17359 8245 17368 8279
rect 17316 8236 17368 8245
rect 19432 8236 19484 8288
rect 21640 8279 21692 8288
rect 21640 8245 21649 8279
rect 21649 8245 21683 8279
rect 21683 8245 21692 8279
rect 21640 8236 21692 8245
rect 24032 8236 24084 8288
rect 39672 8483 39724 8492
rect 39672 8449 39681 8483
rect 39681 8449 39715 8483
rect 39715 8449 39724 8483
rect 39672 8440 39724 8449
rect 40408 8440 40460 8492
rect 43536 8440 43588 8492
rect 40224 8415 40276 8424
rect 40224 8381 40233 8415
rect 40233 8381 40267 8415
rect 40267 8381 40276 8415
rect 40224 8372 40276 8381
rect 36084 8236 36136 8288
rect 36728 8236 36780 8288
rect 37740 8236 37792 8288
rect 38292 8236 38344 8288
rect 41420 8415 41472 8424
rect 41420 8381 41429 8415
rect 41429 8381 41463 8415
rect 41463 8381 41472 8415
rect 41420 8372 41472 8381
rect 42248 8415 42300 8424
rect 42248 8381 42257 8415
rect 42257 8381 42291 8415
rect 42291 8381 42300 8415
rect 42248 8372 42300 8381
rect 42524 8372 42576 8424
rect 45560 8415 45612 8424
rect 45560 8381 45569 8415
rect 45569 8381 45603 8415
rect 45603 8381 45612 8415
rect 45560 8372 45612 8381
rect 47952 8483 48004 8492
rect 47952 8449 47961 8483
rect 47961 8449 47995 8483
rect 47995 8449 48004 8483
rect 47952 8440 48004 8449
rect 49056 8483 49108 8492
rect 49056 8449 49065 8483
rect 49065 8449 49099 8483
rect 49099 8449 49108 8483
rect 49056 8440 49108 8449
rect 49332 8483 49384 8492
rect 49332 8449 49341 8483
rect 49341 8449 49375 8483
rect 49375 8449 49384 8483
rect 49332 8440 49384 8449
rect 51172 8619 51224 8628
rect 51172 8585 51181 8619
rect 51181 8585 51215 8619
rect 51215 8585 51224 8619
rect 51172 8576 51224 8585
rect 52920 8576 52972 8628
rect 55220 8576 55272 8628
rect 47768 8415 47820 8424
rect 47768 8381 47777 8415
rect 47777 8381 47811 8415
rect 47811 8381 47820 8415
rect 47768 8372 47820 8381
rect 49240 8415 49292 8424
rect 49240 8381 49258 8415
rect 49258 8381 49292 8415
rect 49240 8372 49292 8381
rect 49608 8415 49660 8424
rect 49608 8381 49617 8415
rect 49617 8381 49651 8415
rect 49651 8381 49660 8415
rect 49608 8372 49660 8381
rect 49884 8372 49936 8424
rect 41512 8304 41564 8356
rect 40868 8279 40920 8288
rect 40868 8245 40877 8279
rect 40877 8245 40911 8279
rect 40911 8245 40920 8279
rect 40868 8236 40920 8245
rect 42156 8236 42208 8288
rect 42340 8236 42392 8288
rect 45376 8236 45428 8288
rect 50252 8415 50304 8424
rect 50252 8381 50261 8415
rect 50261 8381 50295 8415
rect 50295 8381 50304 8415
rect 50252 8372 50304 8381
rect 52828 8440 52880 8492
rect 57796 8576 57848 8628
rect 54852 8483 54904 8492
rect 54852 8449 54861 8483
rect 54861 8449 54895 8483
rect 54895 8449 54904 8483
rect 54852 8440 54904 8449
rect 56324 8440 56376 8492
rect 48320 8279 48372 8288
rect 48320 8245 48329 8279
rect 48329 8245 48363 8279
rect 48363 8245 48372 8279
rect 48320 8236 48372 8245
rect 50160 8304 50212 8356
rect 51264 8304 51316 8356
rect 54668 8372 54720 8424
rect 55128 8415 55180 8424
rect 55128 8381 55137 8415
rect 55137 8381 55171 8415
rect 55171 8381 55180 8415
rect 55128 8372 55180 8381
rect 55312 8372 55364 8424
rect 56140 8372 56192 8424
rect 51908 8279 51960 8288
rect 51908 8245 51917 8279
rect 51917 8245 51951 8279
rect 51951 8245 51960 8279
rect 51908 8236 51960 8245
rect 54024 8236 54076 8288
rect 57704 8236 57756 8288
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 22616 8134 22668 8186
rect 22680 8134 22732 8186
rect 22744 8134 22796 8186
rect 22808 8134 22860 8186
rect 22872 8134 22924 8186
rect 37060 8134 37112 8186
rect 37124 8134 37176 8186
rect 37188 8134 37240 8186
rect 37252 8134 37304 8186
rect 37316 8134 37368 8186
rect 51504 8134 51556 8186
rect 51568 8134 51620 8186
rect 51632 8134 51684 8186
rect 51696 8134 51748 8186
rect 51760 8134 51812 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 3976 8032 4028 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6276 8032 6328 8084
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 3700 7828 3752 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4344 7828 4396 7880
rect 7748 7964 7800 8016
rect 5816 7828 5868 7880
rect 6092 7828 6144 7880
rect 8760 8032 8812 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10784 8032 10836 8084
rect 11796 8032 11848 8084
rect 12164 8032 12216 8084
rect 8852 7964 8904 8016
rect 13360 8032 13412 8084
rect 17960 8075 18012 8084
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 4712 7760 4764 7812
rect 8300 7828 8352 7880
rect 8484 7828 8536 7880
rect 8668 7828 8720 7880
rect 9496 7828 9548 7880
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 13084 7896 13136 7948
rect 14832 7896 14884 7948
rect 15108 7896 15160 7948
rect 15200 7939 15252 7948
rect 15200 7905 15209 7939
rect 15209 7905 15243 7939
rect 15243 7905 15252 7939
rect 15200 7896 15252 7905
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 19340 7964 19392 8016
rect 22284 7964 22336 8016
rect 24124 7964 24176 8016
rect 25320 7964 25372 8016
rect 25780 8007 25832 8016
rect 25780 7973 25789 8007
rect 25789 7973 25823 8007
rect 25823 7973 25832 8007
rect 25780 7964 25832 7973
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 29368 7939 29420 7948
rect 29368 7905 29377 7939
rect 29377 7905 29411 7939
rect 29411 7905 29420 7939
rect 29368 7896 29420 7905
rect 4068 7692 4120 7744
rect 5448 7692 5500 7744
rect 7380 7692 7432 7744
rect 7472 7692 7524 7744
rect 9588 7803 9640 7812
rect 9588 7769 9597 7803
rect 9597 7769 9631 7803
rect 9631 7769 9640 7803
rect 9588 7760 9640 7769
rect 12716 7828 12768 7880
rect 17776 7828 17828 7880
rect 20536 7828 20588 7880
rect 20812 7828 20864 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 23572 7871 23624 7880
rect 23572 7837 23581 7871
rect 23581 7837 23615 7871
rect 23615 7837 23624 7871
rect 23572 7828 23624 7837
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 26700 7828 26752 7880
rect 18144 7760 18196 7812
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 19156 7692 19208 7744
rect 20628 7692 20680 7744
rect 23020 7735 23072 7744
rect 23020 7701 23029 7735
rect 23029 7701 23063 7735
rect 23063 7701 23072 7735
rect 23020 7692 23072 7701
rect 24032 7735 24084 7744
rect 24032 7701 24041 7735
rect 24041 7701 24075 7735
rect 24075 7701 24084 7735
rect 24032 7692 24084 7701
rect 25964 7735 26016 7744
rect 25964 7701 25973 7735
rect 25973 7701 26007 7735
rect 26007 7701 26016 7735
rect 25964 7692 26016 7701
rect 27620 7692 27672 7744
rect 28724 7735 28776 7744
rect 28724 7701 28733 7735
rect 28733 7701 28767 7735
rect 28767 7701 28776 7735
rect 28724 7692 28776 7701
rect 29460 7692 29512 7744
rect 33416 8032 33468 8084
rect 38476 8032 38528 8084
rect 41696 8032 41748 8084
rect 42524 8032 42576 8084
rect 45560 8032 45612 8084
rect 47952 8075 48004 8084
rect 47952 8041 47961 8075
rect 47961 8041 47995 8075
rect 47995 8041 48004 8075
rect 47952 8032 48004 8041
rect 50252 8032 50304 8084
rect 31760 7939 31812 7948
rect 31760 7905 31769 7939
rect 31769 7905 31803 7939
rect 31803 7905 31812 7939
rect 31760 7896 31812 7905
rect 32220 7939 32272 7948
rect 32220 7905 32229 7939
rect 32229 7905 32263 7939
rect 32263 7905 32272 7939
rect 32220 7896 32272 7905
rect 32496 7896 32548 7948
rect 32680 7896 32732 7948
rect 35716 7896 35768 7948
rect 35992 7896 36044 7948
rect 36452 7896 36504 7948
rect 32864 7828 32916 7880
rect 36912 7939 36964 7948
rect 36912 7905 36921 7939
rect 36921 7905 36955 7939
rect 36955 7905 36964 7939
rect 36912 7896 36964 7905
rect 37188 7939 37240 7948
rect 37188 7905 37197 7939
rect 37197 7905 37231 7939
rect 37231 7905 37240 7939
rect 37188 7896 37240 7905
rect 37648 7939 37700 7948
rect 37648 7905 37657 7939
rect 37657 7905 37691 7939
rect 37691 7905 37700 7939
rect 37648 7896 37700 7905
rect 37740 7896 37792 7948
rect 30472 7760 30524 7812
rect 31852 7760 31904 7812
rect 36728 7828 36780 7880
rect 38016 7896 38068 7948
rect 44824 7964 44876 8016
rect 45192 7964 45244 8016
rect 50160 8007 50212 8016
rect 50160 7973 50169 8007
rect 50169 7973 50203 8007
rect 50203 7973 50212 8007
rect 50160 7964 50212 7973
rect 44640 7896 44692 7948
rect 52828 8032 52880 8084
rect 55128 8032 55180 8084
rect 54944 8007 54996 8016
rect 40500 7828 40552 7880
rect 41972 7828 42024 7880
rect 42156 7871 42208 7880
rect 42156 7837 42190 7871
rect 42190 7837 42208 7871
rect 42156 7828 42208 7837
rect 38292 7803 38344 7812
rect 38292 7769 38301 7803
rect 38301 7769 38335 7803
rect 38335 7769 38344 7803
rect 38292 7760 38344 7769
rect 40316 7760 40368 7812
rect 40868 7760 40920 7812
rect 32312 7692 32364 7744
rect 34888 7735 34940 7744
rect 34888 7701 34897 7735
rect 34897 7701 34931 7735
rect 34931 7701 34940 7735
rect 34888 7692 34940 7701
rect 35256 7735 35308 7744
rect 35256 7701 35265 7735
rect 35265 7701 35299 7735
rect 35299 7701 35308 7735
rect 35256 7692 35308 7701
rect 37648 7692 37700 7744
rect 37924 7735 37976 7744
rect 37924 7701 37933 7735
rect 37933 7701 37967 7735
rect 37967 7701 37976 7735
rect 37924 7692 37976 7701
rect 39028 7692 39080 7744
rect 46480 7760 46532 7812
rect 47584 7760 47636 7812
rect 43260 7735 43312 7744
rect 43260 7701 43269 7735
rect 43269 7701 43303 7735
rect 43303 7701 43312 7735
rect 43260 7692 43312 7701
rect 43996 7692 44048 7744
rect 44180 7692 44232 7744
rect 45468 7692 45520 7744
rect 51908 7828 51960 7880
rect 54944 7973 54953 8007
rect 54953 7973 54987 8007
rect 54987 7973 54996 8007
rect 54944 7964 54996 7973
rect 53932 7896 53984 7948
rect 55220 7896 55272 7948
rect 55864 7939 55916 7948
rect 55864 7905 55873 7939
rect 55873 7905 55907 7939
rect 55907 7905 55916 7939
rect 55864 7896 55916 7905
rect 57704 7939 57756 7948
rect 57704 7905 57713 7939
rect 57713 7905 57747 7939
rect 57747 7905 57756 7939
rect 57704 7896 57756 7905
rect 58072 7896 58124 7948
rect 54484 7828 54536 7880
rect 48596 7760 48648 7812
rect 49240 7760 49292 7812
rect 49884 7735 49936 7744
rect 49884 7701 49893 7735
rect 49893 7701 49927 7735
rect 49927 7701 49936 7735
rect 49884 7692 49936 7701
rect 52000 7735 52052 7744
rect 52000 7701 52009 7735
rect 52009 7701 52043 7735
rect 52043 7701 52052 7735
rect 52000 7692 52052 7701
rect 55312 7735 55364 7744
rect 55312 7701 55321 7735
rect 55321 7701 55355 7735
rect 55355 7701 55364 7735
rect 55312 7692 55364 7701
rect 56140 7692 56192 7744
rect 56508 7692 56560 7744
rect 15394 7590 15446 7642
rect 15458 7590 15510 7642
rect 15522 7590 15574 7642
rect 15586 7590 15638 7642
rect 15650 7590 15702 7642
rect 29838 7590 29890 7642
rect 29902 7590 29954 7642
rect 29966 7590 30018 7642
rect 30030 7590 30082 7642
rect 30094 7590 30146 7642
rect 44282 7590 44334 7642
rect 44346 7590 44398 7642
rect 44410 7590 44462 7642
rect 44474 7590 44526 7642
rect 44538 7590 44590 7642
rect 58726 7590 58778 7642
rect 58790 7590 58842 7642
rect 58854 7590 58906 7642
rect 58918 7590 58970 7642
rect 58982 7590 59034 7642
rect 3424 7420 3476 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 4528 7463 4580 7472
rect 4528 7429 4537 7463
rect 4537 7429 4571 7463
rect 4571 7429 4580 7463
rect 4528 7420 4580 7429
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4712 7352 4764 7404
rect 4896 7284 4948 7336
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 4344 7216 4396 7268
rect 6000 7488 6052 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 9588 7488 9640 7540
rect 11244 7488 11296 7540
rect 14280 7488 14332 7540
rect 14832 7488 14884 7540
rect 14924 7488 14976 7540
rect 16580 7488 16632 7540
rect 20628 7488 20680 7540
rect 8668 7420 8720 7472
rect 7748 7352 7800 7404
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 7288 7284 7340 7336
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 8300 7284 8352 7336
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 3700 7148 3752 7200
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 15844 7352 15896 7404
rect 16580 7352 16632 7404
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17776 7352 17828 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 20812 7463 20864 7472
rect 20812 7429 20821 7463
rect 20821 7429 20855 7463
rect 20855 7429 20864 7463
rect 20812 7420 20864 7429
rect 21364 7420 21416 7472
rect 21640 7420 21692 7472
rect 24124 7420 24176 7472
rect 24676 7463 24728 7472
rect 24676 7429 24685 7463
rect 24685 7429 24719 7463
rect 24719 7429 24728 7463
rect 24676 7420 24728 7429
rect 23020 7352 23072 7404
rect 24032 7352 24084 7404
rect 25964 7488 26016 7540
rect 28448 7531 28500 7540
rect 28448 7497 28457 7531
rect 28457 7497 28491 7531
rect 28491 7497 28500 7531
rect 28448 7488 28500 7497
rect 28724 7488 28776 7540
rect 29644 7488 29696 7540
rect 30564 7488 30616 7540
rect 31576 7488 31628 7540
rect 32404 7531 32456 7540
rect 32404 7497 32413 7531
rect 32413 7497 32447 7531
rect 32447 7497 32456 7531
rect 32404 7488 32456 7497
rect 34244 7531 34296 7540
rect 34244 7497 34253 7531
rect 34253 7497 34287 7531
rect 34287 7497 34296 7531
rect 34244 7488 34296 7497
rect 34520 7488 34572 7540
rect 35256 7488 35308 7540
rect 35808 7488 35860 7540
rect 36452 7488 36504 7540
rect 36820 7531 36872 7540
rect 36820 7497 36829 7531
rect 36829 7497 36863 7531
rect 36863 7497 36872 7531
rect 36820 7488 36872 7497
rect 38384 7531 38436 7540
rect 38384 7497 38393 7531
rect 38393 7497 38427 7531
rect 38427 7497 38436 7531
rect 38384 7488 38436 7497
rect 38476 7488 38528 7540
rect 37740 7420 37792 7472
rect 38108 7420 38160 7472
rect 40684 7420 40736 7472
rect 28816 7352 28868 7404
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 15108 7284 15160 7336
rect 18236 7284 18288 7336
rect 18972 7284 19024 7336
rect 29736 7352 29788 7404
rect 7380 7148 7432 7200
rect 7656 7148 7708 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8484 7148 8536 7200
rect 8668 7148 8720 7200
rect 12440 7148 12492 7200
rect 14096 7148 14148 7200
rect 15200 7148 15252 7200
rect 16028 7148 16080 7200
rect 16672 7148 16724 7200
rect 24860 7216 24912 7268
rect 26608 7259 26660 7268
rect 26608 7225 26617 7259
rect 26617 7225 26651 7259
rect 26651 7225 26660 7259
rect 26608 7216 26660 7225
rect 30196 7216 30248 7268
rect 17960 7148 18012 7200
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 21272 7148 21324 7200
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 26792 7148 26844 7200
rect 27620 7148 27672 7200
rect 29460 7148 29512 7200
rect 30380 7191 30432 7200
rect 30380 7157 30389 7191
rect 30389 7157 30423 7191
rect 30423 7157 30432 7191
rect 30380 7148 30432 7157
rect 30564 7191 30616 7200
rect 30564 7157 30573 7191
rect 30573 7157 30607 7191
rect 30607 7157 30616 7191
rect 30564 7148 30616 7157
rect 31116 7327 31168 7336
rect 31116 7293 31125 7327
rect 31125 7293 31159 7327
rect 31159 7293 31168 7327
rect 31116 7284 31168 7293
rect 33416 7327 33468 7336
rect 33416 7293 33425 7327
rect 33425 7293 33459 7327
rect 33459 7293 33468 7327
rect 33416 7284 33468 7293
rect 34888 7352 34940 7404
rect 35624 7352 35676 7404
rect 35900 7284 35952 7336
rect 36084 7327 36136 7336
rect 36084 7293 36093 7327
rect 36093 7293 36127 7327
rect 36127 7293 36136 7327
rect 36084 7284 36136 7293
rect 36544 7352 36596 7404
rect 37188 7352 37240 7404
rect 37924 7352 37976 7404
rect 38476 7352 38528 7404
rect 40408 7352 40460 7404
rect 36728 7284 36780 7336
rect 38016 7284 38068 7336
rect 38200 7284 38252 7336
rect 38384 7284 38436 7336
rect 40132 7327 40184 7336
rect 40132 7293 40141 7327
rect 40141 7293 40175 7327
rect 40175 7293 40184 7327
rect 40132 7284 40184 7293
rect 40500 7327 40552 7336
rect 40500 7293 40509 7327
rect 40509 7293 40543 7327
rect 40543 7293 40552 7327
rect 40500 7284 40552 7293
rect 41420 7488 41472 7540
rect 41512 7531 41564 7540
rect 41512 7497 41521 7531
rect 41521 7497 41555 7531
rect 41555 7497 41564 7531
rect 41512 7488 41564 7497
rect 42248 7488 42300 7540
rect 43536 7488 43588 7540
rect 46756 7531 46808 7540
rect 46756 7497 46765 7531
rect 46765 7497 46799 7531
rect 46799 7497 46808 7531
rect 46756 7488 46808 7497
rect 47584 7531 47636 7540
rect 47584 7497 47593 7531
rect 47593 7497 47627 7531
rect 47627 7497 47636 7531
rect 47584 7488 47636 7497
rect 48596 7531 48648 7540
rect 48596 7497 48605 7531
rect 48605 7497 48639 7531
rect 48639 7497 48648 7531
rect 48596 7488 48648 7497
rect 49148 7488 49200 7540
rect 52000 7488 52052 7540
rect 53472 7531 53524 7540
rect 53472 7497 53481 7531
rect 53481 7497 53515 7531
rect 53515 7497 53524 7531
rect 53472 7488 53524 7497
rect 54024 7488 54076 7540
rect 54116 7531 54168 7540
rect 54116 7497 54125 7531
rect 54125 7497 54159 7531
rect 54159 7497 54168 7531
rect 54116 7488 54168 7497
rect 56784 7488 56836 7540
rect 57612 7531 57664 7540
rect 57612 7497 57621 7531
rect 57621 7497 57655 7531
rect 57655 7497 57664 7531
rect 57612 7488 57664 7497
rect 57888 7531 57940 7540
rect 57888 7497 57897 7531
rect 57897 7497 57931 7531
rect 57931 7497 57940 7531
rect 57888 7488 57940 7497
rect 41972 7420 42024 7472
rect 43996 7420 44048 7472
rect 44088 7420 44140 7472
rect 52552 7420 52604 7472
rect 55588 7420 55640 7472
rect 41420 7395 41472 7404
rect 41420 7361 41429 7395
rect 41429 7361 41463 7395
rect 41463 7361 41472 7395
rect 41420 7352 41472 7361
rect 42708 7352 42760 7404
rect 41696 7284 41748 7336
rect 43444 7284 43496 7336
rect 45376 7352 45428 7404
rect 48320 7352 48372 7404
rect 48688 7352 48740 7404
rect 49884 7352 49936 7404
rect 50252 7352 50304 7404
rect 48780 7284 48832 7336
rect 52184 7352 52236 7404
rect 55128 7352 55180 7404
rect 58072 7420 58124 7472
rect 57612 7352 57664 7404
rect 55864 7284 55916 7336
rect 56508 7284 56560 7336
rect 32312 7216 32364 7268
rect 32680 7216 32732 7268
rect 39856 7216 39908 7268
rect 44916 7216 44968 7268
rect 32496 7148 32548 7200
rect 33416 7148 33468 7200
rect 35624 7148 35676 7200
rect 36452 7191 36504 7200
rect 36452 7157 36461 7191
rect 36461 7157 36495 7191
rect 36495 7157 36504 7191
rect 36452 7148 36504 7157
rect 38476 7148 38528 7200
rect 38752 7148 38804 7200
rect 39028 7191 39080 7200
rect 39028 7157 39037 7191
rect 39037 7157 39071 7191
rect 39071 7157 39080 7191
rect 39028 7148 39080 7157
rect 44824 7148 44876 7200
rect 45192 7148 45244 7200
rect 46480 7191 46532 7200
rect 46480 7157 46489 7191
rect 46489 7157 46523 7191
rect 46523 7157 46532 7191
rect 46480 7148 46532 7157
rect 47124 7148 47176 7200
rect 58256 7216 58308 7268
rect 52000 7191 52052 7200
rect 52000 7157 52009 7191
rect 52009 7157 52043 7191
rect 52043 7157 52052 7191
rect 52000 7148 52052 7157
rect 52644 7148 52696 7200
rect 52920 7191 52972 7200
rect 52920 7157 52929 7191
rect 52929 7157 52963 7191
rect 52963 7157 52972 7191
rect 52920 7148 52972 7157
rect 54760 7148 54812 7200
rect 55496 7191 55548 7200
rect 55496 7157 55505 7191
rect 55505 7157 55539 7191
rect 55539 7157 55548 7191
rect 55496 7148 55548 7157
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 22616 7046 22668 7098
rect 22680 7046 22732 7098
rect 22744 7046 22796 7098
rect 22808 7046 22860 7098
rect 22872 7046 22924 7098
rect 37060 7046 37112 7098
rect 37124 7046 37176 7098
rect 37188 7046 37240 7098
rect 37252 7046 37304 7098
rect 37316 7046 37368 7098
rect 51504 7046 51556 7098
rect 51568 7046 51620 7098
rect 51632 7046 51684 7098
rect 51696 7046 51748 7098
rect 51760 7046 51812 7098
rect 3424 6944 3476 6996
rect 12256 6944 12308 6996
rect 3332 6851 3384 6860
rect 3332 6817 3341 6851
rect 3341 6817 3375 6851
rect 3375 6817 3384 6851
rect 3332 6808 3384 6817
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5080 6876 5132 6928
rect 12348 6876 12400 6928
rect 13820 6944 13872 6996
rect 20444 6944 20496 6996
rect 13912 6876 13964 6928
rect 21364 6919 21416 6928
rect 6460 6808 6512 6860
rect 7104 6808 7156 6860
rect 7564 6808 7616 6860
rect 7748 6808 7800 6860
rect 4068 6672 4120 6724
rect 3700 6604 3752 6656
rect 3976 6604 4028 6656
rect 4896 6647 4948 6656
rect 4896 6613 4905 6647
rect 4905 6613 4939 6647
rect 4939 6613 4948 6647
rect 4896 6604 4948 6613
rect 6368 6604 6420 6656
rect 6828 6604 6880 6656
rect 7104 6604 7156 6656
rect 8576 6808 8628 6860
rect 8208 6740 8260 6792
rect 9128 6740 9180 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 12440 6740 12492 6792
rect 9036 6672 9088 6724
rect 9128 6604 9180 6656
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 11060 6672 11112 6724
rect 12256 6715 12308 6724
rect 12256 6681 12265 6715
rect 12265 6681 12299 6715
rect 12299 6681 12308 6715
rect 12256 6672 12308 6681
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 11796 6604 11848 6656
rect 12164 6604 12216 6656
rect 14280 6604 14332 6656
rect 14740 6740 14792 6792
rect 16672 6740 16724 6792
rect 17960 6808 18012 6860
rect 19248 6851 19300 6860
rect 19248 6817 19257 6851
rect 19257 6817 19291 6851
rect 19291 6817 19300 6851
rect 19248 6808 19300 6817
rect 19616 6808 19668 6860
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 21364 6885 21373 6919
rect 21373 6885 21407 6919
rect 21407 6885 21416 6919
rect 21364 6876 21416 6885
rect 20260 6851 20312 6860
rect 20260 6817 20294 6851
rect 20294 6817 20312 6851
rect 20260 6808 20312 6817
rect 23572 6944 23624 6996
rect 24676 6944 24728 6996
rect 23664 6808 23716 6860
rect 23756 6808 23808 6860
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 15936 6604 15988 6656
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 17776 6672 17828 6724
rect 17316 6604 17368 6656
rect 19340 6672 19392 6724
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 24308 6808 24360 6860
rect 24860 6808 24912 6860
rect 25780 6944 25832 6996
rect 26516 6944 26568 6996
rect 30380 6944 30432 6996
rect 31116 6944 31168 6996
rect 25688 6808 25740 6860
rect 26608 6808 26660 6860
rect 26792 6851 26844 6860
rect 26792 6817 26801 6851
rect 26801 6817 26835 6851
rect 26835 6817 26844 6851
rect 26792 6808 26844 6817
rect 30196 6876 30248 6928
rect 34980 6919 35032 6928
rect 34980 6885 34989 6919
rect 34989 6885 35023 6919
rect 35023 6885 35032 6919
rect 34980 6876 35032 6885
rect 35716 6876 35768 6928
rect 35900 6876 35952 6928
rect 36360 6876 36412 6928
rect 36820 6876 36872 6928
rect 37188 6876 37240 6928
rect 27804 6851 27856 6860
rect 27804 6817 27813 6851
rect 27813 6817 27847 6851
rect 27847 6817 27856 6851
rect 27804 6808 27856 6817
rect 29000 6808 29052 6860
rect 30472 6851 30524 6860
rect 30472 6817 30481 6851
rect 30481 6817 30515 6851
rect 30515 6817 30524 6851
rect 30472 6808 30524 6817
rect 30564 6808 30616 6860
rect 21916 6740 21968 6749
rect 25044 6783 25096 6792
rect 25044 6749 25053 6783
rect 25053 6749 25087 6783
rect 25087 6749 25096 6783
rect 25044 6740 25096 6749
rect 25136 6740 25188 6792
rect 26056 6783 26108 6792
rect 26056 6749 26065 6783
rect 26065 6749 26099 6783
rect 26099 6749 26108 6783
rect 26056 6740 26108 6749
rect 22468 6672 22520 6724
rect 19708 6604 19760 6656
rect 20904 6604 20956 6656
rect 23940 6604 23992 6656
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 25136 6604 25188 6656
rect 27160 6647 27212 6656
rect 27160 6613 27169 6647
rect 27169 6613 27203 6647
rect 27203 6613 27212 6647
rect 27160 6604 27212 6613
rect 28816 6604 28868 6656
rect 32496 6740 32548 6792
rect 35624 6808 35676 6860
rect 33600 6740 33652 6792
rect 33416 6672 33468 6724
rect 33692 6715 33744 6724
rect 33692 6681 33701 6715
rect 33701 6681 33735 6715
rect 33735 6681 33744 6715
rect 33692 6672 33744 6681
rect 35992 6783 36044 6792
rect 35992 6749 36001 6783
rect 36001 6749 36035 6783
rect 36035 6749 36044 6783
rect 35992 6740 36044 6749
rect 36268 6851 36320 6860
rect 36268 6817 36277 6851
rect 36277 6817 36311 6851
rect 36311 6817 36320 6851
rect 36268 6808 36320 6817
rect 41420 6944 41472 6996
rect 42708 6944 42760 6996
rect 45468 6987 45520 6996
rect 45468 6953 45477 6987
rect 45477 6953 45511 6987
rect 45511 6953 45520 6987
rect 45468 6944 45520 6953
rect 40408 6851 40460 6860
rect 40408 6817 40417 6851
rect 40417 6817 40451 6851
rect 40451 6817 40460 6851
rect 40408 6808 40460 6817
rect 43996 6919 44048 6928
rect 43996 6885 44005 6919
rect 44005 6885 44039 6919
rect 44039 6885 44048 6919
rect 43996 6876 44048 6885
rect 45192 6876 45244 6928
rect 54392 6944 54444 6996
rect 55588 6987 55640 6996
rect 55588 6953 55597 6987
rect 55597 6953 55631 6987
rect 55631 6953 55640 6987
rect 55588 6944 55640 6953
rect 53196 6876 53248 6928
rect 35256 6672 35308 6724
rect 37556 6672 37608 6724
rect 38660 6715 38712 6724
rect 38660 6681 38669 6715
rect 38669 6681 38703 6715
rect 38703 6681 38712 6715
rect 38660 6672 38712 6681
rect 31024 6604 31076 6656
rect 31760 6604 31812 6656
rect 33508 6604 33560 6656
rect 35440 6647 35492 6656
rect 35440 6613 35449 6647
rect 35449 6613 35483 6647
rect 35483 6613 35492 6647
rect 35440 6604 35492 6613
rect 36084 6604 36136 6656
rect 38292 6604 38344 6656
rect 38568 6604 38620 6656
rect 39120 6604 39172 6656
rect 40132 6740 40184 6792
rect 42524 6808 42576 6860
rect 42616 6851 42668 6860
rect 42616 6817 42625 6851
rect 42625 6817 42659 6851
rect 42659 6817 42668 6851
rect 42616 6808 42668 6817
rect 43260 6851 43312 6860
rect 43260 6817 43269 6851
rect 43269 6817 43303 6851
rect 43303 6817 43312 6851
rect 43260 6808 43312 6817
rect 46664 6851 46716 6860
rect 46664 6817 46673 6851
rect 46673 6817 46707 6851
rect 46707 6817 46716 6851
rect 46664 6808 46716 6817
rect 47860 6808 47912 6860
rect 48504 6808 48556 6860
rect 42064 6783 42116 6792
rect 42064 6749 42073 6783
rect 42073 6749 42107 6783
rect 42107 6749 42116 6783
rect 42064 6740 42116 6749
rect 43076 6783 43128 6792
rect 43076 6749 43085 6783
rect 43085 6749 43119 6783
rect 43119 6749 43128 6783
rect 43076 6740 43128 6749
rect 45652 6740 45704 6792
rect 46756 6740 46808 6792
rect 47308 6740 47360 6792
rect 52460 6808 52512 6860
rect 52644 6808 52696 6860
rect 45836 6672 45888 6724
rect 46480 6672 46532 6724
rect 46664 6672 46716 6724
rect 51908 6783 51960 6792
rect 51908 6749 51917 6783
rect 51917 6749 51951 6783
rect 51951 6749 51960 6783
rect 51908 6740 51960 6749
rect 55496 6808 55548 6860
rect 56600 6876 56652 6928
rect 56784 6851 56836 6860
rect 56784 6817 56793 6851
rect 56793 6817 56827 6851
rect 56827 6817 56836 6851
rect 56784 6808 56836 6817
rect 57888 6808 57940 6860
rect 41236 6604 41288 6656
rect 42800 6604 42852 6656
rect 43628 6647 43680 6656
rect 43628 6613 43637 6647
rect 43637 6613 43671 6647
rect 43671 6613 43680 6647
rect 43628 6604 43680 6613
rect 44824 6604 44876 6656
rect 45744 6647 45796 6656
rect 45744 6613 45753 6647
rect 45753 6613 45787 6647
rect 45787 6613 45796 6647
rect 45744 6604 45796 6613
rect 47492 6604 47544 6656
rect 49884 6672 49936 6724
rect 48044 6604 48096 6656
rect 48320 6604 48372 6656
rect 49056 6604 49108 6656
rect 49792 6604 49844 6656
rect 50252 6604 50304 6656
rect 51172 6672 51224 6724
rect 50804 6604 50856 6656
rect 52000 6604 52052 6656
rect 52276 6604 52328 6656
rect 53104 6604 53156 6656
rect 54116 6604 54168 6656
rect 55956 6604 56008 6656
rect 56784 6604 56836 6656
rect 56968 6647 57020 6656
rect 56968 6613 56977 6647
rect 56977 6613 57011 6647
rect 57011 6613 57020 6647
rect 56968 6604 57020 6613
rect 57980 6672 58032 6724
rect 57520 6647 57572 6656
rect 57520 6613 57529 6647
rect 57529 6613 57563 6647
rect 57563 6613 57572 6647
rect 57520 6604 57572 6613
rect 58348 6647 58400 6656
rect 58348 6613 58357 6647
rect 58357 6613 58391 6647
rect 58391 6613 58400 6647
rect 58348 6604 58400 6613
rect 15394 6502 15446 6554
rect 15458 6502 15510 6554
rect 15522 6502 15574 6554
rect 15586 6502 15638 6554
rect 15650 6502 15702 6554
rect 29838 6502 29890 6554
rect 29902 6502 29954 6554
rect 29966 6502 30018 6554
rect 30030 6502 30082 6554
rect 30094 6502 30146 6554
rect 44282 6502 44334 6554
rect 44346 6502 44398 6554
rect 44410 6502 44462 6554
rect 44474 6502 44526 6554
rect 44538 6502 44590 6554
rect 58726 6502 58778 6554
rect 58790 6502 58842 6554
rect 58854 6502 58906 6554
rect 58918 6502 58970 6554
rect 58982 6502 59034 6554
rect 7748 6400 7800 6452
rect 8208 6400 8260 6452
rect 8576 6400 8628 6452
rect 10048 6400 10100 6452
rect 11612 6400 11664 6452
rect 13912 6400 13964 6452
rect 14280 6400 14332 6452
rect 6000 6375 6052 6384
rect 6000 6341 6009 6375
rect 6009 6341 6043 6375
rect 6043 6341 6052 6375
rect 6000 6332 6052 6341
rect 7564 6332 7616 6384
rect 10232 6375 10284 6384
rect 5448 6264 5500 6316
rect 7380 6264 7432 6316
rect 9036 6264 9088 6316
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 3976 6128 4028 6180
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 5724 6196 5776 6248
rect 7012 6196 7064 6248
rect 9588 6264 9640 6316
rect 10232 6341 10266 6375
rect 10266 6341 10284 6375
rect 10232 6332 10284 6341
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 11336 6171 11388 6180
rect 11336 6137 11345 6171
rect 11345 6137 11379 6171
rect 11379 6137 11388 6171
rect 11336 6128 11388 6137
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 3240 6060 3292 6112
rect 3516 6103 3568 6112
rect 3516 6069 3525 6103
rect 3525 6069 3559 6103
rect 3559 6069 3568 6103
rect 3516 6060 3568 6069
rect 4436 6103 4488 6112
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 7196 6060 7248 6112
rect 8024 6060 8076 6112
rect 11704 6060 11756 6112
rect 14740 6400 14792 6452
rect 16764 6400 16816 6452
rect 17316 6400 17368 6452
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 18788 6400 18840 6452
rect 19616 6400 19668 6452
rect 19708 6443 19760 6452
rect 19708 6409 19717 6443
rect 19717 6409 19751 6443
rect 19751 6409 19760 6443
rect 19708 6400 19760 6409
rect 16672 6307 16724 6316
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 18420 6264 18472 6316
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 13636 6171 13688 6180
rect 13636 6137 13645 6171
rect 13645 6137 13679 6171
rect 13679 6137 13688 6171
rect 13636 6128 13688 6137
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 19524 6264 19576 6316
rect 19892 6332 19944 6384
rect 22284 6332 22336 6384
rect 20260 6264 20312 6316
rect 20812 6307 20864 6316
rect 20812 6273 20830 6307
rect 20830 6273 20864 6307
rect 20812 6264 20864 6273
rect 21364 6264 21416 6316
rect 25136 6400 25188 6452
rect 26056 6400 26108 6452
rect 23940 6332 23992 6384
rect 25320 6332 25372 6384
rect 37188 6400 37240 6452
rect 24768 6307 24820 6316
rect 24768 6273 24777 6307
rect 24777 6273 24811 6307
rect 24811 6273 24820 6307
rect 24768 6264 24820 6273
rect 26516 6264 26568 6316
rect 27160 6264 27212 6316
rect 28816 6307 28868 6316
rect 28816 6273 28839 6307
rect 28839 6273 28868 6307
rect 28816 6264 28868 6273
rect 31024 6332 31076 6384
rect 21640 6171 21692 6180
rect 21640 6137 21649 6171
rect 21649 6137 21683 6171
rect 21683 6137 21692 6171
rect 21640 6128 21692 6137
rect 23664 6128 23716 6180
rect 21088 6060 21140 6112
rect 21180 6060 21232 6112
rect 23020 6060 23072 6112
rect 25044 6060 25096 6112
rect 27620 6060 27672 6112
rect 30196 6060 30248 6112
rect 31116 6307 31168 6316
rect 31116 6273 31134 6307
rect 31134 6273 31168 6307
rect 31116 6264 31168 6273
rect 31392 6239 31444 6248
rect 31392 6205 31401 6239
rect 31401 6205 31435 6239
rect 31435 6205 31444 6239
rect 31392 6196 31444 6205
rect 32220 6332 32272 6384
rect 33232 6307 33284 6316
rect 35256 6332 35308 6384
rect 35440 6375 35492 6384
rect 35440 6341 35474 6375
rect 35474 6341 35492 6375
rect 35440 6332 35492 6341
rect 35532 6332 35584 6384
rect 36268 6332 36320 6384
rect 33232 6273 33250 6307
rect 33250 6273 33284 6307
rect 33232 6264 33284 6273
rect 34428 6239 34480 6248
rect 34428 6205 34437 6239
rect 34437 6205 34471 6239
rect 34471 6205 34480 6239
rect 36452 6264 36504 6316
rect 37464 6264 37516 6316
rect 41236 6400 41288 6452
rect 42064 6400 42116 6452
rect 34428 6196 34480 6205
rect 36176 6196 36228 6248
rect 40500 6332 40552 6384
rect 43076 6400 43128 6452
rect 43628 6332 43680 6384
rect 39120 6307 39172 6316
rect 39120 6273 39143 6307
rect 39143 6273 39172 6307
rect 39120 6264 39172 6273
rect 40408 6264 40460 6316
rect 45744 6400 45796 6452
rect 48780 6443 48832 6452
rect 48780 6409 48789 6443
rect 48789 6409 48823 6443
rect 48823 6409 48832 6443
rect 48780 6400 48832 6409
rect 44088 6332 44140 6384
rect 44824 6332 44876 6384
rect 38660 6196 38712 6248
rect 40868 6239 40920 6248
rect 40868 6205 40877 6239
rect 40877 6205 40911 6239
rect 40911 6205 40920 6239
rect 40868 6196 40920 6205
rect 41696 6239 41748 6248
rect 41696 6205 41705 6239
rect 41705 6205 41739 6239
rect 41739 6205 41748 6239
rect 41696 6196 41748 6205
rect 33600 6128 33652 6180
rect 38752 6128 38804 6180
rect 45192 6264 45244 6316
rect 48320 6264 48372 6316
rect 47124 6239 47176 6248
rect 47124 6205 47133 6239
rect 47133 6205 47167 6239
rect 47167 6205 47176 6239
rect 47124 6196 47176 6205
rect 32772 6060 32824 6112
rect 36544 6103 36596 6112
rect 36544 6069 36553 6103
rect 36553 6069 36587 6103
rect 36587 6069 36596 6103
rect 36544 6060 36596 6069
rect 36912 6060 36964 6112
rect 39764 6060 39816 6112
rect 41144 6060 41196 6112
rect 43352 6060 43404 6112
rect 44824 6103 44876 6112
rect 44824 6069 44833 6103
rect 44833 6069 44867 6103
rect 44867 6069 44876 6103
rect 44824 6060 44876 6069
rect 46204 6060 46256 6112
rect 46572 6103 46624 6112
rect 46572 6069 46581 6103
rect 46581 6069 46615 6103
rect 46615 6069 46624 6103
rect 46572 6060 46624 6069
rect 47676 6060 47728 6112
rect 48136 6128 48188 6180
rect 49608 6264 49660 6316
rect 51080 6239 51132 6248
rect 51080 6205 51089 6239
rect 51089 6205 51123 6239
rect 51123 6205 51132 6239
rect 51080 6196 51132 6205
rect 51908 6400 51960 6452
rect 53104 6400 53156 6452
rect 53196 6400 53248 6452
rect 54116 6443 54168 6452
rect 54116 6409 54125 6443
rect 54125 6409 54159 6443
rect 54159 6409 54168 6443
rect 54116 6400 54168 6409
rect 52552 6264 52604 6316
rect 52828 6264 52880 6316
rect 54944 6307 54996 6316
rect 54944 6273 54953 6307
rect 54953 6273 54987 6307
rect 54987 6273 54996 6307
rect 54944 6264 54996 6273
rect 57520 6400 57572 6452
rect 57888 6400 57940 6452
rect 57704 6307 57756 6316
rect 57704 6273 57713 6307
rect 57713 6273 57747 6307
rect 57747 6273 57756 6307
rect 57704 6264 57756 6273
rect 55220 6239 55272 6248
rect 55220 6205 55229 6239
rect 55229 6205 55263 6239
rect 55263 6205 55272 6239
rect 55220 6196 55272 6205
rect 55588 6196 55640 6248
rect 48504 6103 48556 6112
rect 48504 6069 48513 6103
rect 48513 6069 48547 6103
rect 48547 6069 48556 6103
rect 48504 6060 48556 6069
rect 49792 6103 49844 6112
rect 49792 6069 49801 6103
rect 49801 6069 49835 6103
rect 49835 6069 49844 6103
rect 49792 6060 49844 6069
rect 55864 6060 55916 6112
rect 56692 6196 56744 6248
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 22616 5958 22668 6010
rect 22680 5958 22732 6010
rect 22744 5958 22796 6010
rect 22808 5958 22860 6010
rect 22872 5958 22924 6010
rect 37060 5958 37112 6010
rect 37124 5958 37176 6010
rect 37188 5958 37240 6010
rect 37252 5958 37304 6010
rect 37316 5958 37368 6010
rect 51504 5958 51556 6010
rect 51568 5958 51620 6010
rect 51632 5958 51684 6010
rect 51696 5958 51748 6010
rect 51760 5958 51812 6010
rect 3976 5856 4028 5908
rect 5448 5856 5500 5908
rect 6184 5856 6236 5908
rect 6828 5856 6880 5908
rect 7380 5856 7432 5908
rect 9680 5856 9732 5908
rect 11980 5856 12032 5908
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 7748 5720 7800 5772
rect 8024 5763 8076 5772
rect 8024 5729 8033 5763
rect 8033 5729 8067 5763
rect 8067 5729 8076 5763
rect 8024 5720 8076 5729
rect 8760 5720 8812 5772
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 1768 5652 1820 5704
rect 2688 5652 2740 5704
rect 2780 5652 2832 5704
rect 4436 5652 4488 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 7012 5695 7064 5704
rect 7012 5661 7030 5695
rect 7030 5661 7064 5695
rect 7012 5652 7064 5661
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8024 5584 8076 5636
rect 10232 5720 10284 5772
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 11704 5720 11756 5772
rect 12808 5788 12860 5840
rect 12900 5788 12952 5840
rect 13636 5788 13688 5840
rect 14464 5788 14516 5840
rect 14096 5720 14148 5772
rect 14924 5856 14976 5908
rect 16396 5856 16448 5908
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 19432 5856 19484 5908
rect 20444 5856 20496 5908
rect 20812 5856 20864 5908
rect 22284 5899 22336 5908
rect 22284 5865 22293 5899
rect 22293 5865 22327 5899
rect 22327 5865 22336 5899
rect 22284 5856 22336 5865
rect 22468 5899 22520 5908
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 23020 5856 23072 5908
rect 28540 5856 28592 5908
rect 18696 5788 18748 5840
rect 19892 5788 19944 5840
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 10140 5652 10192 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 12808 5584 12860 5636
rect 13360 5627 13412 5636
rect 13360 5593 13369 5627
rect 13369 5593 13403 5627
rect 13403 5593 13412 5627
rect 13360 5584 13412 5593
rect 13728 5584 13780 5636
rect 14556 5652 14608 5704
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 15936 5720 15988 5772
rect 17960 5720 18012 5772
rect 18328 5763 18380 5772
rect 18328 5729 18337 5763
rect 18337 5729 18371 5763
rect 18371 5729 18380 5763
rect 18328 5720 18380 5729
rect 16304 5652 16356 5704
rect 21180 5720 21232 5772
rect 22928 5720 22980 5772
rect 24584 5788 24636 5840
rect 4344 5516 4396 5568
rect 7564 5516 7616 5568
rect 8668 5516 8720 5568
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 11888 5516 11940 5568
rect 13820 5516 13872 5568
rect 15752 5584 15804 5636
rect 16212 5584 16264 5636
rect 14556 5516 14608 5568
rect 19432 5559 19484 5568
rect 19432 5525 19441 5559
rect 19441 5525 19475 5559
rect 19475 5525 19484 5559
rect 19432 5516 19484 5525
rect 19524 5516 19576 5568
rect 20260 5516 20312 5568
rect 21088 5584 21140 5636
rect 24032 5652 24084 5704
rect 25872 5788 25924 5840
rect 21364 5516 21416 5568
rect 24768 5584 24820 5636
rect 25320 5584 25372 5636
rect 25596 5652 25648 5704
rect 26700 5652 26752 5704
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 26976 5652 27028 5661
rect 27804 5652 27856 5704
rect 30380 5856 30432 5908
rect 33416 5856 33468 5908
rect 38108 5856 38160 5908
rect 38292 5856 38344 5908
rect 38476 5899 38528 5908
rect 38476 5865 38485 5899
rect 38485 5865 38519 5899
rect 38519 5865 38528 5899
rect 38476 5856 38528 5865
rect 38660 5856 38712 5908
rect 41144 5899 41196 5908
rect 41144 5865 41153 5899
rect 41153 5865 41187 5899
rect 41187 5865 41196 5899
rect 41144 5856 41196 5865
rect 41696 5856 41748 5908
rect 43628 5856 43680 5908
rect 32128 5831 32180 5840
rect 32128 5797 32137 5831
rect 32137 5797 32171 5831
rect 32171 5797 32180 5831
rect 32128 5788 32180 5797
rect 30196 5720 30248 5772
rect 33508 5788 33560 5840
rect 33876 5788 33928 5840
rect 35624 5831 35676 5840
rect 35624 5797 35633 5831
rect 35633 5797 35667 5831
rect 35667 5797 35676 5831
rect 35624 5788 35676 5797
rect 38568 5788 38620 5840
rect 41880 5788 41932 5840
rect 42064 5788 42116 5840
rect 47860 5831 47912 5840
rect 47860 5797 47869 5831
rect 47869 5797 47903 5831
rect 47903 5797 47912 5831
rect 47860 5788 47912 5797
rect 33324 5720 33376 5772
rect 22928 5516 22980 5568
rect 25780 5516 25832 5568
rect 27620 5516 27672 5568
rect 28264 5516 28316 5568
rect 28540 5516 28592 5568
rect 29644 5652 29696 5704
rect 30932 5652 30984 5704
rect 31576 5695 31628 5704
rect 31576 5661 31585 5695
rect 31585 5661 31619 5695
rect 31619 5661 31628 5695
rect 31576 5652 31628 5661
rect 31760 5695 31812 5704
rect 31760 5661 31778 5695
rect 31778 5661 31812 5695
rect 31760 5652 31812 5661
rect 32772 5695 32824 5704
rect 32772 5661 32781 5695
rect 32781 5661 32815 5695
rect 32815 5661 32824 5695
rect 38752 5720 38804 5772
rect 32772 5652 32824 5661
rect 33508 5652 33560 5704
rect 36912 5652 36964 5704
rect 37556 5652 37608 5704
rect 40132 5720 40184 5772
rect 40224 5720 40276 5772
rect 45192 5763 45244 5772
rect 45192 5729 45201 5763
rect 45201 5729 45235 5763
rect 45235 5729 45244 5763
rect 45192 5720 45244 5729
rect 47124 5720 47176 5772
rect 47768 5720 47820 5772
rect 51080 5856 51132 5908
rect 53380 5856 53432 5908
rect 55220 5856 55272 5908
rect 56692 5899 56744 5908
rect 56692 5865 56701 5899
rect 56701 5865 56735 5899
rect 56735 5865 56744 5899
rect 56692 5856 56744 5865
rect 56784 5899 56836 5908
rect 56784 5865 56793 5899
rect 56793 5865 56827 5899
rect 56827 5865 56836 5899
rect 56784 5856 56836 5865
rect 58440 5899 58492 5908
rect 58440 5865 58449 5899
rect 58449 5865 58483 5899
rect 58483 5865 58492 5899
rect 58440 5856 58492 5865
rect 50252 5763 50304 5772
rect 50252 5729 50261 5763
rect 50261 5729 50295 5763
rect 50295 5729 50304 5763
rect 50252 5720 50304 5729
rect 29276 5584 29328 5636
rect 36544 5584 36596 5636
rect 40776 5652 40828 5704
rect 37924 5627 37976 5636
rect 37924 5593 37933 5627
rect 37933 5593 37967 5627
rect 37967 5593 37976 5627
rect 37924 5584 37976 5593
rect 39764 5584 39816 5636
rect 43352 5652 43404 5704
rect 47308 5695 47360 5704
rect 47308 5661 47317 5695
rect 47317 5661 47351 5695
rect 47351 5661 47360 5695
rect 47308 5652 47360 5661
rect 48872 5652 48924 5704
rect 49700 5695 49752 5704
rect 49700 5661 49718 5695
rect 49718 5661 49752 5695
rect 49700 5652 49752 5661
rect 50160 5652 50212 5704
rect 50436 5652 50488 5704
rect 52828 5652 52880 5704
rect 57704 5720 57756 5772
rect 56692 5652 56744 5704
rect 44180 5627 44232 5636
rect 44180 5593 44189 5627
rect 44189 5593 44223 5627
rect 44223 5593 44232 5627
rect 44180 5584 44232 5593
rect 46020 5584 46072 5636
rect 52276 5584 52328 5636
rect 52736 5584 52788 5636
rect 54024 5584 54076 5636
rect 55680 5584 55732 5636
rect 56508 5584 56560 5636
rect 58256 5695 58308 5704
rect 58256 5661 58265 5695
rect 58265 5661 58299 5695
rect 58299 5661 58308 5695
rect 58256 5652 58308 5661
rect 29000 5559 29052 5568
rect 29000 5525 29009 5559
rect 29009 5525 29043 5559
rect 29043 5525 29052 5559
rect 29000 5516 29052 5525
rect 29368 5559 29420 5568
rect 29368 5525 29377 5559
rect 29377 5525 29411 5559
rect 29411 5525 29420 5559
rect 29368 5516 29420 5525
rect 32680 5516 32732 5568
rect 32864 5516 32916 5568
rect 33600 5559 33652 5568
rect 33600 5525 33609 5559
rect 33609 5525 33643 5559
rect 33643 5525 33652 5559
rect 33600 5516 33652 5525
rect 37096 5559 37148 5568
rect 37096 5525 37105 5559
rect 37105 5525 37139 5559
rect 37139 5525 37148 5559
rect 37096 5516 37148 5525
rect 38752 5516 38804 5568
rect 41144 5516 41196 5568
rect 41788 5516 41840 5568
rect 42156 5516 42208 5568
rect 42708 5516 42760 5568
rect 44824 5516 44876 5568
rect 47952 5516 48004 5568
rect 49608 5516 49660 5568
rect 51080 5516 51132 5568
rect 57520 5559 57572 5568
rect 57520 5525 57529 5559
rect 57529 5525 57563 5559
rect 57563 5525 57572 5559
rect 57520 5516 57572 5525
rect 15394 5414 15446 5466
rect 15458 5414 15510 5466
rect 15522 5414 15574 5466
rect 15586 5414 15638 5466
rect 15650 5414 15702 5466
rect 29838 5414 29890 5466
rect 29902 5414 29954 5466
rect 29966 5414 30018 5466
rect 30030 5414 30082 5466
rect 30094 5414 30146 5466
rect 44282 5414 44334 5466
rect 44346 5414 44398 5466
rect 44410 5414 44462 5466
rect 44474 5414 44526 5466
rect 44538 5414 44590 5466
rect 58726 5414 58778 5466
rect 58790 5414 58842 5466
rect 58854 5414 58906 5466
rect 58918 5414 58970 5466
rect 58982 5414 59034 5466
rect 2688 5312 2740 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 6368 5312 6420 5364
rect 7380 5312 7432 5364
rect 7748 5312 7800 5364
rect 3516 5244 3568 5296
rect 5172 5244 5224 5296
rect 5632 5244 5684 5296
rect 10140 5312 10192 5364
rect 11060 5312 11112 5364
rect 11152 5312 11204 5364
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 2964 5040 3016 5092
rect 3332 5040 3384 5092
rect 6000 5108 6052 5160
rect 8668 5287 8720 5296
rect 8668 5253 8697 5287
rect 8697 5253 8720 5287
rect 8668 5244 8720 5253
rect 8852 5244 8904 5296
rect 7104 5176 7156 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 13360 5244 13412 5296
rect 14648 5312 14700 5364
rect 16120 5355 16172 5364
rect 16120 5321 16129 5355
rect 16129 5321 16163 5355
rect 16163 5321 16172 5355
rect 16120 5312 16172 5321
rect 19892 5312 19944 5364
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 17960 5176 18012 5228
rect 11060 5108 11112 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 11704 5151 11756 5160
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 4620 4972 4672 5024
rect 4988 4972 5040 5024
rect 5172 4972 5224 5024
rect 7380 4972 7432 5024
rect 7840 4972 7892 5024
rect 12072 5040 12124 5092
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 12164 4972 12216 5024
rect 12348 4972 12400 5024
rect 17224 5151 17276 5160
rect 17224 5117 17233 5151
rect 17233 5117 17267 5151
rect 17267 5117 17276 5151
rect 17224 5108 17276 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19248 5151 19300 5160
rect 19248 5117 19257 5151
rect 19257 5117 19291 5151
rect 19291 5117 19300 5151
rect 19248 5108 19300 5117
rect 19800 5176 19852 5228
rect 21364 5312 21416 5364
rect 22192 5244 22244 5296
rect 23940 5244 23992 5296
rect 18972 5040 19024 5092
rect 19432 5040 19484 5092
rect 20720 5108 20772 5160
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 21548 5040 21600 5092
rect 24860 5176 24912 5228
rect 25596 5219 25648 5228
rect 25596 5185 25630 5219
rect 25630 5185 25648 5219
rect 25596 5176 25648 5185
rect 24676 5108 24728 5160
rect 26976 5312 27028 5364
rect 27988 5355 28040 5364
rect 27988 5321 27997 5355
rect 27997 5321 28031 5355
rect 28031 5321 28040 5355
rect 27988 5312 28040 5321
rect 29276 5312 29328 5364
rect 29644 5312 29696 5364
rect 30288 5312 30340 5364
rect 31116 5312 31168 5364
rect 31300 5355 31352 5364
rect 31300 5321 31309 5355
rect 31309 5321 31343 5355
rect 31343 5321 31352 5355
rect 31300 5312 31352 5321
rect 32128 5312 32180 5364
rect 27344 5244 27396 5296
rect 27620 5108 27672 5160
rect 15936 4972 15988 5024
rect 16120 4972 16172 5024
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 18512 4972 18564 5024
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 21916 5015 21968 5024
rect 21916 4981 21925 5015
rect 21925 4981 21959 5015
rect 21959 4981 21968 5015
rect 21916 4972 21968 4981
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 25228 5015 25280 5024
rect 25228 4981 25237 5015
rect 25237 4981 25271 5015
rect 25271 4981 25280 5015
rect 25228 4972 25280 4981
rect 25320 4972 25372 5024
rect 27712 4972 27764 5024
rect 27804 4972 27856 5024
rect 28724 4972 28776 5024
rect 28816 4972 28868 5024
rect 32588 5244 32640 5296
rect 34888 5287 34940 5296
rect 34888 5253 34897 5287
rect 34897 5253 34931 5287
rect 34931 5253 34940 5287
rect 34888 5244 34940 5253
rect 35992 5312 36044 5364
rect 36084 5355 36136 5364
rect 36084 5321 36093 5355
rect 36093 5321 36127 5355
rect 36127 5321 36136 5355
rect 36084 5312 36136 5321
rect 37096 5312 37148 5364
rect 37648 5355 37700 5364
rect 37648 5321 37657 5355
rect 37657 5321 37691 5355
rect 37691 5321 37700 5355
rect 37648 5312 37700 5321
rect 40500 5312 40552 5364
rect 41788 5312 41840 5364
rect 44180 5312 44232 5364
rect 45192 5312 45244 5364
rect 45652 5355 45704 5364
rect 45652 5321 45661 5355
rect 45661 5321 45695 5355
rect 45695 5321 45704 5355
rect 45652 5312 45704 5321
rect 46572 5312 46624 5364
rect 36452 5244 36504 5296
rect 36728 5287 36780 5296
rect 36728 5253 36737 5287
rect 36737 5253 36771 5287
rect 36771 5253 36780 5287
rect 36728 5244 36780 5253
rect 29368 5176 29420 5228
rect 31300 5176 31352 5228
rect 32128 5176 32180 5228
rect 32864 5176 32916 5228
rect 33232 5219 33284 5228
rect 33232 5185 33241 5219
rect 33241 5185 33275 5219
rect 33275 5185 33284 5219
rect 33232 5176 33284 5185
rect 33600 5176 33652 5228
rect 33876 5176 33928 5228
rect 35808 5176 35860 5228
rect 36176 5176 36228 5228
rect 30196 5151 30248 5160
rect 30196 5117 30205 5151
rect 30205 5117 30239 5151
rect 30239 5117 30248 5151
rect 30196 5108 30248 5117
rect 31392 5108 31444 5160
rect 32312 5108 32364 5160
rect 32404 5108 32456 5160
rect 34428 5108 34480 5160
rect 38660 5176 38712 5228
rect 42800 5287 42852 5296
rect 42800 5253 42809 5287
rect 42809 5253 42843 5287
rect 42843 5253 42852 5287
rect 42800 5244 42852 5253
rect 41236 5176 41288 5228
rect 42616 5176 42668 5228
rect 37740 5151 37792 5160
rect 37740 5117 37749 5151
rect 37749 5117 37783 5151
rect 37783 5117 37792 5151
rect 37740 5108 37792 5117
rect 33508 5040 33560 5092
rect 33600 5040 33652 5092
rect 33784 5040 33836 5092
rect 38752 5108 38804 5160
rect 34612 4972 34664 5024
rect 35808 4972 35860 5024
rect 36912 4972 36964 5024
rect 37556 4972 37608 5024
rect 38016 4972 38068 5024
rect 40868 5040 40920 5092
rect 41052 5151 41104 5160
rect 41052 5117 41061 5151
rect 41061 5117 41095 5151
rect 41095 5117 41104 5151
rect 41052 5108 41104 5117
rect 42708 5151 42760 5160
rect 42708 5117 42717 5151
rect 42717 5117 42751 5151
rect 42751 5117 42760 5151
rect 42708 5108 42760 5117
rect 45008 5040 45060 5092
rect 47492 5244 47544 5296
rect 47768 5176 47820 5228
rect 40500 4972 40552 5024
rect 41328 4972 41380 5024
rect 42156 4972 42208 5024
rect 43536 4972 43588 5024
rect 45376 4972 45428 5024
rect 46204 5151 46256 5160
rect 46204 5117 46213 5151
rect 46213 5117 46247 5151
rect 46247 5117 46256 5151
rect 46204 5108 46256 5117
rect 47676 5108 47728 5160
rect 50436 5244 50488 5296
rect 51080 5355 51132 5364
rect 51080 5321 51089 5355
rect 51089 5321 51123 5355
rect 51123 5321 51132 5355
rect 51080 5312 51132 5321
rect 52552 5312 52604 5364
rect 54024 5355 54076 5364
rect 54024 5321 54033 5355
rect 54033 5321 54067 5355
rect 54067 5321 54076 5355
rect 54024 5312 54076 5321
rect 54944 5355 54996 5364
rect 54944 5321 54953 5355
rect 54953 5321 54987 5355
rect 54987 5321 54996 5355
rect 54944 5312 54996 5321
rect 55680 5355 55732 5364
rect 55680 5321 55689 5355
rect 55689 5321 55723 5355
rect 55723 5321 55732 5355
rect 55680 5312 55732 5321
rect 57520 5312 57572 5364
rect 57612 5355 57664 5364
rect 57612 5321 57621 5355
rect 57621 5321 57655 5355
rect 57655 5321 57664 5355
rect 57612 5312 57664 5321
rect 52644 5244 52696 5296
rect 53104 5244 53156 5296
rect 50160 5176 50212 5228
rect 50896 5219 50948 5228
rect 50896 5185 50905 5219
rect 50905 5185 50939 5219
rect 50939 5185 50948 5219
rect 50896 5176 50948 5185
rect 53380 5219 53432 5228
rect 53380 5185 53389 5219
rect 53389 5185 53423 5219
rect 53423 5185 53432 5219
rect 53380 5176 53432 5185
rect 57336 5244 57388 5296
rect 50344 5108 50396 5160
rect 53012 5108 53064 5160
rect 46204 4972 46256 5024
rect 46480 5015 46532 5024
rect 46480 4981 46489 5015
rect 46489 4981 46523 5015
rect 46523 4981 46532 5015
rect 46480 4972 46532 4981
rect 48872 5015 48924 5024
rect 48872 4981 48881 5015
rect 48881 4981 48915 5015
rect 48915 4981 48924 5015
rect 55220 5040 55272 5092
rect 55956 5176 56008 5228
rect 56968 5219 57020 5228
rect 56968 5185 56977 5219
rect 56977 5185 57011 5219
rect 57011 5185 57020 5219
rect 56968 5176 57020 5185
rect 57152 5176 57204 5228
rect 56140 5108 56192 5160
rect 56600 5108 56652 5160
rect 48872 4972 48924 4981
rect 51172 4972 51224 5024
rect 52552 4972 52604 5024
rect 53748 5015 53800 5024
rect 53748 4981 53757 5015
rect 53757 4981 53791 5015
rect 53791 4981 53800 5015
rect 53748 4972 53800 4981
rect 53840 4972 53892 5024
rect 55404 5015 55456 5024
rect 55404 4981 55413 5015
rect 55413 4981 55447 5015
rect 55447 4981 55456 5015
rect 55404 4972 55456 4981
rect 57796 4972 57848 5024
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 22616 4870 22668 4922
rect 22680 4870 22732 4922
rect 22744 4870 22796 4922
rect 22808 4870 22860 4922
rect 22872 4870 22924 4922
rect 37060 4870 37112 4922
rect 37124 4870 37176 4922
rect 37188 4870 37240 4922
rect 37252 4870 37304 4922
rect 37316 4870 37368 4922
rect 51504 4870 51556 4922
rect 51568 4870 51620 4922
rect 51632 4870 51684 4922
rect 51696 4870 51748 4922
rect 51760 4870 51812 4922
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 2596 4768 2648 4820
rect 4620 4768 4672 4820
rect 6092 4768 6144 4820
rect 6184 4768 6236 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 8944 4768 8996 4820
rect 9404 4768 9456 4820
rect 9772 4768 9824 4820
rect 4988 4700 5040 4752
rect 3240 4632 3292 4684
rect 8300 4700 8352 4752
rect 9680 4700 9732 4752
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 8760 4632 8812 4684
rect 9036 4632 9088 4684
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 3148 4564 3200 4616
rect 4620 4564 4672 4616
rect 5908 4564 5960 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7104 4564 7156 4616
rect 5172 4496 5224 4548
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 10508 4564 10560 4616
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 15200 4700 15252 4752
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 20076 4768 20128 4820
rect 20444 4768 20496 4820
rect 24124 4768 24176 4820
rect 24216 4768 24268 4820
rect 24308 4768 24360 4820
rect 15844 4632 15896 4684
rect 7748 4496 7800 4548
rect 11152 4496 11204 4548
rect 11428 4496 11480 4548
rect 13084 4496 13136 4548
rect 13912 4564 13964 4616
rect 16212 4564 16264 4616
rect 7932 4428 7984 4480
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 9128 4428 9180 4480
rect 11060 4428 11112 4480
rect 11520 4428 11572 4480
rect 11704 4428 11756 4480
rect 12992 4428 13044 4480
rect 15292 4496 15344 4548
rect 15752 4496 15804 4548
rect 16672 4496 16724 4548
rect 21364 4632 21416 4684
rect 24032 4675 24084 4684
rect 24032 4641 24041 4675
rect 24041 4641 24075 4675
rect 24075 4641 24084 4675
rect 24032 4632 24084 4641
rect 18512 4564 18564 4616
rect 18052 4496 18104 4548
rect 19248 4496 19300 4548
rect 20812 4607 20864 4616
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 21916 4564 21968 4616
rect 25688 4700 25740 4752
rect 26516 4768 26568 4820
rect 27620 4811 27672 4820
rect 27620 4777 27629 4811
rect 27629 4777 27663 4811
rect 27663 4777 27672 4811
rect 27620 4768 27672 4777
rect 27712 4768 27764 4820
rect 28816 4700 28868 4752
rect 24676 4632 24728 4684
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 26976 4632 27028 4684
rect 24308 4564 24360 4616
rect 25044 4607 25096 4616
rect 25044 4573 25053 4607
rect 25053 4573 25087 4607
rect 25087 4573 25096 4607
rect 25044 4564 25096 4573
rect 26056 4607 26108 4616
rect 26056 4573 26065 4607
rect 26065 4573 26099 4607
rect 26099 4573 26108 4607
rect 26056 4564 26108 4573
rect 26608 4607 26660 4616
rect 26608 4573 26617 4607
rect 26617 4573 26651 4607
rect 26651 4573 26660 4607
rect 26608 4564 26660 4573
rect 28264 4607 28316 4616
rect 19616 4539 19668 4548
rect 19616 4505 19625 4539
rect 19625 4505 19659 4539
rect 19659 4505 19668 4539
rect 19616 4496 19668 4505
rect 20260 4496 20312 4548
rect 26332 4496 26384 4548
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 28356 4607 28408 4616
rect 28356 4573 28365 4607
rect 28365 4573 28399 4607
rect 28399 4573 28408 4607
rect 28356 4564 28408 4573
rect 28080 4496 28132 4548
rect 30748 4700 30800 4752
rect 31484 4700 31536 4752
rect 32588 4700 32640 4752
rect 36176 4700 36228 4752
rect 36452 4743 36504 4752
rect 36452 4709 36461 4743
rect 36461 4709 36495 4743
rect 36495 4709 36504 4743
rect 36452 4700 36504 4709
rect 37740 4768 37792 4820
rect 37924 4768 37976 4820
rect 38016 4811 38068 4820
rect 38016 4777 38025 4811
rect 38025 4777 38059 4811
rect 38059 4777 38068 4811
rect 38016 4768 38068 4777
rect 38844 4811 38896 4820
rect 38844 4777 38853 4811
rect 38853 4777 38887 4811
rect 38887 4777 38896 4811
rect 38844 4768 38896 4777
rect 39672 4768 39724 4820
rect 41880 4768 41932 4820
rect 42708 4768 42760 4820
rect 46020 4811 46072 4820
rect 46020 4777 46029 4811
rect 46029 4777 46063 4811
rect 46063 4777 46072 4811
rect 46020 4768 46072 4777
rect 46480 4768 46532 4820
rect 48504 4768 48556 4820
rect 50160 4768 50212 4820
rect 51356 4768 51408 4820
rect 52552 4768 52604 4820
rect 57152 4768 57204 4820
rect 57704 4768 57756 4820
rect 31300 4632 31352 4684
rect 29184 4496 29236 4548
rect 30196 4496 30248 4548
rect 14096 4428 14148 4480
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 14556 4428 14608 4480
rect 16120 4428 16172 4480
rect 18880 4428 18932 4480
rect 19432 4428 19484 4480
rect 21088 4428 21140 4480
rect 23480 4471 23532 4480
rect 23480 4437 23489 4471
rect 23489 4437 23523 4471
rect 23523 4437 23532 4471
rect 23480 4428 23532 4437
rect 23940 4471 23992 4480
rect 23940 4437 23949 4471
rect 23949 4437 23983 4471
rect 23983 4437 23992 4471
rect 23940 4428 23992 4437
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 26884 4471 26936 4480
rect 26884 4437 26893 4471
rect 26893 4437 26927 4471
rect 26927 4437 26936 4471
rect 26884 4428 26936 4437
rect 28632 4471 28684 4480
rect 28632 4437 28641 4471
rect 28641 4437 28675 4471
rect 28675 4437 28684 4471
rect 28632 4428 28684 4437
rect 28724 4428 28776 4480
rect 32036 4496 32088 4548
rect 33784 4632 33836 4684
rect 32864 4564 32916 4616
rect 33508 4564 33560 4616
rect 33876 4607 33928 4616
rect 33876 4573 33885 4607
rect 33885 4573 33919 4607
rect 33919 4573 33928 4607
rect 33876 4564 33928 4573
rect 35624 4632 35676 4684
rect 36544 4632 36596 4684
rect 37004 4675 37056 4684
rect 37004 4641 37013 4675
rect 37013 4641 37047 4675
rect 37047 4641 37056 4675
rect 37004 4632 37056 4641
rect 32772 4496 32824 4548
rect 34152 4539 34204 4548
rect 34152 4505 34161 4539
rect 34161 4505 34195 4539
rect 34195 4505 34204 4539
rect 34152 4496 34204 4505
rect 31944 4428 31996 4480
rect 32588 4471 32640 4480
rect 32588 4437 32597 4471
rect 32597 4437 32631 4471
rect 32631 4437 32640 4471
rect 32588 4428 32640 4437
rect 35164 4539 35216 4548
rect 35164 4505 35173 4539
rect 35173 4505 35207 4539
rect 35207 4505 35216 4539
rect 35164 4496 35216 4505
rect 35716 4564 35768 4616
rect 36176 4564 36228 4616
rect 36820 4607 36872 4616
rect 40224 4632 40276 4684
rect 41052 4700 41104 4752
rect 41236 4743 41288 4752
rect 41236 4709 41245 4743
rect 41245 4709 41279 4743
rect 41279 4709 41288 4743
rect 41236 4700 41288 4709
rect 41328 4632 41380 4684
rect 41972 4632 42024 4684
rect 44180 4632 44232 4684
rect 44824 4632 44876 4684
rect 48688 4700 48740 4752
rect 49424 4700 49476 4752
rect 36820 4573 36854 4607
rect 36854 4573 36872 4607
rect 36820 4564 36872 4573
rect 35900 4496 35952 4548
rect 40408 4607 40460 4616
rect 40408 4573 40417 4607
rect 40417 4573 40451 4607
rect 40451 4573 40460 4607
rect 40408 4564 40460 4573
rect 40592 4496 40644 4548
rect 38292 4471 38344 4480
rect 38292 4437 38301 4471
rect 38301 4437 38335 4471
rect 38335 4437 38344 4471
rect 38292 4428 38344 4437
rect 39856 4471 39908 4480
rect 39856 4437 39865 4471
rect 39865 4437 39899 4471
rect 39899 4437 39908 4471
rect 39856 4428 39908 4437
rect 41788 4607 41840 4616
rect 41788 4573 41797 4607
rect 41797 4573 41831 4607
rect 41831 4573 41840 4607
rect 41788 4564 41840 4573
rect 42616 4564 42668 4616
rect 44088 4564 44140 4616
rect 44640 4607 44692 4616
rect 44640 4573 44649 4607
rect 44649 4573 44683 4607
rect 44683 4573 44692 4607
rect 44640 4564 44692 4573
rect 44916 4564 44968 4616
rect 45928 4607 45980 4616
rect 45928 4573 45937 4607
rect 45937 4573 45971 4607
rect 45971 4573 45980 4607
rect 45928 4564 45980 4573
rect 50804 4700 50856 4752
rect 55956 4700 56008 4752
rect 56508 4743 56560 4752
rect 56508 4709 56517 4743
rect 56517 4709 56551 4743
rect 56551 4709 56560 4743
rect 56508 4700 56560 4709
rect 47308 4607 47360 4616
rect 47308 4573 47317 4607
rect 47317 4573 47351 4607
rect 47351 4573 47360 4607
rect 47308 4564 47360 4573
rect 47492 4607 47544 4616
rect 47492 4573 47501 4607
rect 47501 4573 47535 4607
rect 47535 4573 47544 4607
rect 47492 4564 47544 4573
rect 51172 4632 51224 4684
rect 52460 4632 52512 4684
rect 54024 4632 54076 4684
rect 49700 4564 49752 4616
rect 51448 4607 51500 4616
rect 51448 4573 51457 4607
rect 51457 4573 51491 4607
rect 51491 4573 51500 4607
rect 51448 4564 51500 4573
rect 52000 4564 52052 4616
rect 52092 4607 52144 4616
rect 52092 4573 52101 4607
rect 52101 4573 52135 4607
rect 52135 4573 52144 4607
rect 52092 4564 52144 4573
rect 53104 4607 53156 4616
rect 53104 4573 53113 4607
rect 53113 4573 53147 4607
rect 53147 4573 53156 4607
rect 53104 4564 53156 4573
rect 54116 4607 54168 4616
rect 54116 4573 54125 4607
rect 54125 4573 54159 4607
rect 54159 4573 54168 4607
rect 54116 4564 54168 4573
rect 51356 4496 51408 4548
rect 55496 4607 55548 4616
rect 55496 4573 55505 4607
rect 55505 4573 55539 4607
rect 55539 4573 55548 4607
rect 55496 4564 55548 4573
rect 55680 4607 55732 4616
rect 55680 4573 55689 4607
rect 55689 4573 55723 4607
rect 55723 4573 55732 4607
rect 55680 4564 55732 4573
rect 55772 4607 55824 4616
rect 55772 4573 55781 4607
rect 55781 4573 55815 4607
rect 55815 4573 55824 4607
rect 55772 4564 55824 4573
rect 57796 4564 57848 4616
rect 58164 4607 58216 4616
rect 58164 4573 58173 4607
rect 58173 4573 58207 4607
rect 58207 4573 58216 4607
rect 58164 4564 58216 4573
rect 43812 4428 43864 4480
rect 45008 4471 45060 4480
rect 45008 4437 45017 4471
rect 45017 4437 45051 4471
rect 45051 4437 45060 4471
rect 45008 4428 45060 4437
rect 45284 4471 45336 4480
rect 45284 4437 45293 4471
rect 45293 4437 45327 4471
rect 45327 4437 45336 4471
rect 45284 4428 45336 4437
rect 46756 4471 46808 4480
rect 46756 4437 46765 4471
rect 46765 4437 46799 4471
rect 46799 4437 46808 4471
rect 46756 4428 46808 4437
rect 49608 4428 49660 4480
rect 50528 4428 50580 4480
rect 50804 4471 50856 4480
rect 50804 4437 50813 4471
rect 50813 4437 50847 4471
rect 50847 4437 50856 4471
rect 50804 4428 50856 4437
rect 50896 4471 50948 4480
rect 50896 4437 50905 4471
rect 50905 4437 50939 4471
rect 50939 4437 50948 4471
rect 50896 4428 50948 4437
rect 52736 4471 52788 4480
rect 52736 4437 52745 4471
rect 52745 4437 52779 4471
rect 52779 4437 52788 4471
rect 52736 4428 52788 4437
rect 53196 4471 53248 4480
rect 53196 4437 53205 4471
rect 53205 4437 53239 4471
rect 53239 4437 53248 4471
rect 53196 4428 53248 4437
rect 53564 4471 53616 4480
rect 53564 4437 53573 4471
rect 53573 4437 53607 4471
rect 53607 4437 53616 4471
rect 53564 4428 53616 4437
rect 56600 4496 56652 4548
rect 57428 4496 57480 4548
rect 56048 4428 56100 4480
rect 56416 4471 56468 4480
rect 56416 4437 56425 4471
rect 56425 4437 56459 4471
rect 56459 4437 56468 4471
rect 56416 4428 56468 4437
rect 57060 4428 57112 4480
rect 15394 4326 15446 4378
rect 15458 4326 15510 4378
rect 15522 4326 15574 4378
rect 15586 4326 15638 4378
rect 15650 4326 15702 4378
rect 29838 4326 29890 4378
rect 29902 4326 29954 4378
rect 29966 4326 30018 4378
rect 30030 4326 30082 4378
rect 30094 4326 30146 4378
rect 44282 4326 44334 4378
rect 44346 4326 44398 4378
rect 44410 4326 44462 4378
rect 44474 4326 44526 4378
rect 44538 4326 44590 4378
rect 58726 4326 58778 4378
rect 58790 4326 58842 4378
rect 58854 4326 58906 4378
rect 58918 4326 58970 4378
rect 58982 4326 59034 4378
rect 2872 4224 2924 4276
rect 3608 4224 3660 4276
rect 4620 4224 4672 4276
rect 5080 4224 5132 4276
rect 2228 4156 2280 4208
rect 3516 4156 3568 4208
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 5632 4156 5684 4208
rect 4252 4088 4304 4140
rect 7104 4156 7156 4208
rect 2964 4020 3016 4072
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 4160 4020 4212 4072
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 6828 4088 6880 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7012 4088 7064 4140
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 7932 4267 7984 4276
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 9404 4224 9456 4276
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 11428 4224 11480 4276
rect 11704 4224 11756 4276
rect 14372 4224 14424 4276
rect 15844 4224 15896 4276
rect 16396 4267 16448 4276
rect 16396 4233 16405 4267
rect 16405 4233 16439 4267
rect 16439 4233 16448 4267
rect 16396 4224 16448 4233
rect 17224 4224 17276 4276
rect 7656 4156 7708 4208
rect 9036 4156 9088 4208
rect 10600 4199 10652 4208
rect 10600 4165 10609 4199
rect 10609 4165 10643 4199
rect 10643 4165 10652 4199
rect 10600 4156 10652 4165
rect 14004 4156 14056 4208
rect 15292 4156 15344 4208
rect 17500 4224 17552 4276
rect 19616 4224 19668 4276
rect 20904 4224 20956 4276
rect 24308 4224 24360 4276
rect 24400 4224 24452 4276
rect 27620 4224 27672 4276
rect 20536 4199 20588 4208
rect 20536 4165 20545 4199
rect 20545 4165 20579 4199
rect 20579 4165 20588 4199
rect 20536 4156 20588 4165
rect 7564 4088 7616 4140
rect 7748 4088 7800 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8576 4088 8628 4140
rect 9312 4088 9364 4140
rect 9864 4088 9916 4140
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 5816 4063 5868 4072
rect 4988 4020 5040 4029
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 5816 4020 5868 4029
rect 6184 4020 6236 4072
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 7196 4020 7248 4072
rect 12348 4088 12400 4140
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 12808 4020 12860 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 5080 3952 5132 4004
rect 5632 3952 5684 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 6368 3884 6420 3936
rect 7564 3884 7616 3936
rect 10600 3952 10652 4004
rect 9128 3884 9180 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11520 3884 11572 3936
rect 13636 4020 13688 4072
rect 13636 3884 13688 3936
rect 15384 4020 15436 4072
rect 15936 4020 15988 4072
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 20812 4088 20864 4140
rect 21640 4131 21692 4140
rect 21640 4097 21649 4131
rect 21649 4097 21683 4131
rect 21683 4097 21692 4131
rect 21640 4088 21692 4097
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 19064 4020 19116 4072
rect 19432 4020 19484 4072
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 22284 4088 22336 4097
rect 23940 4156 23992 4208
rect 13912 3952 13964 4004
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 15016 3884 15068 3936
rect 16856 3952 16908 4004
rect 17868 3952 17920 4004
rect 19892 3952 19944 4004
rect 20352 3952 20404 4004
rect 20536 3952 20588 4004
rect 21824 3952 21876 4004
rect 24492 4020 24544 4072
rect 27344 4199 27396 4208
rect 27344 4165 27353 4199
rect 27353 4165 27387 4199
rect 27387 4165 27396 4199
rect 27344 4156 27396 4165
rect 32588 4224 32640 4276
rect 32680 4224 32732 4276
rect 37464 4224 37516 4276
rect 38292 4224 38344 4276
rect 40408 4224 40460 4276
rect 40500 4267 40552 4276
rect 40500 4233 40509 4267
rect 40509 4233 40543 4267
rect 40543 4233 40552 4267
rect 40500 4224 40552 4233
rect 44180 4224 44232 4276
rect 44272 4224 44324 4276
rect 44824 4224 44876 4276
rect 45928 4224 45980 4276
rect 46756 4224 46808 4276
rect 47952 4267 48004 4276
rect 47952 4233 47961 4267
rect 47961 4233 47995 4267
rect 47995 4233 48004 4267
rect 47952 4224 48004 4233
rect 49700 4224 49752 4276
rect 49884 4224 49936 4276
rect 50804 4267 50856 4276
rect 50804 4233 50813 4267
rect 50813 4233 50847 4267
rect 50847 4233 50856 4267
rect 50804 4224 50856 4233
rect 50896 4224 50948 4276
rect 51448 4224 51500 4276
rect 27252 4131 27304 4140
rect 27252 4097 27261 4131
rect 27261 4097 27295 4131
rect 27295 4097 27304 4131
rect 27252 4088 27304 4097
rect 27528 4088 27580 4140
rect 28724 4088 28776 4140
rect 28816 4088 28868 4140
rect 29460 4131 29512 4140
rect 29460 4097 29469 4131
rect 29469 4097 29503 4131
rect 29503 4097 29512 4131
rect 29460 4088 29512 4097
rect 29644 4088 29696 4140
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 21456 3927 21508 3936
rect 21456 3893 21465 3927
rect 21465 3893 21499 3927
rect 21499 3893 21508 3927
rect 21456 3884 21508 3893
rect 24308 3927 24360 3936
rect 24308 3893 24317 3927
rect 24317 3893 24351 3927
rect 24351 3893 24360 3927
rect 24308 3884 24360 3893
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 25780 4063 25832 4072
rect 25780 4029 25789 4063
rect 25789 4029 25823 4063
rect 25823 4029 25832 4063
rect 25780 4020 25832 4029
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 26056 3952 26108 4004
rect 29736 4020 29788 4072
rect 30380 4020 30432 4072
rect 30840 4020 30892 4072
rect 26700 3884 26752 3936
rect 27068 3927 27120 3936
rect 27068 3893 27077 3927
rect 27077 3893 27111 3927
rect 27111 3893 27120 3927
rect 27068 3884 27120 3893
rect 27344 3927 27396 3936
rect 27344 3893 27353 3927
rect 27353 3893 27387 3927
rect 27387 3893 27396 3927
rect 27344 3884 27396 3893
rect 27804 3927 27856 3936
rect 27804 3893 27813 3927
rect 27813 3893 27847 3927
rect 27847 3893 27856 3927
rect 27804 3884 27856 3893
rect 30932 3884 30984 3936
rect 31300 4063 31352 4072
rect 31300 4029 31309 4063
rect 31309 4029 31343 4063
rect 31343 4029 31352 4063
rect 31300 4020 31352 4029
rect 31760 4063 31812 4072
rect 31760 4029 31769 4063
rect 31769 4029 31803 4063
rect 31803 4029 31812 4063
rect 31760 4020 31812 4029
rect 31944 4063 31996 4072
rect 31944 4029 31953 4063
rect 31953 4029 31987 4063
rect 31987 4029 31996 4063
rect 31944 4020 31996 4029
rect 32496 4131 32548 4140
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 32864 4088 32916 4140
rect 33232 4131 33284 4140
rect 33232 4097 33241 4131
rect 33241 4097 33275 4131
rect 33275 4097 33284 4131
rect 33232 4088 33284 4097
rect 33784 4131 33836 4140
rect 33784 4097 33793 4131
rect 33793 4097 33827 4131
rect 33827 4097 33836 4131
rect 33784 4088 33836 4097
rect 33968 4131 34020 4140
rect 33968 4097 33977 4131
rect 33977 4097 34011 4131
rect 34011 4097 34020 4131
rect 33968 4088 34020 4097
rect 35992 4088 36044 4140
rect 36268 4088 36320 4140
rect 33600 4020 33652 4072
rect 33876 4020 33928 4072
rect 34704 4020 34756 4072
rect 35348 4020 35400 4072
rect 36084 4020 36136 4072
rect 36820 4020 36872 4072
rect 37096 4131 37148 4140
rect 37096 4097 37105 4131
rect 37105 4097 37139 4131
rect 37139 4097 37148 4131
rect 37096 4088 37148 4097
rect 37832 4063 37884 4072
rect 37832 4029 37841 4063
rect 37841 4029 37875 4063
rect 37875 4029 37884 4063
rect 37832 4020 37884 4029
rect 35624 3952 35676 4004
rect 34060 3884 34112 3936
rect 34520 3927 34572 3936
rect 34520 3893 34529 3927
rect 34529 3893 34563 3927
rect 34563 3893 34572 3927
rect 34520 3884 34572 3893
rect 36636 3884 36688 3936
rect 37464 3884 37516 3936
rect 39856 4156 39908 4208
rect 40132 4156 40184 4208
rect 41236 4199 41288 4208
rect 38660 4088 38712 4140
rect 41236 4165 41245 4199
rect 41245 4165 41279 4199
rect 41279 4165 41288 4199
rect 41236 4156 41288 4165
rect 42984 4156 43036 4208
rect 45284 4156 45336 4208
rect 39580 4020 39632 4072
rect 40224 3952 40276 4004
rect 41052 4063 41104 4072
rect 41052 4029 41061 4063
rect 41061 4029 41095 4063
rect 41095 4029 41104 4063
rect 41052 4020 41104 4029
rect 41604 4088 41656 4140
rect 42156 4020 42208 4072
rect 42616 4063 42668 4072
rect 42616 4029 42625 4063
rect 42625 4029 42659 4063
rect 42659 4029 42668 4063
rect 42616 4020 42668 4029
rect 43812 4131 43864 4140
rect 43812 4097 43821 4131
rect 43821 4097 43855 4131
rect 43855 4097 43864 4131
rect 43812 4088 43864 4097
rect 44272 4131 44324 4140
rect 44272 4097 44281 4131
rect 44281 4097 44315 4131
rect 44315 4097 44324 4131
rect 44272 4088 44324 4097
rect 44640 4131 44692 4140
rect 44640 4097 44649 4131
rect 44649 4097 44683 4131
rect 44683 4097 44692 4131
rect 44640 4088 44692 4097
rect 45192 4088 45244 4140
rect 46204 4088 46256 4140
rect 45744 4020 45796 4072
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 47216 4131 47268 4140
rect 47216 4097 47225 4131
rect 47225 4097 47259 4131
rect 47259 4097 47268 4131
rect 47216 4088 47268 4097
rect 49792 4156 49844 4208
rect 53932 4156 53984 4208
rect 48412 4088 48464 4140
rect 48596 4131 48648 4140
rect 48596 4097 48605 4131
rect 48605 4097 48639 4131
rect 48639 4097 48648 4131
rect 48596 4088 48648 4097
rect 40316 3884 40368 3936
rect 41236 3884 41288 3936
rect 44456 3952 44508 4004
rect 45836 3952 45888 4004
rect 47308 3952 47360 4004
rect 47584 4020 47636 4072
rect 47860 4063 47912 4072
rect 47860 4029 47869 4063
rect 47869 4029 47903 4063
rect 47903 4029 47912 4063
rect 47860 4020 47912 4029
rect 49608 4088 49660 4140
rect 50344 4088 50396 4140
rect 50528 4088 50580 4140
rect 51264 4088 51316 4140
rect 52736 4088 52788 4140
rect 55312 4224 55364 4276
rect 55496 4224 55548 4276
rect 56416 4224 56468 4276
rect 55864 4156 55916 4208
rect 54760 4131 54812 4140
rect 54760 4097 54769 4131
rect 54769 4097 54803 4131
rect 54803 4097 54812 4131
rect 54760 4088 54812 4097
rect 55956 4131 56008 4140
rect 55956 4097 55965 4131
rect 55965 4097 55999 4131
rect 55999 4097 56008 4131
rect 55956 4088 56008 4097
rect 56968 4156 57020 4208
rect 51080 4020 51132 4072
rect 52644 4020 52696 4072
rect 52920 4063 52972 4072
rect 52920 4029 52929 4063
rect 52929 4029 52963 4063
rect 52963 4029 52972 4063
rect 52920 4020 52972 4029
rect 53104 4020 53156 4072
rect 41604 3927 41656 3936
rect 41604 3893 41613 3927
rect 41613 3893 41647 3927
rect 41647 3893 41656 3927
rect 41604 3884 41656 3893
rect 42248 3927 42300 3936
rect 42248 3893 42257 3927
rect 42257 3893 42291 3927
rect 42291 3893 42300 3927
rect 42248 3884 42300 3893
rect 45284 3884 45336 3936
rect 48320 3927 48372 3936
rect 48320 3893 48329 3927
rect 48329 3893 48363 3927
rect 48363 3893 48372 3927
rect 48320 3884 48372 3893
rect 48688 3927 48740 3936
rect 48688 3893 48697 3927
rect 48697 3893 48731 3927
rect 48731 3893 48740 3927
rect 48688 3884 48740 3893
rect 52552 3952 52604 4004
rect 54024 4020 54076 4072
rect 54116 4020 54168 4072
rect 54852 4020 54904 4072
rect 55036 4063 55088 4072
rect 55036 4029 55045 4063
rect 55045 4029 55079 4063
rect 55079 4029 55088 4063
rect 55036 4020 55088 4029
rect 55588 4020 55640 4072
rect 55772 4063 55824 4072
rect 55772 4029 55781 4063
rect 55781 4029 55815 4063
rect 55815 4029 55824 4063
rect 55772 4020 55824 4029
rect 55956 3952 56008 4004
rect 49700 3884 49752 3936
rect 51908 3927 51960 3936
rect 51908 3893 51917 3927
rect 51917 3893 51951 3927
rect 51951 3893 51960 3927
rect 51908 3884 51960 3893
rect 54024 3927 54076 3936
rect 54024 3893 54033 3927
rect 54033 3893 54067 3927
rect 54067 3893 54076 3927
rect 54024 3884 54076 3893
rect 56692 4063 56744 4072
rect 56692 4029 56701 4063
rect 56701 4029 56735 4063
rect 56735 4029 56744 4063
rect 56692 4020 56744 4029
rect 57244 4020 57296 4072
rect 57520 3884 57572 3936
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 22616 3782 22668 3834
rect 22680 3782 22732 3834
rect 22744 3782 22796 3834
rect 22808 3782 22860 3834
rect 22872 3782 22924 3834
rect 37060 3782 37112 3834
rect 37124 3782 37176 3834
rect 37188 3782 37240 3834
rect 37252 3782 37304 3834
rect 37316 3782 37368 3834
rect 51504 3782 51556 3834
rect 51568 3782 51620 3834
rect 51632 3782 51684 3834
rect 51696 3782 51748 3834
rect 51760 3782 51812 3834
rect 4160 3612 4212 3664
rect 5356 3655 5408 3664
rect 5356 3621 5365 3655
rect 5365 3621 5399 3655
rect 5399 3621 5408 3655
rect 5356 3612 5408 3621
rect 5448 3612 5500 3664
rect 2136 3587 2188 3596
rect 2136 3553 2145 3587
rect 2145 3553 2179 3587
rect 2179 3553 2188 3587
rect 2136 3544 2188 3553
rect 3148 3544 3200 3596
rect 3240 3544 3292 3596
rect 4620 3544 4672 3596
rect 4804 3587 4856 3596
rect 4804 3553 4813 3587
rect 4813 3553 4847 3587
rect 4847 3553 4856 3587
rect 4804 3544 4856 3553
rect 4896 3544 4948 3596
rect 5080 3587 5132 3596
rect 5080 3553 5104 3587
rect 5104 3553 5132 3587
rect 5080 3544 5132 3553
rect 6736 3680 6788 3732
rect 6828 3680 6880 3732
rect 7104 3612 7156 3664
rect 8208 3612 8260 3664
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 13544 3680 13596 3732
rect 14096 3680 14148 3732
rect 3516 3476 3568 3528
rect 5908 3476 5960 3528
rect 7932 3544 7984 3596
rect 9036 3587 9088 3596
rect 9036 3553 9045 3587
rect 9045 3553 9079 3587
rect 9079 3553 9088 3587
rect 9036 3544 9088 3553
rect 9128 3544 9180 3596
rect 11244 3612 11296 3664
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 3424 3408 3476 3460
rect 7288 3451 7340 3460
rect 7288 3417 7297 3451
rect 7297 3417 7331 3451
rect 7331 3417 7340 3451
rect 7288 3408 7340 3417
rect 15752 3680 15804 3732
rect 16396 3680 16448 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 17868 3680 17920 3732
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 12808 3476 12860 3528
rect 11428 3408 11480 3460
rect 14004 3476 14056 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15200 3476 15252 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 20352 3612 20404 3664
rect 18788 3544 18840 3596
rect 19156 3544 19208 3596
rect 22284 3680 22336 3732
rect 16580 3476 16632 3528
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 4068 3340 4120 3392
rect 6920 3340 6972 3392
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 11336 3340 11388 3392
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12440 3340 12492 3349
rect 12716 3340 12768 3392
rect 19064 3476 19116 3528
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 20260 3476 20312 3528
rect 21088 3519 21140 3528
rect 21088 3485 21097 3519
rect 21097 3485 21131 3519
rect 21131 3485 21140 3519
rect 21088 3476 21140 3485
rect 21364 3476 21416 3528
rect 13912 3383 13964 3392
rect 13912 3349 13921 3383
rect 13921 3349 13955 3383
rect 13955 3349 13964 3383
rect 13912 3340 13964 3349
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 15200 3340 15252 3392
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 21456 3408 21508 3460
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 24768 3680 24820 3732
rect 26056 3680 26108 3732
rect 26700 3680 26752 3732
rect 28724 3723 28776 3732
rect 28724 3689 28733 3723
rect 28733 3689 28767 3723
rect 28767 3689 28776 3723
rect 28724 3680 28776 3689
rect 29460 3680 29512 3732
rect 30932 3680 30984 3732
rect 36084 3723 36136 3732
rect 36084 3689 36093 3723
rect 36093 3689 36127 3723
rect 36127 3689 36136 3723
rect 36084 3680 36136 3689
rect 36176 3723 36228 3732
rect 36176 3689 36185 3723
rect 36185 3689 36219 3723
rect 36219 3689 36228 3723
rect 36176 3680 36228 3689
rect 23020 3476 23072 3528
rect 24400 3476 24452 3528
rect 25228 3476 25280 3528
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 30104 3587 30156 3596
rect 30104 3553 30113 3587
rect 30113 3553 30147 3587
rect 30147 3553 30156 3587
rect 30104 3544 30156 3553
rect 31760 3612 31812 3664
rect 37832 3680 37884 3732
rect 37924 3680 37976 3732
rect 42156 3680 42208 3732
rect 42892 3723 42944 3732
rect 42892 3689 42901 3723
rect 42901 3689 42935 3723
rect 42935 3689 42944 3723
rect 42892 3680 42944 3689
rect 42984 3680 43036 3732
rect 32036 3544 32088 3596
rect 32496 3544 32548 3596
rect 33600 3544 33652 3596
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 17224 3340 17276 3349
rect 17684 3383 17736 3392
rect 17684 3349 17693 3383
rect 17693 3349 17727 3383
rect 17727 3349 17736 3383
rect 17684 3340 17736 3349
rect 18236 3340 18288 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 21548 3383 21600 3392
rect 21548 3349 21557 3383
rect 21557 3349 21591 3383
rect 21591 3349 21600 3383
rect 21548 3340 21600 3349
rect 22652 3340 22704 3392
rect 24124 3383 24176 3392
rect 24124 3349 24133 3383
rect 24133 3349 24167 3383
rect 24167 3349 24176 3383
rect 24124 3340 24176 3349
rect 24308 3408 24360 3460
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 25228 3340 25280 3392
rect 25780 3340 25832 3392
rect 26792 3383 26844 3392
rect 26792 3349 26801 3383
rect 26801 3349 26835 3383
rect 26835 3349 26844 3383
rect 26792 3340 26844 3349
rect 28540 3408 28592 3460
rect 29092 3408 29144 3460
rect 34520 3476 34572 3528
rect 38108 3587 38160 3596
rect 38108 3553 38117 3587
rect 38117 3553 38151 3587
rect 38151 3553 38160 3587
rect 38108 3544 38160 3553
rect 38384 3544 38436 3596
rect 38476 3544 38528 3596
rect 37648 3476 37700 3528
rect 38660 3476 38712 3528
rect 39948 3587 40000 3596
rect 39948 3553 39957 3587
rect 39957 3553 39991 3587
rect 39991 3553 40000 3587
rect 39948 3544 40000 3553
rect 40132 3587 40184 3596
rect 40132 3553 40141 3587
rect 40141 3553 40175 3587
rect 40175 3553 40184 3587
rect 40132 3544 40184 3553
rect 28264 3340 28316 3392
rect 29276 3340 29328 3392
rect 29368 3340 29420 3392
rect 29736 3340 29788 3392
rect 33232 3408 33284 3460
rect 37464 3408 37516 3460
rect 39396 3519 39448 3528
rect 39396 3485 39405 3519
rect 39405 3485 39439 3519
rect 39439 3485 39448 3519
rect 39396 3476 39448 3485
rect 42064 3612 42116 3664
rect 43076 3587 43128 3596
rect 43076 3553 43085 3587
rect 43085 3553 43119 3587
rect 43119 3553 43128 3587
rect 43076 3544 43128 3553
rect 45744 3680 45796 3732
rect 47860 3680 47912 3732
rect 48596 3680 48648 3732
rect 49056 3680 49108 3732
rect 44180 3544 44232 3596
rect 47768 3612 47820 3664
rect 45008 3544 45060 3596
rect 45100 3544 45152 3596
rect 45376 3544 45428 3596
rect 46848 3587 46900 3596
rect 46848 3553 46857 3587
rect 46857 3553 46891 3587
rect 46891 3553 46900 3587
rect 46848 3544 46900 3553
rect 47308 3544 47360 3596
rect 41972 3519 42024 3528
rect 41972 3485 41981 3519
rect 41981 3485 42015 3519
rect 42015 3485 42024 3519
rect 41972 3476 42024 3485
rect 41788 3408 41840 3460
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 43996 3476 44048 3528
rect 42892 3451 42944 3460
rect 42892 3417 42901 3451
rect 42901 3417 42935 3451
rect 42935 3417 42944 3451
rect 42892 3408 42944 3417
rect 43812 3408 43864 3460
rect 46204 3476 46256 3528
rect 47032 3519 47084 3528
rect 47032 3485 47050 3519
rect 47050 3485 47084 3519
rect 47032 3476 47084 3485
rect 48136 3519 48188 3528
rect 48136 3485 48145 3519
rect 48145 3485 48179 3519
rect 48179 3485 48188 3519
rect 48136 3476 48188 3485
rect 48872 3544 48924 3596
rect 51356 3680 51408 3732
rect 52000 3680 52052 3732
rect 53196 3680 53248 3732
rect 53932 3680 53984 3732
rect 55036 3680 55088 3732
rect 55220 3680 55272 3732
rect 49884 3544 49936 3596
rect 50344 3544 50396 3596
rect 50712 3519 50764 3528
rect 50712 3485 50721 3519
rect 50721 3485 50755 3519
rect 50755 3485 50764 3519
rect 50712 3476 50764 3485
rect 31116 3383 31168 3392
rect 31116 3349 31125 3383
rect 31125 3349 31159 3383
rect 31159 3349 31168 3383
rect 31116 3340 31168 3349
rect 31392 3383 31444 3392
rect 31392 3349 31401 3383
rect 31401 3349 31435 3383
rect 31435 3349 31444 3383
rect 31392 3340 31444 3349
rect 33508 3340 33560 3392
rect 35992 3340 36044 3392
rect 37556 3340 37608 3392
rect 39856 3340 39908 3392
rect 40684 3383 40736 3392
rect 40684 3349 40693 3383
rect 40693 3349 40727 3383
rect 40727 3349 40736 3383
rect 40684 3340 40736 3349
rect 43168 3340 43220 3392
rect 49424 3408 49476 3460
rect 50252 3408 50304 3460
rect 51908 3476 51960 3528
rect 52000 3519 52052 3528
rect 52000 3485 52009 3519
rect 52009 3485 52043 3519
rect 52043 3485 52052 3519
rect 52000 3476 52052 3485
rect 58532 3612 58584 3664
rect 57244 3544 57296 3596
rect 52828 3476 52880 3528
rect 54852 3519 54904 3528
rect 54852 3485 54861 3519
rect 54861 3485 54895 3519
rect 54895 3485 54904 3519
rect 54852 3476 54904 3485
rect 57060 3519 57112 3528
rect 57060 3485 57069 3519
rect 57069 3485 57103 3519
rect 57103 3485 57112 3519
rect 57060 3476 57112 3485
rect 57152 3519 57204 3528
rect 57152 3485 57161 3519
rect 57161 3485 57195 3519
rect 57195 3485 57204 3519
rect 57152 3476 57204 3485
rect 57888 3408 57940 3460
rect 44180 3340 44232 3392
rect 44824 3383 44876 3392
rect 44824 3349 44833 3383
rect 44833 3349 44867 3383
rect 44867 3349 44876 3383
rect 44824 3340 44876 3349
rect 45008 3383 45060 3392
rect 45008 3349 45017 3383
rect 45017 3349 45051 3383
rect 45051 3349 45060 3383
rect 45008 3340 45060 3349
rect 45652 3383 45704 3392
rect 45652 3349 45661 3383
rect 45661 3349 45695 3383
rect 45695 3349 45704 3383
rect 45652 3340 45704 3349
rect 46204 3340 46256 3392
rect 47492 3340 47544 3392
rect 48412 3340 48464 3392
rect 49700 3340 49752 3392
rect 51724 3340 51776 3392
rect 54116 3340 54168 3392
rect 15394 3238 15446 3290
rect 15458 3238 15510 3290
rect 15522 3238 15574 3290
rect 15586 3238 15638 3290
rect 15650 3238 15702 3290
rect 29838 3238 29890 3290
rect 29902 3238 29954 3290
rect 29966 3238 30018 3290
rect 30030 3238 30082 3290
rect 30094 3238 30146 3290
rect 44282 3238 44334 3290
rect 44346 3238 44398 3290
rect 44410 3238 44462 3290
rect 44474 3238 44526 3290
rect 44538 3238 44590 3290
rect 58726 3238 58778 3290
rect 58790 3238 58842 3290
rect 58854 3238 58906 3290
rect 58918 3238 58970 3290
rect 58982 3238 59034 3290
rect 1860 3179 1912 3188
rect 1860 3145 1869 3179
rect 1869 3145 1903 3179
rect 1903 3145 1912 3179
rect 1860 3136 1912 3145
rect 2136 3136 2188 3188
rect 4068 3136 4120 3188
rect 1768 3000 1820 3052
rect 3240 3000 3292 3052
rect 4344 3068 4396 3120
rect 4620 3136 4672 3188
rect 5264 3136 5316 3188
rect 5908 3136 5960 3188
rect 6368 3136 6420 3188
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 6920 3136 6972 3188
rect 7564 3179 7616 3188
rect 7564 3145 7573 3179
rect 7573 3145 7607 3179
rect 7607 3145 7616 3179
rect 7564 3136 7616 3145
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 2320 2932 2372 2984
rect 4988 2932 5040 2984
rect 5540 2864 5592 2916
rect 9772 3136 9824 3188
rect 10876 3136 10928 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 11704 3136 11756 3188
rect 14556 3136 14608 3188
rect 15844 3136 15896 3188
rect 17684 3136 17736 3188
rect 17960 3136 18012 3188
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 18328 3179 18380 3188
rect 18328 3145 18337 3179
rect 18337 3145 18371 3179
rect 18371 3145 18380 3179
rect 18328 3136 18380 3145
rect 18420 3136 18472 3188
rect 18788 3136 18840 3188
rect 20812 3136 20864 3188
rect 21548 3136 21600 3188
rect 21824 3136 21876 3188
rect 6460 3000 6512 3052
rect 7288 3000 7340 3052
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8208 3000 8260 3052
rect 9680 3068 9732 3120
rect 6644 2932 6696 2984
rect 10048 3000 10100 3052
rect 13820 3068 13872 3120
rect 11244 2932 11296 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 14096 3000 14148 3052
rect 21732 3068 21784 3120
rect 14924 3000 14976 3052
rect 18052 3000 18104 3052
rect 21456 3000 21508 3052
rect 22008 3000 22060 3052
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 15292 2932 15344 2984
rect 16212 2932 16264 2984
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 9036 2796 9088 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 12348 2839 12400 2848
rect 12348 2805 12357 2839
rect 12357 2805 12391 2839
rect 12391 2805 12400 2839
rect 12348 2796 12400 2805
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 14648 2796 14700 2848
rect 15016 2796 15068 2848
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 23020 3136 23072 3188
rect 24124 3136 24176 3188
rect 27252 3136 27304 3188
rect 27528 3136 27580 3188
rect 23020 3000 23072 3052
rect 23756 3000 23808 3052
rect 26240 3068 26292 3120
rect 29092 3179 29144 3188
rect 29092 3145 29101 3179
rect 29101 3145 29135 3179
rect 29135 3145 29144 3179
rect 29092 3136 29144 3145
rect 30840 3136 30892 3188
rect 31760 3136 31812 3188
rect 33508 3136 33560 3188
rect 28264 3068 28316 3120
rect 18604 2864 18656 2916
rect 20260 2864 20312 2916
rect 21548 2864 21600 2916
rect 23480 2932 23532 2984
rect 23572 2932 23624 2984
rect 24124 2932 24176 2984
rect 25780 2932 25832 2984
rect 27620 3000 27672 3052
rect 26608 2932 26660 2984
rect 29000 3000 29052 3052
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 29184 3000 29236 3009
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 29092 2932 29144 2984
rect 30196 2932 30248 2984
rect 33508 3043 33560 3052
rect 33508 3009 33517 3043
rect 33517 3009 33551 3043
rect 33551 3009 33560 3043
rect 33508 3000 33560 3009
rect 34612 3136 34664 3188
rect 36360 3136 36412 3188
rect 38476 3136 38528 3188
rect 40684 3136 40736 3188
rect 41604 3136 41656 3188
rect 41880 3136 41932 3188
rect 43076 3136 43128 3188
rect 43536 3136 43588 3188
rect 44732 3136 44784 3188
rect 45008 3136 45060 3188
rect 47216 3136 47268 3188
rect 48320 3136 48372 3188
rect 49424 3136 49476 3188
rect 50712 3136 50764 3188
rect 54024 3136 54076 3188
rect 54116 3179 54168 3188
rect 54116 3145 54125 3179
rect 54125 3145 54159 3179
rect 54159 3145 54168 3179
rect 54116 3136 54168 3145
rect 55956 3179 56008 3188
rect 55956 3145 55965 3179
rect 55965 3145 55999 3179
rect 55999 3145 56008 3179
rect 55956 3136 56008 3145
rect 35440 3000 35492 3052
rect 35624 3000 35676 3052
rect 35992 3000 36044 3052
rect 36360 3000 36412 3052
rect 22284 2839 22336 2848
rect 22284 2805 22293 2839
rect 22293 2805 22327 2839
rect 22327 2805 22336 2839
rect 22284 2796 22336 2805
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 32036 2864 32088 2916
rect 27712 2796 27764 2848
rect 31760 2796 31812 2848
rect 33508 2864 33560 2916
rect 35348 2975 35400 2984
rect 35348 2941 35357 2975
rect 35357 2941 35391 2975
rect 35391 2941 35400 2975
rect 35348 2932 35400 2941
rect 35716 2975 35768 2984
rect 35716 2941 35725 2975
rect 35725 2941 35759 2975
rect 35759 2941 35768 2975
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 38660 3000 38712 3052
rect 43352 3043 43404 3052
rect 43352 3009 43361 3043
rect 43361 3009 43395 3043
rect 43395 3009 43404 3043
rect 43352 3000 43404 3009
rect 43996 3000 44048 3052
rect 44088 3043 44140 3052
rect 44088 3009 44097 3043
rect 44097 3009 44131 3043
rect 44131 3009 44140 3043
rect 44088 3000 44140 3009
rect 44456 3000 44508 3052
rect 44640 3000 44692 3052
rect 44824 3111 44876 3120
rect 44824 3077 44858 3111
rect 44858 3077 44876 3111
rect 44824 3068 44876 3077
rect 45100 3068 45152 3120
rect 45284 3000 45336 3052
rect 46940 3000 46992 3052
rect 50344 3068 50396 3120
rect 53564 3068 53616 3120
rect 48872 3000 48924 3052
rect 49608 3000 49660 3052
rect 35716 2932 35768 2941
rect 37648 2932 37700 2984
rect 38476 2932 38528 2984
rect 34152 2796 34204 2848
rect 35992 2796 36044 2848
rect 36360 2796 36412 2848
rect 37464 2796 37516 2848
rect 40684 2932 40736 2984
rect 40132 2864 40184 2916
rect 45836 2932 45888 2984
rect 48044 2932 48096 2984
rect 50712 2932 50764 2984
rect 52368 3043 52420 3052
rect 52368 3009 52377 3043
rect 52377 3009 52411 3043
rect 52411 3009 52420 3043
rect 52368 3000 52420 3009
rect 52828 3000 52880 3052
rect 57520 3136 57572 3188
rect 57704 3136 57756 3188
rect 57888 3179 57940 3188
rect 57888 3145 57897 3179
rect 57897 3145 57931 3179
rect 57931 3145 57940 3179
rect 57888 3136 57940 3145
rect 54484 3000 54536 3052
rect 52552 2975 52604 2984
rect 52552 2941 52561 2975
rect 52561 2941 52595 2975
rect 52595 2941 52604 2975
rect 52552 2932 52604 2941
rect 53932 2932 53984 2984
rect 55036 2932 55088 2984
rect 57704 3043 57756 3052
rect 57704 3009 57713 3043
rect 57713 3009 57747 3043
rect 57747 3009 57756 3043
rect 57704 3000 57756 3009
rect 42248 2864 42300 2916
rect 40408 2796 40460 2848
rect 41972 2796 42024 2848
rect 43720 2839 43772 2848
rect 43720 2805 43729 2839
rect 43729 2805 43763 2839
rect 43763 2805 43772 2839
rect 43720 2796 43772 2805
rect 43996 2796 44048 2848
rect 45560 2796 45612 2848
rect 47032 2796 47084 2848
rect 48320 2839 48372 2848
rect 48320 2805 48329 2839
rect 48329 2805 48363 2839
rect 48363 2805 48372 2839
rect 48320 2796 48372 2805
rect 48412 2796 48464 2848
rect 52184 2864 52236 2916
rect 50252 2839 50304 2848
rect 50252 2805 50261 2839
rect 50261 2805 50295 2839
rect 50295 2805 50304 2839
rect 50252 2796 50304 2805
rect 53380 2796 53432 2848
rect 55404 2796 55456 2848
rect 57980 2864 58032 2916
rect 57428 2796 57480 2848
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 22616 2694 22668 2746
rect 22680 2694 22732 2746
rect 22744 2694 22796 2746
rect 22808 2694 22860 2746
rect 22872 2694 22924 2746
rect 37060 2694 37112 2746
rect 37124 2694 37176 2746
rect 37188 2694 37240 2746
rect 37252 2694 37304 2746
rect 37316 2694 37368 2746
rect 51504 2694 51556 2746
rect 51568 2694 51620 2746
rect 51632 2694 51684 2746
rect 51696 2694 51748 2746
rect 51760 2694 51812 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 7748 2592 7800 2644
rect 8024 2592 8076 2644
rect 9864 2592 9916 2644
rect 12440 2592 12492 2644
rect 14004 2592 14056 2644
rect 14280 2592 14332 2644
rect 17592 2592 17644 2644
rect 21548 2592 21600 2644
rect 21640 2592 21692 2644
rect 22376 2592 22428 2644
rect 23480 2592 23532 2644
rect 23756 2592 23808 2644
rect 26424 2592 26476 2644
rect 26884 2592 26936 2644
rect 27436 2635 27488 2644
rect 27436 2601 27445 2635
rect 27445 2601 27479 2635
rect 27479 2601 27488 2635
rect 27436 2592 27488 2601
rect 28632 2592 28684 2644
rect 29000 2592 29052 2644
rect 31392 2592 31444 2644
rect 33784 2592 33836 2644
rect 7564 2456 7616 2508
rect 9956 2456 10008 2508
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4896 2388 4948 2440
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 2044 2320 2096 2372
rect 5264 2363 5316 2372
rect 5264 2329 5273 2363
rect 5273 2329 5307 2363
rect 5307 2329 5316 2363
rect 5264 2320 5316 2329
rect 7012 2388 7064 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9772 2388 9824 2440
rect 20720 2524 20772 2576
rect 12164 2456 12216 2508
rect 12348 2388 12400 2440
rect 14188 2456 14240 2508
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 14556 2456 14608 2465
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 15844 2499 15896 2508
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 17868 2456 17920 2508
rect 13912 2388 13964 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17224 2388 17276 2440
rect 19432 2388 19484 2440
rect 20260 2388 20312 2440
rect 22468 2456 22520 2508
rect 22100 2388 22152 2440
rect 8392 2320 8444 2372
rect 14372 2320 14424 2372
rect 20720 2363 20772 2372
rect 20720 2329 20729 2363
rect 20729 2329 20763 2363
rect 20763 2329 20772 2363
rect 20720 2320 20772 2329
rect 22284 2320 22336 2372
rect 23204 2388 23256 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2388 25280 2440
rect 26792 2431 26844 2440
rect 26792 2397 26801 2431
rect 26801 2397 26835 2431
rect 26835 2397 26844 2431
rect 26792 2388 26844 2397
rect 27620 2456 27672 2508
rect 25780 2363 25832 2372
rect 25780 2329 25789 2363
rect 25789 2329 25823 2363
rect 25823 2329 25832 2363
rect 25780 2320 25832 2329
rect 27712 2431 27764 2440
rect 27712 2397 27721 2431
rect 27721 2397 27755 2431
rect 27755 2397 27764 2431
rect 27712 2388 27764 2397
rect 29736 2456 29788 2508
rect 30104 2499 30156 2508
rect 30104 2465 30113 2499
rect 30113 2465 30147 2499
rect 30147 2465 30156 2499
rect 30104 2456 30156 2465
rect 31116 2456 31168 2508
rect 35716 2592 35768 2644
rect 35992 2592 36044 2644
rect 37004 2592 37056 2644
rect 35440 2524 35492 2576
rect 43352 2592 43404 2644
rect 44456 2592 44508 2644
rect 45652 2592 45704 2644
rect 49792 2635 49844 2644
rect 49792 2601 49801 2635
rect 49801 2601 49835 2635
rect 49835 2601 49844 2635
rect 49792 2592 49844 2601
rect 51172 2592 51224 2644
rect 51908 2592 51960 2644
rect 55312 2592 55364 2644
rect 34428 2456 34480 2508
rect 35716 2456 35768 2508
rect 29276 2388 29328 2440
rect 31760 2431 31812 2440
rect 31760 2397 31769 2431
rect 31769 2397 31803 2431
rect 31803 2397 31812 2431
rect 31760 2388 31812 2397
rect 32036 2388 32088 2440
rect 7656 2252 7708 2304
rect 30748 2363 30800 2372
rect 30748 2329 30757 2363
rect 30757 2329 30791 2363
rect 30791 2329 30800 2363
rect 30748 2320 30800 2329
rect 28816 2252 28868 2304
rect 33232 2388 33284 2440
rect 34060 2388 34112 2440
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 35256 2388 35308 2440
rect 37096 2431 37148 2440
rect 37096 2397 37105 2431
rect 37105 2397 37139 2431
rect 37139 2397 37148 2431
rect 37096 2388 37148 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 32404 2320 32456 2372
rect 35624 2320 35676 2372
rect 35900 2252 35952 2304
rect 36820 2252 36872 2304
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 39856 2431 39908 2440
rect 39856 2397 39865 2431
rect 39865 2397 39899 2431
rect 39899 2397 39908 2431
rect 39856 2388 39908 2397
rect 39120 2320 39172 2372
rect 41328 2456 41380 2508
rect 40408 2388 40460 2440
rect 42248 2431 42300 2440
rect 42248 2397 42257 2431
rect 42257 2397 42291 2431
rect 42291 2397 42300 2431
rect 42248 2388 42300 2397
rect 43720 2431 43772 2440
rect 43720 2397 43729 2431
rect 43729 2397 43763 2431
rect 43763 2397 43772 2431
rect 43720 2388 43772 2397
rect 40592 2320 40644 2372
rect 42524 2320 42576 2372
rect 43444 2320 43496 2372
rect 44272 2388 44324 2440
rect 45560 2499 45612 2508
rect 45560 2465 45569 2499
rect 45569 2465 45603 2499
rect 45603 2465 45612 2499
rect 45560 2456 45612 2465
rect 43812 2252 43864 2304
rect 47032 2499 47084 2508
rect 47032 2465 47041 2499
rect 47041 2465 47075 2499
rect 47075 2465 47084 2499
rect 47032 2456 47084 2465
rect 49240 2456 49292 2508
rect 52000 2456 52052 2508
rect 52460 2456 52512 2508
rect 53748 2456 53800 2508
rect 48320 2388 48372 2440
rect 47308 2320 47360 2372
rect 46756 2252 46808 2304
rect 49700 2388 49752 2440
rect 50252 2431 50304 2440
rect 50252 2397 50261 2431
rect 50261 2397 50295 2431
rect 50295 2397 50304 2431
rect 50252 2388 50304 2397
rect 52184 2431 52236 2440
rect 52184 2397 52193 2431
rect 52193 2397 52227 2431
rect 52227 2397 52236 2431
rect 52184 2388 52236 2397
rect 51356 2320 51408 2372
rect 52736 2431 52788 2440
rect 52736 2397 52745 2431
rect 52745 2397 52779 2431
rect 52779 2397 52788 2431
rect 52736 2388 52788 2397
rect 55404 2456 55456 2508
rect 55772 2592 55824 2644
rect 57152 2635 57204 2644
rect 57152 2601 57161 2635
rect 57161 2601 57195 2635
rect 57195 2601 57204 2635
rect 57152 2592 57204 2601
rect 57704 2592 57756 2644
rect 55772 2456 55824 2508
rect 55680 2431 55732 2440
rect 55680 2397 55689 2431
rect 55689 2397 55723 2431
rect 55723 2397 55732 2431
rect 55680 2388 55732 2397
rect 57612 2456 57664 2508
rect 57980 2456 58032 2508
rect 57520 2431 57572 2440
rect 57520 2397 57529 2431
rect 57529 2397 57563 2431
rect 57563 2397 57572 2431
rect 57520 2388 57572 2397
rect 58348 2320 58400 2372
rect 50988 2252 51040 2304
rect 15394 2150 15446 2202
rect 15458 2150 15510 2202
rect 15522 2150 15574 2202
rect 15586 2150 15638 2202
rect 15650 2150 15702 2202
rect 29838 2150 29890 2202
rect 29902 2150 29954 2202
rect 29966 2150 30018 2202
rect 30030 2150 30082 2202
rect 30094 2150 30146 2202
rect 44282 2150 44334 2202
rect 44346 2150 44398 2202
rect 44410 2150 44462 2202
rect 44474 2150 44526 2202
rect 44538 2150 44590 2202
rect 58726 2150 58778 2202
rect 58790 2150 58842 2202
rect 58854 2150 58906 2202
rect 58918 2150 58970 2202
rect 58982 2150 59034 2202
rect 34612 2048 34664 2100
rect 39672 2048 39724 2100
rect 33048 1368 33100 1420
rect 37096 1368 37148 1420
<< metal2 >>
rect 15394 21788 15702 21797
rect 15394 21786 15400 21788
rect 15456 21786 15480 21788
rect 15536 21786 15560 21788
rect 15616 21786 15640 21788
rect 15696 21786 15702 21788
rect 15456 21734 15458 21786
rect 15638 21734 15640 21786
rect 15394 21732 15400 21734
rect 15456 21732 15480 21734
rect 15536 21732 15560 21734
rect 15616 21732 15640 21734
rect 15696 21732 15702 21734
rect 15394 21723 15702 21732
rect 29838 21788 30146 21797
rect 29838 21786 29844 21788
rect 29900 21786 29924 21788
rect 29980 21786 30004 21788
rect 30060 21786 30084 21788
rect 30140 21786 30146 21788
rect 29900 21734 29902 21786
rect 30082 21734 30084 21786
rect 29838 21732 29844 21734
rect 29900 21732 29924 21734
rect 29980 21732 30004 21734
rect 30060 21732 30084 21734
rect 30140 21732 30146 21734
rect 29838 21723 30146 21732
rect 44282 21788 44590 21797
rect 44282 21786 44288 21788
rect 44344 21786 44368 21788
rect 44424 21786 44448 21788
rect 44504 21786 44528 21788
rect 44584 21786 44590 21788
rect 44344 21734 44346 21786
rect 44526 21734 44528 21786
rect 44282 21732 44288 21734
rect 44344 21732 44368 21734
rect 44424 21732 44448 21734
rect 44504 21732 44528 21734
rect 44584 21732 44590 21734
rect 44282 21723 44590 21732
rect 58726 21788 59034 21797
rect 58726 21786 58732 21788
rect 58788 21786 58812 21788
rect 58868 21786 58892 21788
rect 58948 21786 58972 21788
rect 59028 21786 59034 21788
rect 58788 21734 58790 21786
rect 58970 21734 58972 21786
rect 58726 21732 58732 21734
rect 58788 21732 58812 21734
rect 58868 21732 58892 21734
rect 58948 21732 58972 21734
rect 59028 21732 59034 21734
rect 58726 21723 59034 21732
rect 38384 21548 38436 21554
rect 38384 21490 38436 21496
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 30748 21480 30800 21486
rect 30748 21422 30800 21428
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 32956 21480 33008 21486
rect 32956 21422 33008 21428
rect 33416 21480 33468 21486
rect 33416 21422 33468 21428
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4172 20398 4200 20742
rect 5000 20534 5028 21286
rect 5184 21010 5212 21286
rect 5644 21146 5672 21422
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 8680 21010 8708 21286
rect 8956 21146 8984 21286
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4264 19854 4292 20334
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18290 3556 19110
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2148 16590 2176 18158
rect 4172 17882 4200 19246
rect 4264 18290 4292 19790
rect 4448 19786 4476 20198
rect 4436 19780 4488 19786
rect 4436 19722 4488 19728
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4632 18970 4660 19246
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2148 16114 2176 16526
rect 2608 16182 2636 16934
rect 2976 16590 3004 17478
rect 3528 17338 3556 17614
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3252 16250 3280 17070
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16250 3832 16390
rect 3988 16250 4016 17206
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 14414 2176 16050
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2240 13938 2268 14758
rect 2700 14414 2728 15302
rect 3252 15162 3280 15438
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15162 3832 15302
rect 3988 15162 4016 16186
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 14006 2544 14214
rect 2884 14074 2912 14894
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2056 12986 2084 13874
rect 3528 13802 3556 14758
rect 3804 14074 3832 14758
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3988 13938 4016 15098
rect 4172 14958 4200 17682
rect 4448 17678 4476 18770
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 15978 4384 16526
rect 4632 16522 4660 17070
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14618 4200 14894
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4356 14482 4384 15438
rect 4724 14958 4752 18838
rect 5184 16998 5212 20946
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 5644 20058 5672 20878
rect 6564 20330 6592 20878
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 6552 20324 6604 20330
rect 6552 20266 6604 20272
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 18358 5304 19110
rect 6472 18970 6500 19246
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5828 18154 5856 18566
rect 6380 18290 6408 18702
rect 6472 18630 6500 18770
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5460 17746 5488 18022
rect 6380 17882 6408 18226
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5276 16674 5304 17070
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 5184 16646 5304 16674
rect 5184 16590 5212 16646
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4724 14074 4752 14894
rect 5080 14408 5132 14414
rect 5184 14396 5212 16526
rect 5460 16454 5488 16526
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5132 14368 5212 14396
rect 5080 14350 5132 14356
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4724 13870 4752 14010
rect 5276 14006 5304 15302
rect 5736 14958 5764 15302
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5368 14482 5396 14826
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 1872 12442 1900 12786
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 12442 3740 12582
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 4172 12238 4200 12786
rect 4448 12434 4476 12786
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 4264 12406 4476 12434
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3344 11150 3372 12038
rect 3620 11354 3648 12038
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2884 10266 2912 10610
rect 3160 10266 3188 10610
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 8430 2268 9590
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 7410 2268 8366
rect 2792 7886 2820 9998
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 3068 9722 3096 9930
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3252 9654 3280 11018
rect 3344 10538 3372 11086
rect 3896 10674 3924 11086
rect 3988 11082 4016 11630
rect 4172 11354 4200 12174
rect 4264 12102 4292 12406
rect 5184 12306 5212 12582
rect 5552 12442 5580 12718
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4264 11898 4292 12038
rect 4540 11898 4568 12038
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11354 4384 11494
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 11150 4384 11290
rect 4540 11234 4568 11698
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4448 11206 4568 11234
rect 4448 11150 4476 11206
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 4080 9654 4108 10610
rect 4264 10538 4292 10950
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3344 8498 3372 8910
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8566 3832 8774
rect 3896 8634 3924 9522
rect 4356 9178 4384 10610
rect 4448 10538 4476 11086
rect 4724 11014 4752 11630
rect 4816 11082 4844 11766
rect 5644 11762 5672 12174
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11150 4936 11494
rect 5000 11150 5028 11698
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4816 10810 4844 11018
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5644 10674 5672 10950
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 6914 2268 7346
rect 1964 6886 2268 6914
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1780 4826 1808 5646
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1780 4146 1808 4762
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 800 980 3431
rect 1688 3369 1716 3878
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1780 3058 1808 4082
rect 1858 3224 1914 3233
rect 1858 3159 1860 3168
rect 1912 3159 1914 3168
rect 1860 3130 1912 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1964 2650 1992 6886
rect 3344 6866 3372 8434
rect 3804 7886 3832 8502
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3896 8090 3924 8366
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3436 7002 3464 7414
rect 3712 7206 3740 7822
rect 3988 7410 4016 8026
rect 4356 7886 4384 8434
rect 4540 8362 4568 9318
rect 5000 9178 5028 9522
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8362 5396 8842
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7410 4108 7686
rect 4540 7478 4568 8298
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4724 7410 4752 7754
rect 5460 7750 5488 9522
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5552 9178 5580 9454
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5552 8974 5580 9114
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 8090 5580 8502
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3712 6662 3740 7142
rect 3988 6662 4016 7346
rect 4080 6730 4108 7346
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4356 6866 4384 7210
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4724 6798 4752 7346
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2700 5710 2728 6054
rect 2792 5710 2820 6054
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2700 5370 2728 5646
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4826 2636 4966
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 4214 2268 4422
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2976 4078 3004 5034
rect 3252 4690 3280 6054
rect 3344 5098 3372 6190
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5302 3556 6054
rect 3988 5914 4016 6122
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3160 4010 3188 4558
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3252 3720 3280 4626
rect 3528 4214 3556 5102
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4282 3648 4422
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3160 3692 3280 3720
rect 2134 3632 2190 3641
rect 3160 3602 3188 3692
rect 2134 3567 2136 3576
rect 2188 3567 2190 3576
rect 3148 3596 3200 3602
rect 2136 3538 2188 3544
rect 3148 3538 3200 3544
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 2148 3194 2176 3538
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 3252 3058 3280 3538
rect 3528 3534 3556 4150
rect 3792 4072 3844 4078
rect 3790 4040 3792 4049
rect 3844 4040 3846 4049
rect 3790 3975 3846 3984
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 1688 1170 1716 2314
rect 1504 1142 1716 1170
rect 1504 800 1532 1142
rect 2056 800 2084 2314
rect 2332 1578 2360 2926
rect 2332 1550 2636 1578
rect 2608 800 2636 1550
rect 3160 870 3280 898
rect 3160 800 3188 870
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3252 762 3280 870
rect 3436 762 3464 3402
rect 4080 3398 4108 6666
rect 4908 6662 4936 7278
rect 5092 6934 5120 7278
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5710 4476 6054
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4356 5370 4384 5510
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4826 4660 4966
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4252 4480 4304 4486
rect 4250 4448 4252 4457
rect 4344 4480 4396 4486
rect 4304 4448 4306 4457
rect 4344 4422 4396 4428
rect 4250 4383 4306 4392
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4172 3670 4200 4014
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3194 4108 3334
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3792 2440 3844 2446
rect 3712 2400 3792 2428
rect 3712 800 3740 2400
rect 3792 2382 3844 2388
rect 4264 800 4292 4082
rect 4356 3126 4384 4422
rect 4632 4282 4660 4558
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4908 3924 4936 6598
rect 5460 6322 5488 7686
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5030 5028 6190
rect 5460 5914 5488 6258
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5644 5386 5672 9522
rect 5736 6254 5764 14894
rect 5828 14074 5856 14962
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6012 12442 6040 16934
rect 6288 16726 6316 16934
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6288 16250 6316 16662
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6104 15162 6132 15302
rect 6196 15162 6224 15438
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6184 14544 6236 14550
rect 6288 14498 6316 16186
rect 6380 15162 6408 16730
rect 6472 15434 6500 18566
rect 7024 17678 7052 19314
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7116 18154 7144 18906
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7116 16998 7144 18090
rect 7300 17746 7328 19722
rect 7576 18222 7604 20334
rect 7668 20058 7696 20334
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7668 19514 7696 19722
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7760 19310 7788 20742
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8036 20330 8156 20346
rect 8036 20324 8168 20330
rect 8036 20318 8116 20324
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 8036 18970 8064 20318
rect 8116 20266 8168 20272
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8588 18766 8616 20538
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8772 20058 8800 20334
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 9048 19700 9076 20742
rect 9140 20602 9168 20878
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9128 19712 9180 19718
rect 9048 19672 9128 19700
rect 9128 19654 9180 19660
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7392 18086 7420 18158
rect 8680 18086 8708 19110
rect 8864 18358 8892 19246
rect 9140 18630 9168 19654
rect 9416 19242 9444 20946
rect 9508 20466 9536 21422
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9784 19854 9812 20742
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10152 20058 10180 20402
rect 10796 20398 10824 21014
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10888 20534 10916 20878
rect 10876 20528 10928 20534
rect 11060 20528 11112 20534
rect 10876 20470 10928 20476
rect 10980 20476 11060 20482
rect 10980 20470 11112 20476
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9876 19514 9904 19654
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 9140 18306 9168 18566
rect 9232 18426 9260 18566
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9140 18278 9260 18306
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 8680 17882 8708 18022
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 17338 7328 17682
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7300 16590 7328 17274
rect 8312 17202 8340 17478
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8680 17134 8708 17818
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 17270 9168 17682
rect 9232 17542 9260 18278
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7944 16590 7972 16934
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 8772 16590 8800 17070
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 7300 16114 7328 16526
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7484 16250 7512 16458
rect 8116 16448 8168 16454
rect 8036 16396 8116 16402
rect 8036 16390 8168 16396
rect 8036 16374 8156 16390
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6748 15706 6776 15982
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6564 14618 6592 14894
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6236 14492 6316 14498
rect 6184 14486 6316 14492
rect 6196 14470 6316 14486
rect 6656 14482 6684 15438
rect 7932 15360 7984 15366
rect 8036 15348 8064 16374
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 8864 15638 8892 15846
rect 8944 15700 8996 15706
rect 8996 15660 9076 15688
rect 8944 15642 8996 15648
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 7984 15320 8064 15348
rect 7932 15302 7984 15308
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6288 14278 6316 14470
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12986 6500 13262
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5828 10266 5856 10610
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 7886 5856 8434
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 6012 7546 6040 12378
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6288 11558 6316 12242
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6104 10198 6132 10542
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6564 10130 6592 14214
rect 6656 14074 6684 14418
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8498 6132 8774
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6104 7886 6132 8434
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6196 7546 6224 9386
rect 6288 9042 6316 9862
rect 6748 9654 6776 13874
rect 7116 13682 7144 14758
rect 6932 13654 7144 13682
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10062 6868 10406
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 9382 6868 9998
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8090 6316 8978
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6012 6390 6040 7482
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 6100 5764 6190
rect 5736 6072 5856 6100
rect 5552 5358 5672 5386
rect 5172 5296 5224 5302
rect 5170 5264 5172 5273
rect 5224 5264 5226 5273
rect 5170 5199 5226 5208
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 5000 4078 5028 4694
rect 5184 4554 5212 4966
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5184 4434 5212 4490
rect 5092 4282 5120 4422
rect 5184 4406 5396 4434
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 4908 3896 5028 3924
rect 4710 3768 4766 3777
rect 4710 3703 4766 3712
rect 4620 3596 4672 3602
rect 4724 3584 4752 3703
rect 4894 3632 4950 3641
rect 4804 3596 4856 3602
rect 4724 3556 4804 3584
rect 4620 3538 4672 3544
rect 4894 3567 4896 3576
rect 4804 3538 4856 3544
rect 4948 3567 4950 3576
rect 4896 3538 4948 3544
rect 4632 3194 4660 3538
rect 5000 3482 5028 3896
rect 5092 3602 5120 3946
rect 5368 3670 5396 4406
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4908 3454 5028 3482
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4908 2446 4936 3454
rect 5264 3188 5316 3194
rect 5460 3176 5488 3606
rect 5316 3148 5488 3176
rect 5264 3130 5316 3136
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5000 1578 5028 2926
rect 5552 2922 5580 5358
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5644 4214 5672 5238
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5644 4010 5672 4150
rect 5828 4078 5856 6072
rect 6012 5166 6040 6326
rect 6196 5914 6224 7482
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6182 5536 6238 5545
rect 6104 5494 6182 5522
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6104 4826 6132 5494
rect 6182 5471 6238 5480
rect 6380 5370 6408 6598
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6182 5128 6238 5137
rect 6182 5063 6238 5072
rect 6196 4826 6224 5063
rect 6380 4826 6408 5306
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5920 3534 5948 4558
rect 6104 4146 6132 4762
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 3194 5948 3470
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 6196 2446 6224 4014
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3194 6408 3878
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6472 3058 6500 6802
rect 6840 6662 6868 9318
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6840 5710 6868 5850
rect 6828 5704 6880 5710
rect 6748 5664 6828 5692
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6564 2774 6592 4558
rect 6748 3777 6776 5664
rect 6828 5646 6880 5652
rect 6932 4146 6960 13654
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12102 7144 13126
rect 7760 12434 7788 15098
rect 7944 13938 7972 15302
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14414 8064 14758
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8588 14006 8616 14894
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7760 12406 7972 12434
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7944 12050 7972 12406
rect 8036 12238 8064 12854
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 8680 12434 8708 14554
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 14074 8984 14214
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9048 12434 9076 15660
rect 9140 14074 9168 17206
rect 9232 17066 9260 17478
rect 9416 17338 9444 19178
rect 9508 17678 9536 19314
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9784 17882 9812 18226
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9416 16658 9444 17274
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9600 15366 9628 17818
rect 9692 17746 9720 17818
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 16726 9720 17478
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 14618 9628 15302
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9508 12434 9536 13942
rect 8680 12406 8800 12434
rect 9048 12406 9260 12434
rect 9508 12406 9628 12434
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8772 12102 8800 12406
rect 8760 12096 8812 12102
rect 7576 11762 7604 12038
rect 7760 11898 7788 12038
rect 7944 12022 8064 12050
rect 8760 12038 8812 12044
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 8036 11558 8064 12022
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9654 7696 9930
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7116 6866 7144 9522
rect 7760 9518 7788 10202
rect 7944 10062 7972 11494
rect 8036 10470 8064 11494
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8772 11218 8800 12038
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8772 10606 8800 11154
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10674 8892 10950
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8760 10600 8812 10606
rect 8956 10554 8984 11494
rect 9232 11234 9260 12406
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11762 9536 12038
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11354 9352 11494
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9232 11206 9352 11234
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8760 10542 8812 10548
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8588 10062 8616 10542
rect 8864 10526 8984 10554
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 7944 9586 7972 9998
rect 8864 9994 8892 10526
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8956 10062 8984 10406
rect 9048 10198 9076 10950
rect 9140 10266 9168 11086
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 9140 10062 9168 10202
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9654 8340 9862
rect 8680 9722 8708 9930
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 8680 9178 8708 9658
rect 8864 9518 8892 9930
rect 9140 9722 9168 9998
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9232 9518 9260 11018
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7760 8634 7788 8978
rect 8864 8906 8892 9454
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7760 8022 7788 8570
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7024 5710 7052 6190
rect 7116 5930 7144 6598
rect 7208 6118 7236 7278
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7116 5902 7236 5930
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7116 5234 7144 5714
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 4214 7144 4558
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6734 3768 6790 3777
rect 6840 3738 6868 4082
rect 6734 3703 6736 3712
rect 6788 3703 6790 3712
rect 6828 3732 6880 3738
rect 6736 3674 6788 3680
rect 6828 3674 6880 3680
rect 6920 3392 6972 3398
rect 6642 3360 6698 3369
rect 7024 3380 7052 4082
rect 7116 4078 7144 4150
rect 7208 4078 7236 5902
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7116 3670 7144 4014
rect 7104 3664 7156 3670
rect 7300 3641 7328 7278
rect 7392 7206 7420 7686
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5914 7420 6258
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 5030 7420 5306
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7104 3606 7156 3612
rect 7286 3632 7342 3641
rect 7286 3567 7342 3576
rect 7300 3466 7328 3567
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 6972 3352 7052 3380
rect 6920 3334 6972 3340
rect 6642 3295 6698 3304
rect 6656 3194 6684 3295
rect 6918 3224 6974 3233
rect 6644 3188 6696 3194
rect 6918 3159 6920 3168
rect 6644 3130 6696 3136
rect 6972 3159 6974 3168
rect 6920 3130 6972 3136
rect 6656 2990 6684 3130
rect 7300 3058 7328 3402
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6472 2746 6592 2774
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 4816 1550 5028 1578
rect 4816 800 4844 1550
rect 5276 1170 5304 2314
rect 5276 1142 5396 1170
rect 5368 800 5396 1142
rect 6472 800 6500 2746
rect 7392 2446 7420 4422
rect 7484 4162 7512 7686
rect 7760 7410 7788 7958
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8312 7342 8340 7822
rect 8116 7336 8168 7342
rect 8114 7304 8116 7313
rect 8300 7336 8352 7342
rect 8168 7304 8170 7313
rect 8300 7278 8352 7284
rect 8114 7239 8170 7248
rect 8496 7206 8524 7822
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7576 6390 7604 6802
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7576 4282 7604 5510
rect 7668 5250 7696 7142
rect 7760 6866 7788 7142
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 8588 6866 8616 8298
rect 8680 7886 8708 8434
rect 8772 8090 8800 8434
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 7478 8708 7822
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8772 7274 8800 8026
rect 8864 8022 8892 8842
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6458 8248 6734
rect 8588 6458 8616 6802
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 7760 5778 7788 6394
rect 8680 6338 8708 7142
rect 9140 6798 9168 9114
rect 9218 8936 9274 8945
rect 9218 8871 9220 8880
rect 9272 8871 9274 8880
rect 9220 8842 9272 8848
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8588 6310 8708 6338
rect 9048 6322 9076 6666
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6316 9088 6322
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5778 8064 6054
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7760 5370 7788 5714
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7668 5222 7788 5250
rect 7760 4690 7788 5222
rect 7852 5030 7880 5646
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7656 4208 7708 4214
rect 7484 4146 7604 4162
rect 7656 4150 7708 4156
rect 7484 4140 7616 4146
rect 7484 4134 7564 4140
rect 7484 3058 7512 4134
rect 7564 4082 7616 4088
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3194 7604 3878
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7024 800 7052 2382
rect 7576 800 7604 2450
rect 7668 2310 7696 4150
rect 7760 4146 7788 4490
rect 8036 4486 8064 5578
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7944 4282 7972 4422
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8312 4146 8340 4694
rect 8588 4146 8616 6310
rect 9036 6258 9088 6264
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5302 8708 5510
rect 8668 5296 8720 5302
rect 8772 5273 8800 5714
rect 8852 5296 8904 5302
rect 8668 5238 8720 5244
rect 8758 5264 8814 5273
rect 8852 5238 8904 5244
rect 8758 5199 8814 5208
rect 8772 4690 8800 5199
rect 8864 5137 8892 5238
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 8956 4826 8984 5170
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9048 4690 9076 4966
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9140 4486 9168 6598
rect 9128 4480 9180 4486
rect 9232 4457 9260 8842
rect 9324 5778 9352 11206
rect 9416 11014 9444 11698
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10266 9444 10950
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9416 10130 9444 10202
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9508 9654 9536 10610
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9508 9489 9536 9590
rect 9494 9480 9550 9489
rect 9494 9415 9550 9424
rect 9600 9058 9628 12406
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9692 11150 9720 11834
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10742 9720 11086
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 9926 9720 10678
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9416 9030 9628 9058
rect 9416 8362 9444 9030
rect 9784 8974 9812 17138
rect 9876 15706 9904 19450
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 14958 9904 15438
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14482 9904 14894
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 12850 9904 14214
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9968 12434 9996 17002
rect 10060 15162 10088 18770
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10244 17746 10272 18022
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 15502 10272 17682
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9968 12406 10088 12434
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9876 11354 9904 11630
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8566 9536 8774
rect 9600 8634 9628 8842
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9416 4826 9444 8298
rect 9508 7886 9536 8502
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7546 9628 7754
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6322 9628 7346
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9692 5914 9720 6734
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9784 4826 9812 8910
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9128 4422 9180 4428
rect 9218 4448 9274 4457
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7944 3194 7972 3538
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2650 7788 2790
rect 8036 2650 8064 3470
rect 8220 3058 8248 3606
rect 9048 3602 9076 4150
rect 9140 3942 9168 4422
rect 9274 4406 9352 4434
rect 9218 4383 9274 4392
rect 9324 4146 9352 4406
rect 9416 4282 9444 4762
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3602 9168 3878
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 9048 2854 9076 3538
rect 9692 3126 9720 4694
rect 9876 4282 9904 11018
rect 9968 10606 9996 11630
rect 10060 11286 10088 12406
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 10060 10266 10088 10610
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 6458 10088 9930
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10152 8498 10180 9007
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10152 8090 10180 8434
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10152 5710 10180 8026
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10244 6390 10272 6598
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10140 5364 10192 5370
rect 10244 5352 10272 5714
rect 10192 5324 10272 5352
rect 10140 5306 10192 5312
rect 10152 4282 10180 5306
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 3194 9812 3334
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 9784 2446 9812 2790
rect 9876 2650 9904 4082
rect 10048 3052 10100 3058
rect 10336 3040 10364 18838
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 17678 10456 18566
rect 10704 18358 10732 19110
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10796 16114 10824 20334
rect 10888 19854 10916 20470
rect 10980 20454 11100 20470
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10980 19514 11008 20454
rect 11532 19786 11560 21286
rect 11624 20602 11652 21286
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11256 18970 11284 19246
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18426 11100 18702
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11348 18086 11376 19246
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18766 11560 19110
rect 11716 18970 11744 20402
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12084 19990 12112 20334
rect 12176 20262 12204 21422
rect 13464 21146 13492 21422
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12268 20602 12296 20742
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12084 19334 12112 19926
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12084 19306 12296 19334
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11716 18426 11744 18906
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18426 12020 18566
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15502 10732 15846
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10888 15094 10916 16390
rect 11532 16250 11560 16526
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16250 11744 16390
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15162 11376 15982
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15706 11560 15846
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 14074 10640 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 11072 13870 11100 15030
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10428 12442 10456 13194
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10796 12374 10824 13806
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 11286 10824 12310
rect 11072 12306 11100 13126
rect 11164 12986 11192 13806
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 13326 11376 13670
rect 11624 13394 11652 16050
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15434 11836 15982
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11900 15162 11928 16050
rect 12176 16046 12204 16662
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 15162 12020 15302
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12850 11284 13126
rect 11348 12986 11376 13262
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11624 12782 11652 13330
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11898 11192 12038
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10796 8090 10824 11222
rect 11256 10742 11284 12582
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10810 11468 11086
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10810 11560 10950
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 9518 10916 10406
rect 11716 9674 11744 14894
rect 11900 14074 11928 15098
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11900 13734 11928 14010
rect 12176 13954 12204 15982
rect 12268 15094 12296 19306
rect 12452 17882 12480 19858
rect 12544 19718 12572 20878
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 19786 12664 20198
rect 12820 20058 12848 20878
rect 13188 20398 13216 20878
rect 13464 20466 13492 21082
rect 14844 21010 14872 21286
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14384 20602 14412 20742
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 13372 19786 13400 20334
rect 13648 20058 13676 20334
rect 13820 20324 13872 20330
rect 13740 20284 13820 20312
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19378 12572 19654
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12544 18086 12572 18702
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12544 17610 12572 18022
rect 12636 17678 12664 19722
rect 13740 19378 13768 20284
rect 13820 20266 13872 20272
rect 14096 20324 14148 20330
rect 14096 20266 14148 20272
rect 14108 20058 14136 20266
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18834 12940 19110
rect 13556 18970 13584 19246
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12728 16998 12756 18158
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12360 15586 12388 16526
rect 12716 16448 12768 16454
rect 12820 16436 12848 18566
rect 12912 16726 12940 18770
rect 13556 18630 13584 18906
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17338 13032 17546
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13188 17202 13216 18566
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13280 17678 13308 18226
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12768 16408 12848 16436
rect 12716 16390 12768 16396
rect 12728 16046 12756 16390
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12900 15904 12952 15910
rect 13004 15892 13032 16934
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16250 13308 16390
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13004 15864 13124 15892
rect 12900 15846 12952 15852
rect 12912 15688 12940 15846
rect 12912 15660 13032 15688
rect 12360 15570 12940 15586
rect 13004 15570 13032 15660
rect 12360 15564 12952 15570
rect 12360 15558 12900 15564
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 14550 12296 14894
rect 12360 14890 12388 15558
rect 12900 15506 12952 15512
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12728 15162 12756 15438
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 11992 13926 12204 13954
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13394 11928 13670
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10810 11836 11086
rect 11900 11014 11928 11290
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11992 9674 12020 13926
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13530 12112 13806
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12918 12204 13330
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 11716 9646 11836 9674
rect 11992 9646 12112 9674
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 8974 11100 9386
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10520 4622 10548 7686
rect 11072 6730 11100 7686
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11256 5778 11284 7482
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5370 11100 5510
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 11072 4486 11100 5102
rect 11164 4554 11192 5306
rect 11348 5166 11376 6122
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11440 5012 11468 8298
rect 11808 8294 11836 9646
rect 12084 9518 12112 9646
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11900 8974 11928 9454
rect 12084 9382 12112 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8498 11928 8910
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 6458 11652 7822
rect 11808 6662 11836 8026
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11716 6118 11744 6598
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5778 11744 6054
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11900 5574 11928 6258
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 5914 12020 6190
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5302 11928 5510
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11256 4984 11468 5012
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10600 4208 10652 4214
rect 10598 4176 10600 4185
rect 10652 4176 10654 4185
rect 10598 4111 10654 4120
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10612 3738 10640 3946
rect 11256 3942 11284 4984
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11440 4282 11468 4490
rect 11716 4486 11744 5102
rect 12084 5098 12112 9318
rect 12268 8974 12296 9862
rect 12360 9382 12388 14554
rect 12728 14074 12756 15098
rect 13004 15026 13032 15506
rect 13096 15026 13124 15864
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13188 14618 13216 15506
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12544 13326 12572 14010
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 13096 12850 13124 13330
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9178 12388 9318
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12176 8090 12204 8434
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6730 12296 6938
rect 12360 6934 12388 8842
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12452 6798 12480 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6254 12204 6598
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11532 3942 11560 4422
rect 11716 4282 11744 4422
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 11256 3670 11284 3878
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10100 3012 10364 3040
rect 10048 2994 10100 3000
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8404 1170 8432 2314
rect 8404 1142 8708 1170
rect 8680 800 8708 1142
rect 9232 800 9260 2382
rect 9968 1170 9996 2450
rect 10796 1850 10824 3470
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 3194 10916 3334
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11256 2990 11284 3606
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 3194 11376 3334
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 10796 1822 10916 1850
rect 9784 1142 9996 1170
rect 9784 800 9812 1142
rect 10888 800 10916 1822
rect 11440 800 11468 3402
rect 11532 3194 11560 3470
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3194 11744 3334
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 12084 2990 12112 5034
rect 12360 5030 12388 5646
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12176 4078 12204 4966
rect 12360 4146 12388 4966
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 1170 12204 2450
rect 12360 2446 12388 2790
rect 12452 2650 12480 3334
rect 12544 3058 12572 12310
rect 13280 12238 13308 13126
rect 13372 12306 13400 15302
rect 13464 13274 13492 17546
rect 13556 15450 13584 18566
rect 13740 18136 13768 19314
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18902 13952 19110
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13820 18148 13872 18154
rect 13740 18108 13820 18136
rect 13636 15564 13688 15570
rect 13740 15552 13768 18108
rect 13820 18090 13872 18096
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13832 15570 13860 16526
rect 13924 16250 13952 16526
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13688 15524 13768 15552
rect 13820 15564 13872 15570
rect 13636 15506 13688 15512
rect 13820 15506 13872 15512
rect 13556 15422 13676 15450
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 13394 13584 14350
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13464 13246 13584 13274
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12820 11354 12848 12106
rect 13464 11354 13492 12922
rect 13556 11830 13584 13246
rect 13648 12986 13676 15422
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14074 13768 14962
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10742 13952 11086
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 12990 10568 13046 10577
rect 12990 10503 12992 10512
rect 13044 10503 13046 10512
rect 12992 10474 13044 10480
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12820 9722 12848 9998
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13004 9586 13032 10474
rect 13372 10266 13400 10610
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 7886 12756 9454
rect 13004 8634 13032 9522
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13358 8528 13414 8537
rect 13464 8498 13492 8774
rect 13358 8463 13360 8472
rect 13412 8463 13414 8472
rect 13452 8492 13504 8498
rect 13360 8434 13412 8440
rect 13452 8434 13504 8440
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 7936 13032 8230
rect 13372 8090 13400 8434
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13084 7948 13136 7954
rect 13004 7908 13084 7936
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12820 5642 12848 5782
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12912 4078 12940 5782
rect 13004 4486 13032 7908
rect 13084 7890 13136 7896
rect 13556 6914 13584 8298
rect 13188 6886 13584 6914
rect 13084 6316 13136 6322
rect 13188 6304 13216 6886
rect 13136 6276 13216 6304
rect 13084 6258 13136 6264
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 5302 13400 5578
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12820 3534 12848 4014
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12728 2990 12756 3334
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2854 12848 3470
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11992 1142 12204 1170
rect 11992 800 12020 1142
rect 13096 800 13124 4490
rect 13464 4146 13492 6886
rect 13648 6186 13676 9318
rect 13832 9110 13860 9930
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13832 8362 13860 9046
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5846 13676 6122
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13740 5642 13768 7346
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13832 7002 13860 7278
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6934 13952 7278
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5166 13860 5510
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13636 4072 13688 4078
rect 13556 4020 13636 4026
rect 13556 4014 13688 4020
rect 13556 3998 13676 4014
rect 13556 3738 13584 3998
rect 13832 3992 13860 5102
rect 13924 4622 13952 6394
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14016 4214 14044 18634
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 17882 14136 18566
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14200 14618 14228 19178
rect 14476 18766 14504 20198
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 19514 14596 19654
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14844 19378 14872 20742
rect 15212 20602 15240 21422
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 15394 20700 15702 20709
rect 15394 20698 15400 20700
rect 15456 20698 15480 20700
rect 15536 20698 15560 20700
rect 15616 20698 15640 20700
rect 15696 20698 15702 20700
rect 15456 20646 15458 20698
rect 15638 20646 15640 20698
rect 15394 20644 15400 20646
rect 15456 20644 15480 20646
rect 15536 20644 15560 20646
rect 15616 20644 15640 20646
rect 15696 20644 15702 20646
rect 15394 20635 15702 20644
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15764 20058 15792 20946
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 16040 20602 16068 20742
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15948 19854 15976 20402
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19854 16160 20198
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15394 19612 15702 19621
rect 15394 19610 15400 19612
rect 15456 19610 15480 19612
rect 15536 19610 15560 19612
rect 15616 19610 15640 19612
rect 15696 19610 15702 19612
rect 15456 19558 15458 19610
rect 15638 19558 15640 19610
rect 15394 19556 15400 19558
rect 15456 19556 15480 19558
rect 15536 19556 15560 19558
rect 15616 19556 15640 19558
rect 15696 19556 15702 19558
rect 15394 19547 15702 19556
rect 15764 19514 15792 19722
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18426 14412 18566
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17746 14504 18158
rect 14936 17882 14964 18702
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14752 17338 14780 17682
rect 15304 17678 15332 19246
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15394 18524 15702 18533
rect 15394 18522 15400 18524
rect 15456 18522 15480 18524
rect 15536 18522 15560 18524
rect 15616 18522 15640 18524
rect 15696 18522 15702 18524
rect 15456 18470 15458 18522
rect 15638 18470 15640 18522
rect 15394 18468 15400 18470
rect 15456 18468 15480 18470
rect 15536 18468 15560 18470
rect 15616 18468 15640 18470
rect 15696 18468 15702 18470
rect 15394 18459 15702 18468
rect 15764 18358 15792 18566
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15948 18290 15976 19790
rect 17144 19310 17172 19858
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19514 17632 19722
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17788 19310 17816 20742
rect 18064 20534 18092 21286
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 18248 20058 18276 20742
rect 18616 20602 18644 21422
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18708 20398 18736 20742
rect 19168 20398 19196 21082
rect 22388 21078 22416 21286
rect 22616 21244 22924 21253
rect 22616 21242 22622 21244
rect 22678 21242 22702 21244
rect 22758 21242 22782 21244
rect 22838 21242 22862 21244
rect 22918 21242 22924 21244
rect 22678 21190 22680 21242
rect 22860 21190 22862 21242
rect 22616 21188 22622 21190
rect 22678 21188 22702 21190
rect 22758 21188 22782 21190
rect 22838 21188 22862 21190
rect 22918 21188 22924 21190
rect 22616 21179 22924 21188
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 20602 19288 20742
rect 19812 20602 19840 20878
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17746 16252 18022
rect 16960 17746 16988 18226
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 15394 17436 15702 17445
rect 15394 17434 15400 17436
rect 15456 17434 15480 17436
rect 15536 17434 15560 17436
rect 15616 17434 15640 17436
rect 15696 17434 15702 17436
rect 15456 17382 15458 17434
rect 15638 17382 15640 17434
rect 15394 17380 15400 17382
rect 15456 17380 15480 17382
rect 15536 17380 15560 17382
rect 15616 17380 15640 17382
rect 15696 17380 15702 17382
rect 15394 17371 15702 17380
rect 17420 17338 17448 17546
rect 14740 17332 14792 17338
rect 14660 17292 14740 17320
rect 14660 16046 14688 17292
rect 14740 17274 14792 17280
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17972 17202 18000 18838
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 17882 18092 18566
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17604 16726 17632 16934
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14752 15094 14780 16390
rect 14844 16250 14872 16390
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15212 15706 15240 16526
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 15394 16348 15702 16357
rect 15394 16346 15400 16348
rect 15456 16346 15480 16348
rect 15536 16346 15560 16348
rect 15616 16346 15640 16348
rect 15696 16346 15702 16348
rect 15456 16294 15458 16346
rect 15638 16294 15640 16346
rect 15394 16292 15400 16294
rect 15456 16292 15480 16294
rect 15536 16292 15560 16294
rect 15616 16292 15640 16294
rect 15696 16292 15702 16294
rect 15394 16283 15702 16292
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15706 15608 15846
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 16500 15502 16528 15982
rect 16868 15502 16896 16390
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15394 15260 15702 15269
rect 15394 15258 15400 15260
rect 15456 15258 15480 15260
rect 15536 15258 15560 15260
rect 15616 15258 15640 15260
rect 15696 15258 15702 15260
rect 15456 15206 15458 15258
rect 15638 15206 15640 15258
rect 15394 15204 15400 15206
rect 15456 15204 15480 15206
rect 15536 15204 15560 15206
rect 15616 15204 15640 15206
rect 15696 15204 15702 15206
rect 15394 15195 15702 15204
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 15764 14958 15792 15302
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 13394 14228 14554
rect 14936 13938 14964 14758
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12646 14136 13262
rect 14384 12918 14412 13806
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13394 14504 13670
rect 15212 13530 15240 13806
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14476 13190 14504 13330
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14108 12306 14136 12582
rect 14384 12442 14412 12854
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 10606 14136 11222
rect 14384 11082 14412 11494
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 5778 14136 7142
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 13912 4004 13964 4010
rect 13832 3964 13912 3992
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13648 800 13676 3878
rect 13832 3126 13860 3964
rect 13912 3946 13964 3952
rect 14108 3738 14136 4422
rect 14200 4026 14228 11018
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 7546 14320 8774
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14476 7410 14504 13126
rect 14752 12374 14780 13262
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12986 14872 13126
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14568 10810 14596 11630
rect 15120 11558 15148 13398
rect 15304 13326 15332 14214
rect 15394 14172 15702 14181
rect 15394 14170 15400 14172
rect 15456 14170 15480 14172
rect 15536 14170 15560 14172
rect 15616 14170 15640 14172
rect 15696 14170 15702 14172
rect 15456 14118 15458 14170
rect 15638 14118 15640 14170
rect 15394 14116 15400 14118
rect 15456 14116 15480 14118
rect 15536 14116 15560 14118
rect 15616 14116 15640 14118
rect 15696 14116 15702 14118
rect 15394 14107 15702 14116
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13530 15516 13874
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15394 13084 15702 13093
rect 15394 13082 15400 13084
rect 15456 13082 15480 13084
rect 15536 13082 15560 13084
rect 15616 13082 15640 13084
rect 15696 13082 15702 13084
rect 15456 13030 15458 13082
rect 15638 13030 15640 13082
rect 15394 13028 15400 13030
rect 15456 13028 15480 13030
rect 15536 13028 15560 13030
rect 15616 13028 15640 13030
rect 15696 13028 15702 13030
rect 15394 13019 15702 13028
rect 15764 12714 15792 13330
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 16132 12646 16160 13126
rect 16316 12850 16344 13330
rect 16960 12918 16988 14214
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15394 11996 15702 12005
rect 15394 11994 15400 11996
rect 15456 11994 15480 11996
rect 15536 11994 15560 11996
rect 15616 11994 15640 11996
rect 15696 11994 15702 11996
rect 15456 11942 15458 11994
rect 15638 11942 15640 11994
rect 15394 11940 15400 11942
rect 15456 11940 15480 11942
rect 15536 11940 15560 11942
rect 15616 11940 15640 11942
rect 15696 11940 15702 11942
rect 15394 11931 15702 11940
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14752 10130 14780 10678
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10266 14964 10610
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14740 10124 14792 10130
rect 14660 10084 14740 10112
rect 14660 8838 14688 10084
rect 14740 10066 14792 10072
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9178 14780 9454
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14844 8566 14872 9114
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14844 7954 14872 8502
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14936 7546 14964 8434
rect 15120 7954 15148 11494
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15394 10908 15702 10917
rect 15394 10906 15400 10908
rect 15456 10906 15480 10908
rect 15536 10906 15560 10908
rect 15616 10906 15640 10908
rect 15696 10906 15702 10908
rect 15456 10854 15458 10906
rect 15638 10854 15640 10906
rect 15394 10852 15400 10854
rect 15456 10852 15480 10854
rect 15536 10852 15560 10854
rect 15616 10852 15640 10854
rect 15696 10852 15702 10854
rect 15394 10843 15702 10852
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 10266 15424 10406
rect 15856 10266 15884 10474
rect 16040 10470 16068 12106
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9636 15332 9930
rect 15394 9820 15702 9829
rect 15394 9818 15400 9820
rect 15456 9818 15480 9820
rect 15536 9818 15560 9820
rect 15616 9818 15640 9820
rect 15696 9818 15702 9820
rect 15456 9766 15458 9818
rect 15638 9766 15640 9818
rect 15394 9764 15400 9766
rect 15456 9764 15480 9766
rect 15536 9764 15560 9766
rect 15616 9764 15640 9766
rect 15696 9764 15702 9766
rect 15394 9755 15702 9764
rect 15384 9648 15436 9654
rect 15304 9608 15384 9636
rect 15384 9590 15436 9596
rect 15292 9512 15344 9518
rect 15290 9480 15292 9489
rect 15344 9480 15346 9489
rect 15290 9415 15346 9424
rect 15396 8974 15424 9590
rect 16040 9586 16068 10406
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 9382 16068 9522
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15948 9178 15976 9318
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16040 9058 16068 9318
rect 15948 9030 16068 9058
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15394 8732 15702 8741
rect 15394 8730 15400 8732
rect 15456 8730 15480 8732
rect 15536 8730 15560 8732
rect 15616 8730 15640 8732
rect 15696 8730 15702 8732
rect 15456 8678 15458 8730
rect 15638 8678 15640 8730
rect 15394 8676 15400 8678
rect 15456 8676 15480 8678
rect 15536 8676 15560 8678
rect 15616 8676 15640 8678
rect 15696 8676 15702 8678
rect 15394 8667 15702 8676
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14292 6914 14320 7346
rect 14292 6886 14412 6914
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 6458 14320 6598
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14384 4570 14412 6886
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14844 6746 14872 7482
rect 15120 7342 15148 7890
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15212 7206 15240 7890
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15394 7644 15702 7653
rect 15394 7642 15400 7644
rect 15456 7642 15480 7644
rect 15536 7642 15560 7644
rect 15616 7642 15640 7644
rect 15696 7642 15702 7644
rect 15456 7590 15458 7642
rect 15638 7590 15640 7642
rect 15394 7588 15400 7590
rect 15456 7588 15480 7590
rect 15536 7588 15560 7590
rect 15616 7588 15640 7590
rect 15696 7588 15702 7590
rect 15394 7579 15702 7588
rect 15856 7410 15884 7686
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15948 6914 15976 9030
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15856 6886 15976 6914
rect 14752 6458 14780 6734
rect 14844 6718 14964 6746
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14476 5234 14504 5782
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14568 5574 14596 5646
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14384 4542 14504 4570
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4282 14412 4422
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14200 3998 14320 4026
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13924 2446 13952 3334
rect 14016 2650 14044 3470
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3058 14136 3334
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14200 2514 14228 3878
rect 14292 2650 14320 3998
rect 14476 3074 14504 4542
rect 14568 4486 14596 5510
rect 14660 5370 14688 5714
rect 14844 5710 14872 6598
rect 14936 5914 14964 6718
rect 15394 6556 15702 6565
rect 15394 6554 15400 6556
rect 15456 6554 15480 6556
rect 15536 6554 15560 6556
rect 15616 6554 15640 6556
rect 15696 6554 15702 6556
rect 15456 6502 15458 6554
rect 15638 6502 15640 6554
rect 15394 6500 15400 6502
rect 15456 6500 15480 6502
rect 15536 6500 15560 6502
rect 15616 6500 15640 6502
rect 15696 6500 15702 6502
rect 15394 6491 15702 6500
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15764 5642 15792 6190
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15394 5468 15702 5477
rect 15394 5466 15400 5468
rect 15456 5466 15480 5468
rect 15536 5466 15560 5468
rect 15616 5466 15640 5468
rect 15696 5466 15702 5468
rect 15456 5414 15458 5466
rect 15638 5414 15640 5466
rect 15394 5412 15400 5414
rect 15456 5412 15480 5414
rect 15536 5412 15560 5414
rect 15616 5412 15640 5414
rect 15696 5412 15702 5414
rect 15394 5403 15702 5412
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 3194 14596 4422
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14832 3528 14884 3534
rect 14752 3488 14832 3516
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14384 3046 14504 3074
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14384 2378 14412 3046
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14200 870 14320 898
rect 14200 800 14228 870
rect 3252 734 3464 762
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14292 762 14320 870
rect 14476 762 14504 2926
rect 14568 2514 14596 3130
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14660 2514 14688 2790
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14752 800 14780 3488
rect 14832 3470 14884 3476
rect 14936 3058 14964 3878
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 15028 2854 15056 3878
rect 15212 3534 15240 4694
rect 15856 4690 15884 6886
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 5778 15976 6598
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15948 5030 15976 5714
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15304 4214 15332 4490
rect 15394 4380 15702 4389
rect 15394 4378 15400 4380
rect 15456 4378 15480 4380
rect 15536 4378 15560 4380
rect 15616 4378 15640 4380
rect 15696 4378 15702 4380
rect 15456 4326 15458 4378
rect 15638 4326 15640 4378
rect 15394 4324 15400 4326
rect 15456 4324 15480 4326
rect 15536 4324 15560 4326
rect 15616 4324 15640 4326
rect 15696 4324 15702 4326
rect 15394 4315 15702 4324
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15396 3534 15424 4014
rect 15764 3738 15792 4490
rect 15856 4282 15884 4626
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15948 4078 15976 4966
rect 16040 4826 16068 7142
rect 16132 5370 16160 12582
rect 16316 10266 16344 12582
rect 16408 11830 16436 12582
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 9654 16252 9998
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16316 9382 16344 10202
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 5710 16344 9318
rect 16408 6914 16436 11766
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11218 16620 11494
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16500 10130 16528 11154
rect 16684 11150 16712 12786
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16868 11898 16896 12174
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16684 10606 16712 11086
rect 16776 10674 16804 11698
rect 17052 10742 17080 12038
rect 17144 10810 17172 14826
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 14074 17264 14350
rect 17604 14278 17632 16662
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17696 15162 17724 16594
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 16250 17816 16390
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 18064 15706 18092 16526
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17604 13870 17632 14214
rect 17788 14074 17816 14214
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 11354 17356 11630
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17604 11014 17632 13806
rect 18248 13802 18276 18770
rect 18708 18766 18736 20334
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18340 18426 18368 18566
rect 18432 18426 18460 18566
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18708 18358 18736 18702
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18800 18426 18828 18566
rect 19076 18426 19104 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18340 16998 18368 18158
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18340 15706 18368 15846
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18432 14958 18460 15302
rect 18708 15162 18736 15506
rect 18800 15162 18828 16594
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19076 15638 19104 15914
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18892 15026 18920 15506
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 19168 14958 19196 20334
rect 19812 20330 19840 20538
rect 19800 20324 19852 20330
rect 19800 20266 19852 20272
rect 20088 19854 20116 20878
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20548 20466 20576 20538
rect 21468 20466 21496 20742
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17972 13394 18000 13670
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 18156 13326 18184 13670
rect 18248 13394 18276 13738
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18248 12434 18276 13330
rect 18340 12986 18368 14350
rect 18432 14278 18460 14894
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 14074 18460 14214
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 18616 13530 18644 13806
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18432 12918 18460 13194
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18248 12406 18644 12434
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 17236 10130 17264 10950
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17604 10130 17632 10746
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 16684 9518 16712 10066
rect 17788 9994 17816 10610
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17052 9586 17080 9862
rect 17512 9586 17540 9862
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16684 8974 16712 9454
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16592 8634 16620 8910
rect 16960 8838 16988 9454
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16592 7954 16620 8570
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16592 7410 16620 7482
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16408 6886 16528 6914
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16408 5914 16436 6190
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16132 4486 16160 4966
rect 16224 4622 16252 5578
rect 16500 5234 16528 6886
rect 16684 6798 16712 7142
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6322 16712 6734
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16776 6458 16804 6598
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15212 2446 15240 3334
rect 15394 3292 15702 3301
rect 15394 3290 15400 3292
rect 15456 3290 15480 3292
rect 15536 3290 15560 3292
rect 15616 3290 15640 3292
rect 15696 3290 15702 3292
rect 15456 3238 15458 3290
rect 15638 3238 15640 3290
rect 15394 3236 15400 3238
rect 15456 3236 15480 3238
rect 15536 3236 15560 3238
rect 15616 3236 15640 3238
rect 15696 3236 15702 3238
rect 15394 3227 15702 3236
rect 15856 3194 15884 3470
rect 16028 3392 16080 3398
rect 16026 3360 16028 3369
rect 16080 3360 16082 3369
rect 16026 3295 16082 3304
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 16224 2990 16252 4558
rect 16684 4554 16712 4966
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16408 3738 16436 4218
rect 16868 4010 16896 8298
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 17052 3534 17080 9318
rect 17788 8634 17816 9930
rect 18064 9654 18092 11018
rect 18340 10470 18368 11698
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18616 9382 18644 12406
rect 18708 12170 18736 13466
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19076 12850 19104 12922
rect 19260 12850 19288 13806
rect 19352 13530 19380 19246
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19720 18834 19748 19178
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19904 18222 19932 19654
rect 19984 18828 20036 18834
rect 20088 18816 20116 19790
rect 20364 19718 20392 20334
rect 20640 20058 20668 20334
rect 20812 20324 20864 20330
rect 20732 20284 20812 20312
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20732 19718 20760 20284
rect 20812 20266 20864 20272
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20036 18788 20116 18816
rect 19984 18770 20036 18776
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19628 17338 19656 17614
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19904 17270 19932 18158
rect 20272 17882 20300 18634
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18290 20392 18566
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20548 17746 20576 18158
rect 20732 18154 20760 19654
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18834 21220 19110
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 17882 20760 18090
rect 20720 17876 20772 17882
rect 20640 17836 20720 17864
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16250 19748 16934
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13530 19472 13806
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19340 13184 19392 13190
rect 19536 13138 19564 13330
rect 19628 13326 19656 15302
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19340 13126 19392 13132
rect 19352 12986 19380 13126
rect 19444 13110 19564 13138
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18708 10470 18736 12106
rect 19352 12102 19380 12922
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18984 10810 19012 11086
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 9450 19288 10406
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17328 7954 17356 8230
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17788 7886 17816 8570
rect 17972 8090 18000 8842
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8498 18736 8774
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 7410 17816 7822
rect 18144 7812 18196 7818
rect 18144 7754 18196 7760
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6458 17356 6598
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17236 4282 17264 5102
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17420 3738 17448 7346
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6866 18000 7142
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17788 5914 17816 6666
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17972 5234 18000 5714
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17512 4282 17540 4966
rect 18064 4554 18092 5102
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17880 3738 17908 3946
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 16580 3528 16632 3534
rect 16408 3488 16580 3516
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15304 800 15332 2926
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15394 2204 15702 2213
rect 15394 2202 15400 2204
rect 15456 2202 15480 2204
rect 15536 2202 15560 2204
rect 15616 2202 15640 2204
rect 15696 2202 15702 2204
rect 15456 2150 15458 2202
rect 15638 2150 15640 2202
rect 15394 2148 15400 2150
rect 15456 2148 15480 2150
rect 15536 2148 15560 2150
rect 15616 2148 15640 2150
rect 15696 2148 15702 2150
rect 15394 2139 15702 2148
rect 15856 800 15884 2450
rect 16408 800 16436 3488
rect 16580 3470 16632 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 2446 17264 3334
rect 17604 2650 17632 3470
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 3194 17724 3334
rect 17972 3194 18000 4082
rect 18156 3942 18184 7754
rect 18984 7342 19012 7890
rect 19168 7750 19196 8366
rect 19260 8362 19288 9386
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19352 8022 19380 12038
rect 19444 11762 19472 13110
rect 19524 12436 19576 12442
rect 19628 12434 19656 13126
rect 19720 12832 19748 16186
rect 19904 16114 19932 17206
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 15366 19840 15846
rect 19904 15502 19932 16050
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20180 15570 20208 15982
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 14958 19840 15302
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19800 12844 19852 12850
rect 19720 12804 19800 12832
rect 19800 12786 19852 12792
rect 19904 12714 19932 15438
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 14618 20024 14758
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20088 14074 20116 14962
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 12986 20208 13262
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19628 12406 19840 12434
rect 19524 12378 19576 12384
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19536 11354 19564 12378
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19628 10266 19656 11154
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19628 9722 19656 10202
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19628 9178 19656 9658
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18248 6914 18276 7278
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18340 7018 18368 7142
rect 18340 6990 18552 7018
rect 18248 6886 18460 6914
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 5778 18368 6598
rect 18432 6322 18460 6886
rect 18524 6458 18552 6990
rect 19168 6848 19196 7686
rect 19444 7410 19472 8230
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19248 6860 19300 6866
rect 19168 6820 19248 6848
rect 19248 6802 19300 6808
rect 19340 6724 19392 6730
rect 19536 6712 19564 7346
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19392 6684 19564 6712
rect 19340 6666 19392 6672
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6458 18828 6598
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 19536 6322 19564 6684
rect 19628 6458 19656 6802
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19720 6458 19748 6598
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18708 5846 18736 6190
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 19444 5574 19472 5850
rect 19536 5574 19564 6258
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18524 4622 18552 4966
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 3194 18276 3334
rect 18340 3194 18368 3470
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 3194 18460 3334
rect 18800 3194 18828 3538
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17788 2514 17908 2530
rect 17788 2508 17920 2514
rect 17788 2502 17868 2508
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 16960 800 16988 2382
rect 17512 870 17632 898
rect 17512 800 17540 870
rect 14292 734 14504 762
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 17604 762 17632 870
rect 17788 762 17816 2502
rect 17868 2450 17920 2456
rect 18064 800 18092 2994
rect 18892 2990 18920 4422
rect 18984 4146 19012 5034
rect 19260 4826 19288 5102
rect 19444 5098 19472 5510
rect 19812 5234 19840 12406
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19996 11898 20024 12106
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20272 11830 20300 12854
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11082 20300 11494
rect 20364 11354 20392 16934
rect 20640 16250 20668 17836
rect 20720 17818 20772 17824
rect 20824 17678 20852 18702
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20916 18426 20944 18566
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 15638 20668 16186
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20732 15094 20760 16390
rect 20824 16250 20852 17614
rect 20916 17202 20944 18362
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20720 14408 20772 14414
rect 20640 14356 20720 14362
rect 20640 14350 20772 14356
rect 20640 14334 20760 14350
rect 20640 14074 20668 14334
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20640 12986 20668 14010
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20640 12238 20668 12718
rect 20824 12442 20852 12718
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20640 11626 20668 12174
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 19982 10704 20038 10713
rect 20364 10690 20392 11290
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 19982 10639 19984 10648
rect 20036 10639 20038 10648
rect 20088 10674 20484 10690
rect 20088 10668 20496 10674
rect 20088 10662 20444 10668
rect 19984 10610 20036 10616
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19904 6390 19932 6802
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 19904 5846 19932 6326
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19904 5370 19932 5782
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19260 4146 19288 4490
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19076 3534 19104 4014
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18616 800 18644 2858
rect 19168 800 19196 3538
rect 19352 3534 19380 4966
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4078 19472 4422
rect 19628 4282 19656 4490
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19904 4010 19932 5306
rect 20088 4826 20116 10662
rect 20444 10610 20496 10616
rect 20732 10198 20760 10950
rect 20824 10810 20852 11630
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20916 10266 20944 17138
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 14278 21036 15302
rect 21100 15162 21128 16050
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21008 13326 21036 14214
rect 21100 13326 21128 14214
rect 21192 13394 21220 18770
rect 21376 18290 21404 20198
rect 21468 19922 21496 20402
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21560 19854 21588 20742
rect 22112 20602 22140 20878
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22388 20398 22416 21014
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 21744 20058 21772 20334
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 22296 19446 22324 20334
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 21916 18760 21968 18766
rect 21744 18720 21916 18748
rect 21744 18630 21772 18720
rect 21916 18702 21968 18708
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21836 18426 21864 18566
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 22112 18222 22140 18838
rect 22296 18766 22324 19382
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21284 17542 21312 18158
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 17338 21772 17478
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 15706 21404 16526
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 15162 21496 15438
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21192 12646 21220 13330
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 7868 20484 8910
rect 21192 8498 21220 12582
rect 21836 12434 21864 18022
rect 22112 17678 22140 18158
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22204 17610 22232 18566
rect 22388 18306 22416 20334
rect 22480 19446 22508 20878
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 22616 20156 22924 20165
rect 22616 20154 22622 20156
rect 22678 20154 22702 20156
rect 22758 20154 22782 20156
rect 22838 20154 22862 20156
rect 22918 20154 22924 20156
rect 22678 20102 22680 20154
rect 22860 20102 22862 20154
rect 22616 20100 22622 20102
rect 22678 20100 22702 20102
rect 22758 20100 22782 20102
rect 22838 20100 22862 20102
rect 22918 20100 22924 20102
rect 22616 20091 22924 20100
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19514 22600 19654
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 23492 19310 23520 20334
rect 23584 20058 23612 20402
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23676 19514 23704 20742
rect 24596 20482 24624 20946
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 24676 20800 24728 20806
rect 24728 20760 24808 20788
rect 24676 20742 24728 20748
rect 24674 20496 24730 20505
rect 24596 20454 24674 20482
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 22480 19156 22508 19246
rect 22836 19168 22888 19174
rect 22480 19128 22836 19156
rect 22836 19110 22888 19116
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 22616 19068 22924 19077
rect 22616 19066 22622 19068
rect 22678 19066 22702 19068
rect 22758 19066 22782 19068
rect 22838 19066 22862 19068
rect 22918 19066 22924 19068
rect 22678 19014 22680 19066
rect 22860 19014 22862 19066
rect 22616 19012 22622 19014
rect 22678 19012 22702 19014
rect 22758 19012 22782 19014
rect 22838 19012 22862 19014
rect 22918 19012 22924 19014
rect 22616 19003 22924 19012
rect 22388 18278 22508 18306
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22388 17338 22416 18158
rect 22376 17332 22428 17338
rect 22296 17292 22376 17320
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 21744 12406 21864 12434
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11150 21312 11494
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21456 10192 21508 10198
rect 21560 10146 21588 10950
rect 21508 10140 21588 10146
rect 21456 10134 21588 10140
rect 21468 10118 21588 10134
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21376 9654 21404 9862
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20536 7880 20588 7886
rect 20456 7840 20536 7868
rect 20536 7822 20588 7828
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20640 7546 20668 7686
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20824 7478 20852 7822
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 21284 7206 21312 7822
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 6322 20300 6802
rect 20456 6798 20484 6938
rect 21376 6934 21404 7414
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20456 5914 20484 6734
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20824 5914 20852 6258
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5030 20300 5510
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20272 4554 20300 4966
rect 20456 4826 20484 5850
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 20272 3534 20300 4490
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 20548 4010 20576 4150
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20364 3670 20392 3946
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20272 2922 20300 3470
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20732 2582 20760 5102
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 4146 20852 4558
rect 20916 4282 20944 6598
rect 21376 6322 21404 6870
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21100 5642 21128 6054
rect 21192 5778 21220 6054
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 21376 5574 21404 6258
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5370 21404 5510
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21376 4690 21404 5306
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20824 3194 20852 4082
rect 21100 3534 21128 4422
rect 21468 3942 21496 9998
rect 21560 7290 21588 10118
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 7478 21680 8230
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21560 7262 21680 7290
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21560 5098 21588 7142
rect 21652 6186 21680 7262
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21364 3528 21416 3534
rect 21560 3482 21588 5034
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21364 3470 21416 3476
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 17604 734 17816 762
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19444 762 19472 2382
rect 19628 870 19748 898
rect 19628 762 19656 870
rect 19720 800 19748 870
rect 20272 800 20300 2382
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 1170 20760 2314
rect 20732 1142 20852 1170
rect 20824 800 20852 1142
rect 21376 800 21404 3470
rect 21468 3466 21588 3482
rect 21456 3460 21588 3466
rect 21508 3454 21588 3460
rect 21456 3402 21508 3408
rect 21468 3058 21496 3402
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 3194 21588 3334
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21548 2916 21600 2922
rect 21548 2858 21600 2864
rect 21560 2650 21588 2858
rect 21652 2650 21680 4082
rect 21744 3126 21772 12406
rect 22020 12306 22048 15914
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15570 22140 15846
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22296 14074 22324 17292
rect 22376 17274 22428 17280
rect 22480 15026 22508 18278
rect 22616 17980 22924 17989
rect 22616 17978 22622 17980
rect 22678 17978 22702 17980
rect 22758 17978 22782 17980
rect 22838 17978 22862 17980
rect 22918 17978 22924 17980
rect 22678 17926 22680 17978
rect 22860 17926 22862 17978
rect 22616 17924 22622 17926
rect 22678 17924 22702 17926
rect 22758 17924 22782 17926
rect 22838 17924 22862 17926
rect 22918 17924 22924 17926
rect 22616 17915 22924 17924
rect 22616 16892 22924 16901
rect 22616 16890 22622 16892
rect 22678 16890 22702 16892
rect 22758 16890 22782 16892
rect 22838 16890 22862 16892
rect 22918 16890 22924 16892
rect 22678 16838 22680 16890
rect 22860 16838 22862 16890
rect 22616 16836 22622 16838
rect 22678 16836 22702 16838
rect 22758 16836 22782 16838
rect 22838 16836 22862 16838
rect 22918 16836 22924 16838
rect 22616 16827 22924 16836
rect 23400 16726 23428 19110
rect 23492 18222 23520 19246
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23584 18426 23612 18566
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23492 17746 23520 18158
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23768 16794 23796 19858
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23860 17542 23888 17818
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23400 15910 23428 16662
rect 23768 16046 23796 16730
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 22616 15804 22924 15813
rect 22616 15802 22622 15804
rect 22678 15802 22702 15804
rect 22758 15802 22782 15804
rect 22838 15802 22862 15804
rect 22918 15802 22924 15804
rect 22678 15750 22680 15802
rect 22860 15750 22862 15802
rect 22616 15748 22622 15750
rect 22678 15748 22702 15750
rect 22758 15748 22782 15750
rect 22838 15748 22862 15750
rect 22918 15748 22924 15750
rect 22616 15739 22924 15748
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22388 14618 22416 14894
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22480 14414 22508 14962
rect 22616 14716 22924 14725
rect 22616 14714 22622 14716
rect 22678 14714 22702 14716
rect 22758 14714 22782 14716
rect 22838 14714 22862 14716
rect 22918 14714 22924 14716
rect 22678 14662 22680 14714
rect 22860 14662 22862 14714
rect 22616 14660 22622 14662
rect 22678 14660 22702 14662
rect 22758 14660 22782 14662
rect 22838 14660 22862 14662
rect 22918 14660 22924 14662
rect 22616 14651 22924 14660
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11898 21864 12038
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 22020 9897 22048 12242
rect 22112 12170 22140 13670
rect 22296 13462 22324 14010
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22388 13530 22416 13806
rect 22616 13628 22924 13637
rect 22616 13626 22622 13628
rect 22678 13626 22702 13628
rect 22758 13626 22782 13628
rect 22838 13626 22862 13628
rect 22918 13626 22924 13628
rect 22678 13574 22680 13626
rect 22860 13574 22862 13626
rect 22616 13572 22622 13574
rect 22678 13572 22702 13574
rect 22758 13572 22782 13574
rect 22838 13572 22862 13574
rect 22918 13572 22924 13574
rect 22616 13563 22924 13572
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22204 12434 22232 12650
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 22616 12540 22924 12549
rect 22616 12538 22622 12540
rect 22678 12538 22702 12540
rect 22758 12538 22782 12540
rect 22838 12538 22862 12540
rect 22918 12538 22924 12540
rect 22678 12486 22680 12538
rect 22860 12486 22862 12538
rect 22616 12484 22622 12486
rect 22678 12484 22702 12486
rect 22758 12484 22782 12486
rect 22838 12484 22862 12486
rect 22918 12484 22924 12486
rect 22616 12475 22924 12484
rect 22204 12406 22416 12434
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22112 11642 22140 12106
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11898 22324 12038
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22112 11626 22324 11642
rect 22112 11620 22336 11626
rect 22112 11614 22284 11620
rect 22112 11354 22140 11614
rect 22284 11562 22336 11568
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22388 10810 22416 12406
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 11286 22508 11630
rect 23216 11558 23244 12582
rect 23400 12434 23428 15846
rect 23492 15502 23520 15846
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23584 12986 23612 13126
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23400 12406 23612 12434
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23492 11898 23520 12038
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23584 11694 23612 12406
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 22616 11452 22924 11461
rect 22616 11450 22622 11452
rect 22678 11450 22702 11452
rect 22758 11450 22782 11452
rect 22838 11450 22862 11452
rect 22918 11450 22924 11452
rect 22678 11398 22680 11450
rect 22860 11398 22862 11450
rect 22616 11396 22622 11398
rect 22678 11396 22702 11398
rect 22758 11396 22782 11398
rect 22838 11396 22862 11398
rect 22918 11396 22924 11398
rect 22616 11387 22924 11396
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 23216 11150 23244 11494
rect 23584 11218 23612 11630
rect 23676 11558 23704 13126
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23676 11082 23704 11494
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22112 10130 22140 10746
rect 22480 10606 22508 11018
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22616 10364 22924 10373
rect 22616 10362 22622 10364
rect 22678 10362 22702 10364
rect 22758 10362 22782 10364
rect 22838 10362 22862 10364
rect 22918 10362 22924 10364
rect 22678 10310 22680 10362
rect 22860 10310 22862 10362
rect 22616 10308 22622 10310
rect 22678 10308 22702 10310
rect 22758 10308 22782 10310
rect 22838 10308 22862 10310
rect 22918 10308 22924 10310
rect 22616 10299 22924 10308
rect 23032 10266 23060 10406
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22006 9888 22062 9897
rect 22006 9823 22062 9832
rect 22112 9722 22140 10066
rect 22284 10056 22336 10062
rect 23676 10010 23704 10610
rect 23768 10470 23796 15098
rect 23940 14816 23992 14822
rect 23992 14764 24072 14770
rect 23940 14758 24072 14764
rect 23952 14742 24072 14758
rect 24044 14346 24072 14742
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 24044 13938 24072 14282
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24136 13326 24164 16934
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24228 16250 24256 16390
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24320 15978 24348 16526
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24320 15706 24348 15914
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24412 15094 24440 16390
rect 24596 15570 24624 20454
rect 24674 20431 24730 20440
rect 24780 19718 24808 20760
rect 25056 20058 25084 20810
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25240 19786 25268 20878
rect 25608 20466 25636 21286
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25884 20602 25912 20878
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25884 20466 25912 20538
rect 27264 20534 27292 21286
rect 27816 21146 27844 21422
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 28092 21146 28120 21286
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27908 20534 27936 20810
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24780 18630 24808 19654
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 17134 24808 18566
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24872 16250 24900 17478
rect 25056 17338 25084 17546
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24688 15570 24716 16050
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24596 15162 24624 15506
rect 24964 15434 24992 15846
rect 25056 15706 25084 16526
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24584 15156 24636 15162
rect 24584 15098 24636 15104
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 14074 24900 14214
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12986 24808 13126
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 11898 24072 12174
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24320 11762 24348 12038
rect 24412 11898 24440 12038
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23952 10674 23980 11154
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 22284 9998 22336 10004
rect 22190 9888 22246 9897
rect 22190 9823 22246 9832
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8634 21864 8842
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21928 6798 21956 9454
rect 22112 9178 22140 9454
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21928 4622 21956 4966
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22020 4146 22048 7142
rect 22204 5302 22232 9823
rect 22296 9518 22324 9998
rect 23492 9982 23704 10010
rect 23492 9586 23520 9982
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 8634 22508 9318
rect 22616 9276 22924 9285
rect 22616 9274 22622 9276
rect 22678 9274 22702 9276
rect 22758 9274 22782 9276
rect 22838 9274 22862 9276
rect 22918 9274 22924 9276
rect 22678 9222 22680 9274
rect 22860 9222 22862 9274
rect 22616 9220 22622 9222
rect 22678 9220 22702 9222
rect 22758 9220 22782 9222
rect 22838 9220 22862 9222
rect 22918 9220 22924 9222
rect 22616 9211 22924 9220
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23216 8634 23244 8842
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23492 8430 23520 9522
rect 23584 8498 23612 9862
rect 23768 9178 23796 9862
rect 24136 9518 24164 10542
rect 24320 9994 24348 11698
rect 24504 11354 24532 12106
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24504 10606 24532 11290
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24308 9988 24360 9994
rect 24308 9930 24360 9936
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24412 9518 24440 9862
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23952 9110 23980 9454
rect 23940 9104 23992 9110
rect 23940 9046 23992 9052
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 22616 8188 22924 8197
rect 22616 8186 22622 8188
rect 22678 8186 22702 8188
rect 22758 8186 22782 8188
rect 22838 8186 22862 8188
rect 22918 8186 22924 8188
rect 22678 8134 22680 8186
rect 22860 8134 22862 8186
rect 22616 8132 22622 8134
rect 22678 8132 22702 8134
rect 22758 8132 22782 8134
rect 22838 8132 22862 8134
rect 22918 8132 22924 8134
rect 22616 8123 22924 8132
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22296 6390 22324 7958
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 23032 7410 23060 7686
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22616 7100 22924 7109
rect 22616 7098 22622 7100
rect 22678 7098 22702 7100
rect 22758 7098 22782 7100
rect 22838 7098 22862 7100
rect 22918 7098 22924 7100
rect 22678 7046 22680 7098
rect 22860 7046 22862 7098
rect 22616 7044 22622 7046
rect 22678 7044 22702 7046
rect 22758 7044 22782 7046
rect 22838 7044 22862 7046
rect 22918 7044 22924 7046
rect 22616 7035 22924 7044
rect 23584 7002 23612 7822
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23676 6866 23704 8366
rect 24044 8294 24072 8910
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24044 7750 24072 8230
rect 24136 8022 24164 9454
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7410 24072 7686
rect 24136 7478 24164 7958
rect 24124 7472 24176 7478
rect 24124 7414 24176 7420
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23768 6866 23796 7142
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22296 5914 22324 6326
rect 22480 5914 22508 6666
rect 23676 6186 23704 6802
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23952 6390 23980 6598
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23664 6180 23716 6186
rect 23664 6122 23716 6128
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22616 6012 22924 6021
rect 22616 6010 22622 6012
rect 22678 6010 22702 6012
rect 22758 6010 22782 6012
rect 22838 6010 22862 6012
rect 22918 6010 22924 6012
rect 22678 5958 22680 6010
rect 22860 5958 22862 6010
rect 22616 5956 22622 5958
rect 22678 5956 22702 5958
rect 22758 5956 22782 5958
rect 22838 5956 22862 5958
rect 22918 5956 22924 5958
rect 22616 5947 22924 5956
rect 23032 5914 23060 6054
rect 22284 5908 22336 5914
rect 22284 5850 22336 5856
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5574 22968 5714
rect 22928 5568 22980 5574
rect 22928 5510 22980 5516
rect 23952 5302 23980 6326
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 23940 5296 23992 5302
rect 23940 5238 23992 5244
rect 22616 4924 22924 4933
rect 22616 4922 22622 4924
rect 22678 4922 22702 4924
rect 22758 4922 22782 4924
rect 22838 4922 22862 4924
rect 22918 4922 22924 4924
rect 22678 4870 22680 4922
rect 22860 4870 22862 4922
rect 22616 4868 22622 4870
rect 22678 4868 22702 4870
rect 22758 4868 22782 4870
rect 22838 4868 22862 4870
rect 22918 4868 22924 4870
rect 22616 4859 22924 4868
rect 23952 4486 23980 5238
rect 24044 4690 24072 5646
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24136 4826 24164 5170
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24228 4826 24256 4966
rect 24320 4826 24348 6802
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24032 4684 24084 4690
rect 24032 4626 24084 4632
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24412 4570 24440 6598
rect 24596 5846 24624 11630
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24780 10674 24808 11290
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24872 10130 24900 12310
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24964 11694 24992 12174
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24964 10674 24992 11630
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 25148 10266 25176 17070
rect 25240 13802 25268 18702
rect 25608 18222 25636 20402
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25792 19718 25820 20334
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 19514 25820 19654
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 26160 19310 26188 20266
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25884 18222 25912 18566
rect 26160 18222 26188 19246
rect 26252 18766 26280 20198
rect 26988 19786 27016 20198
rect 27724 20058 27752 20402
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 26976 19780 27028 19786
rect 26976 19722 27028 19728
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 25608 17882 25636 18158
rect 25792 17882 25820 18158
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25608 17218 25636 17818
rect 25792 17678 25820 17818
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 26160 17610 26188 18158
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25884 17338 25912 17478
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25516 17202 25636 17218
rect 25504 17196 25636 17202
rect 25556 17190 25636 17196
rect 25504 17138 25556 17144
rect 25608 16658 25636 17190
rect 26252 16776 26280 18566
rect 26988 18306 27016 19722
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27264 18834 27292 19110
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27080 18426 27108 18566
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 26988 18278 27108 18306
rect 27080 18222 27108 18278
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27080 17746 27108 18158
rect 27068 17740 27120 17746
rect 27068 17682 27120 17688
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26620 16794 26648 17274
rect 26160 16748 26280 16776
rect 26608 16788 26660 16794
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25516 15706 25544 15982
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25516 15162 25544 15642
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25608 15026 25636 16390
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25792 15162 25820 16050
rect 25964 15564 26016 15570
rect 25964 15506 26016 15512
rect 25976 15450 26004 15506
rect 25976 15422 26096 15450
rect 25780 15156 25832 15162
rect 25780 15098 25832 15104
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25424 14074 25452 14350
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 14074 25636 14214
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25792 13938 25820 15098
rect 26068 15026 26096 15422
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 26068 14278 26096 14962
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 25792 13394 25820 13874
rect 26068 13530 26096 14214
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25780 13388 25832 13394
rect 25832 13348 25912 13376
rect 25780 13330 25832 13336
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12782 25820 13126
rect 25884 12986 25912 13348
rect 26160 13002 26188 16748
rect 26608 16730 26660 16736
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26252 16130 26280 16594
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26344 16250 26372 16526
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26252 16102 26372 16130
rect 26344 15570 26372 16102
rect 26620 16046 26648 16730
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26620 15502 26648 15846
rect 26896 15638 26924 17546
rect 26884 15632 26936 15638
rect 26936 15592 27016 15620
rect 26884 15574 26936 15580
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26620 14074 26648 15302
rect 26712 15162 26740 15302
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26332 13388 26384 13394
rect 26252 13348 26332 13376
rect 26252 13190 26280 13348
rect 26332 13330 26384 13336
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 25872 12980 25924 12986
rect 26160 12974 26280 13002
rect 26620 12986 26648 13262
rect 25872 12922 25924 12928
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25792 11898 25820 12718
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25884 12102 25912 12582
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25516 10810 25544 11630
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25240 10198 25268 10678
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25424 10470 25452 10542
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25228 10192 25280 10198
rect 25228 10134 25280 10140
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24688 9110 24716 9318
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 25240 8922 25268 10134
rect 24860 8900 24912 8906
rect 25240 8894 25360 8922
rect 24860 8842 24912 8848
rect 24872 8786 24900 8842
rect 24780 8758 24900 8786
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24688 7002 24716 7414
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24780 6322 24808 8758
rect 25240 8634 25268 8774
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25332 8022 25360 8894
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 25424 7834 25452 10406
rect 25700 9994 25728 10542
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25700 9042 25728 9930
rect 25884 9042 25912 12038
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26160 11082 26188 11494
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 25884 8430 25912 8978
rect 26068 8634 26096 9522
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25780 8016 25832 8022
rect 25780 7958 25832 7964
rect 25332 7806 25452 7834
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24872 6866 24900 7210
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 25056 6118 25084 6734
rect 25148 6662 25176 6734
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6458 25176 6598
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25332 6390 25360 7806
rect 25792 7002 25820 7958
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24780 5216 24808 5578
rect 24860 5228 24912 5234
rect 24780 5188 24860 5216
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24688 4690 24716 5102
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23940 4480 23992 4486
rect 23940 4422 23992 4428
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21836 3194 21864 3946
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21732 3120 21784 3126
rect 21732 3062 21784 3068
rect 22020 3058 22048 4082
rect 22296 3738 22324 4082
rect 22616 3836 22924 3845
rect 22616 3834 22622 3836
rect 22678 3834 22702 3836
rect 22758 3834 22782 3836
rect 22838 3834 22862 3836
rect 22918 3834 22924 3836
rect 22678 3782 22680 3834
rect 22860 3782 22862 3834
rect 22616 3780 22622 3782
rect 22678 3780 22702 3782
rect 22758 3780 22782 3782
rect 22838 3780 22862 3782
rect 22918 3780 22924 3782
rect 22616 3771 22924 3780
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 23492 3602 23520 4422
rect 23952 4214 23980 4422
rect 24320 4282 24348 4558
rect 24412 4542 24532 4570
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4282 24440 4422
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 24504 4078 24532 4542
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22008 3052 22060 3058
rect 22664 3040 22692 3334
rect 23032 3194 23060 3470
rect 24320 3466 24348 3878
rect 24412 3534 24440 3878
rect 24780 3738 24808 5188
rect 24860 5170 24912 5176
rect 25056 4622 25084 6054
rect 25332 5642 25360 6326
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 25608 5234 25636 5646
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 25240 3534 25268 4966
rect 25332 4690 25360 4966
rect 25700 4758 25728 6802
rect 25884 5846 25912 8366
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25976 7546 26004 7686
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 6458 26096 6734
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 25872 5840 25924 5846
rect 25872 5782 25924 5788
rect 25780 5568 25832 5574
rect 25780 5510 25832 5516
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25792 4078 25820 5510
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 26068 4010 26096 4558
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 26068 3738 26096 3946
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 25240 3398 25268 3470
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 24136 3194 24164 3334
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 23020 3052 23072 3058
rect 22664 3012 23020 3040
rect 22008 2994 22060 3000
rect 23020 2994 23072 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22112 1442 22140 2382
rect 22296 2378 22324 2790
rect 22388 2650 22416 2790
rect 22616 2748 22924 2757
rect 22616 2746 22622 2748
rect 22678 2746 22702 2748
rect 22758 2746 22782 2748
rect 22838 2746 22862 2748
rect 22918 2746 22924 2748
rect 22678 2694 22680 2746
rect 22860 2694 22862 2746
rect 22616 2692 22622 2694
rect 22678 2692 22702 2694
rect 22758 2692 22782 2694
rect 22838 2692 22862 2694
rect 22918 2692 22924 2694
rect 22616 2683 22924 2692
rect 23492 2650 23520 2926
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 23032 2502 23244 2530
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 21928 1414 22140 1442
rect 21928 800 21956 1414
rect 22480 800 22508 2450
rect 23032 800 23060 2502
rect 23216 2446 23244 2502
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23584 800 23612 2926
rect 23768 2650 23796 2994
rect 25792 2990 25820 3334
rect 26252 3126 26280 12974
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26528 11898 26556 12106
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26620 11558 26648 12106
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11218 26648 11494
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26712 11098 26740 14758
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26804 13938 26832 14350
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26804 13326 26832 13874
rect 26988 13462 27016 15592
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26988 12238 27016 13398
rect 27068 12708 27120 12714
rect 27068 12650 27120 12656
rect 27080 12238 27108 12650
rect 27264 12442 27292 18566
rect 27448 18358 27476 19110
rect 27908 18698 27936 20470
rect 28092 19854 28120 20742
rect 28368 20602 28396 21422
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28644 20602 28672 20878
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29644 20800 29696 20806
rect 29644 20742 29696 20748
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 29012 20398 29040 20742
rect 28908 20392 28960 20398
rect 28908 20334 28960 20340
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28172 20324 28224 20330
rect 28172 20266 28224 20272
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 28000 18970 28028 19246
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 28184 17338 28212 20266
rect 28920 20058 28948 20334
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 29656 19854 29684 20742
rect 29838 20700 30146 20709
rect 29838 20698 29844 20700
rect 29900 20698 29924 20700
rect 29980 20698 30004 20700
rect 30060 20698 30084 20700
rect 30140 20698 30146 20700
rect 29900 20646 29902 20698
rect 30082 20646 30084 20698
rect 29838 20644 29844 20646
rect 29900 20644 29924 20646
rect 29980 20644 30004 20646
rect 30060 20644 30084 20646
rect 30140 20644 30146 20646
rect 29838 20635 30146 20644
rect 30760 20602 30788 21422
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 31392 21344 31444 21350
rect 31392 21286 31444 21292
rect 31312 21010 31340 21286
rect 31300 21004 31352 21010
rect 31300 20946 31352 20952
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30196 20528 30248 20534
rect 30196 20470 30248 20476
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28276 18766 28304 19110
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28276 17678 28304 18566
rect 28552 18426 28580 19246
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28540 18420 28592 18426
rect 28540 18362 28592 18368
rect 28736 18358 28764 18634
rect 28828 18426 28856 18702
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28724 18352 28776 18358
rect 28724 18294 28776 18300
rect 28920 18086 28948 18702
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18426 29592 18566
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29748 18290 29776 19790
rect 29838 19612 30146 19621
rect 29838 19610 29844 19612
rect 29900 19610 29924 19612
rect 29980 19610 30004 19612
rect 30060 19610 30084 19612
rect 30140 19610 30146 19612
rect 29900 19558 29902 19610
rect 30082 19558 30084 19610
rect 29838 19556 29844 19558
rect 29900 19556 29924 19558
rect 29980 19556 30004 19558
rect 30060 19556 30084 19558
rect 30140 19556 30146 19558
rect 29838 19547 30146 19556
rect 29838 18524 30146 18533
rect 29838 18522 29844 18524
rect 29900 18522 29924 18524
rect 29980 18522 30004 18524
rect 30060 18522 30084 18524
rect 30140 18522 30146 18524
rect 29900 18470 29902 18522
rect 30082 18470 30084 18522
rect 29838 18468 29844 18470
rect 29900 18468 29924 18470
rect 29980 18468 30004 18470
rect 30060 18468 30084 18470
rect 30140 18468 30146 18470
rect 29838 18459 30146 18468
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 28908 18080 28960 18086
rect 28908 18022 28960 18028
rect 28920 17882 28948 18022
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 29196 17542 29224 18158
rect 29748 17746 29776 18226
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 28356 16040 28408 16046
rect 28356 15982 28408 15988
rect 27540 15502 27568 15982
rect 27804 15904 27856 15910
rect 27804 15846 27856 15852
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27816 15162 27844 15846
rect 28368 15706 28396 15982
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27540 13530 27568 13806
rect 27816 13530 27844 13806
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27356 12442 27384 12718
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27344 12436 27396 12442
rect 27344 12378 27396 12384
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 26528 11070 26740 11098
rect 26528 10674 26556 11070
rect 26700 11008 26752 11014
rect 26700 10950 26752 10956
rect 26712 10810 26740 10950
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 27448 10742 27476 12582
rect 27632 11762 27660 12922
rect 27816 12306 27844 13262
rect 27908 12850 27936 14962
rect 28356 14068 28408 14074
rect 28356 14010 28408 14016
rect 28172 13728 28224 13734
rect 28172 13670 28224 13676
rect 28184 12986 28212 13670
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27804 12300 27856 12306
rect 27804 12242 27856 12248
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 27632 10606 27660 10950
rect 27908 10742 27936 10950
rect 27896 10736 27948 10742
rect 27896 10678 27948 10684
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 26884 10192 26936 10198
rect 26884 10134 26936 10140
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 26620 9042 26648 9318
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26700 8356 26752 8362
rect 26700 8298 26752 8304
rect 26712 7886 26740 8298
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26528 7002 26556 7822
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 26620 6866 26648 7210
rect 26792 7200 26844 7206
rect 26792 7142 26844 7148
rect 26804 6866 26832 7142
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26528 4826 26556 6258
rect 26712 5710 26740 6666
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26516 4820 26568 4826
rect 26516 4762 26568 4768
rect 26608 4616 26660 4622
rect 26436 4576 26608 4604
rect 26332 4548 26384 4554
rect 26332 4490 26384 4496
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 24136 800 24164 2926
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24596 1306 24624 2382
rect 24596 1278 24716 1306
rect 24688 800 24716 1278
rect 25240 800 25268 2382
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 25792 800 25820 2314
rect 26344 800 26372 4490
rect 26436 2650 26464 4576
rect 26608 4558 26660 4564
rect 26712 3942 26740 5646
rect 26896 4570 26924 10134
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 26988 5370 27016 5646
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 26988 4690 27016 5306
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26896 4542 27016 4570
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26712 3738 26740 3878
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26792 3392 26844 3398
rect 26792 3334 26844 3340
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26424 2644 26476 2650
rect 26424 2586 26476 2592
rect 19444 734 19656 762
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26620 762 26648 2926
rect 26804 2446 26832 3334
rect 26896 2650 26924 4422
rect 26988 3534 27016 4542
rect 27080 3942 27108 9998
rect 27632 9382 27660 10542
rect 27988 10192 28040 10198
rect 27988 10134 28040 10140
rect 27712 9920 27764 9926
rect 27710 9888 27712 9897
rect 27764 9888 27766 9897
rect 27710 9823 27766 9832
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27632 8906 27660 9318
rect 27724 8974 27752 9454
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 27620 8900 27672 8906
rect 27620 8842 27672 8848
rect 27632 8430 27660 8842
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27632 7750 27660 8366
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27632 7206 27660 7686
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27172 6322 27200 6598
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27632 6118 27660 7142
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27632 5574 27660 6054
rect 27816 5710 27844 6802
rect 27804 5704 27856 5710
rect 27804 5646 27856 5652
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 27356 4214 27384 5238
rect 27632 5166 27660 5510
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27632 4826 27660 5102
rect 27816 5030 27844 5646
rect 28000 5370 28028 10134
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 28092 9654 28120 9862
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 27988 5364 28040 5370
rect 27988 5306 28040 5312
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27724 4826 27752 4966
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27632 4282 27660 4762
rect 28276 4622 28304 5510
rect 28368 4622 28396 14010
rect 28736 12646 28764 17478
rect 29838 17436 30146 17445
rect 29838 17434 29844 17436
rect 29900 17434 29924 17436
rect 29980 17434 30004 17436
rect 30060 17434 30084 17436
rect 30140 17434 30146 17436
rect 29900 17382 29902 17434
rect 30082 17382 30084 17434
rect 29838 17380 29844 17382
rect 29900 17380 29924 17382
rect 29980 17380 30004 17382
rect 30060 17380 30084 17382
rect 30140 17380 30146 17382
rect 29838 17371 30146 17380
rect 29838 16348 30146 16357
rect 29838 16346 29844 16348
rect 29900 16346 29924 16348
rect 29980 16346 30004 16348
rect 30060 16346 30084 16348
rect 30140 16346 30146 16348
rect 29900 16294 29902 16346
rect 30082 16294 30084 16346
rect 29838 16292 29844 16294
rect 29900 16292 29924 16294
rect 29980 16292 30004 16294
rect 30060 16292 30084 16294
rect 30140 16292 30146 16294
rect 29838 16283 30146 16292
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29196 15162 29224 15370
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 29748 14958 29776 15302
rect 29838 15260 30146 15269
rect 29838 15258 29844 15260
rect 29900 15258 29924 15260
rect 29980 15258 30004 15260
rect 30060 15258 30084 15260
rect 30140 15258 30146 15260
rect 29900 15206 29902 15258
rect 30082 15206 30084 15258
rect 29838 15204 29844 15206
rect 29900 15204 29924 15206
rect 29980 15204 30004 15206
rect 30060 15204 30084 15206
rect 30140 15204 30146 15206
rect 29838 15195 30146 15204
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29748 14278 29776 14894
rect 30208 14346 30236 20470
rect 30852 20058 30880 20742
rect 31220 20602 31248 20742
rect 31208 20596 31260 20602
rect 31208 20538 31260 20544
rect 31312 20482 31340 20946
rect 31404 20602 31432 21286
rect 31484 20868 31536 20874
rect 31484 20810 31536 20816
rect 31392 20596 31444 20602
rect 31392 20538 31444 20544
rect 31312 20454 31432 20482
rect 31496 20466 31524 20810
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 31116 19304 31168 19310
rect 31116 19246 31168 19252
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30576 18358 30604 19110
rect 31128 18970 31156 19246
rect 31116 18964 31168 18970
rect 31116 18906 31168 18912
rect 30932 18896 30984 18902
rect 30932 18838 30984 18844
rect 30564 18352 30616 18358
rect 30564 18294 30616 18300
rect 30840 16584 30892 16590
rect 30840 16526 30892 16532
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30300 15094 30328 16390
rect 30852 16250 30880 16526
rect 30840 16244 30892 16250
rect 30840 16186 30892 16192
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30196 14340 30248 14346
rect 30196 14282 30248 14288
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29276 13728 29328 13734
rect 29276 13670 29328 13676
rect 29288 13326 29316 13670
rect 29748 13326 29776 14214
rect 29838 14172 30146 14181
rect 29838 14170 29844 14172
rect 29900 14170 29924 14172
rect 29980 14170 30004 14172
rect 30060 14170 30084 14172
rect 30140 14170 30146 14172
rect 29900 14118 29902 14170
rect 30082 14118 30084 14170
rect 29838 14116 29844 14118
rect 29900 14116 29924 14118
rect 29980 14116 30004 14118
rect 30060 14116 30084 14118
rect 30140 14116 30146 14118
rect 29838 14107 30146 14116
rect 30208 14074 30236 14282
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29092 13252 29144 13258
rect 29092 13194 29144 13200
rect 29104 12986 29132 13194
rect 29748 12986 29776 13262
rect 29838 13084 30146 13093
rect 29838 13082 29844 13084
rect 29900 13082 29924 13084
rect 29980 13082 30004 13084
rect 30060 13082 30084 13084
rect 30140 13082 30146 13084
rect 29900 13030 29902 13082
rect 30082 13030 30084 13082
rect 29838 13028 29844 13030
rect 29900 13028 29924 13030
rect 29980 13028 30004 13030
rect 30060 13028 30084 13030
rect 30140 13028 30146 13030
rect 29838 13019 30146 13028
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 29552 12164 29604 12170
rect 29552 12106 29604 12112
rect 29092 11688 29144 11694
rect 29092 11630 29144 11636
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 29012 11286 29040 11494
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28552 10266 28580 11086
rect 28816 11008 28868 11014
rect 28816 10950 28868 10956
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 28828 9926 28856 10950
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28828 9654 28856 9862
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28460 7546 28488 8434
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 28552 5914 28580 9454
rect 28724 7744 28776 7750
rect 28724 7686 28776 7692
rect 28736 7546 28764 7686
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28828 7410 28856 9590
rect 29012 9110 29040 10406
rect 29104 10130 29132 11630
rect 29460 11552 29512 11558
rect 29460 11494 29512 11500
rect 29472 11354 29500 11494
rect 29460 11348 29512 11354
rect 29460 11290 29512 11296
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 29380 10674 29408 10950
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29276 10464 29328 10470
rect 29276 10406 29328 10412
rect 29288 10266 29316 10406
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29092 10124 29144 10130
rect 29092 10066 29144 10072
rect 29104 9926 29132 10066
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29000 9104 29052 9110
rect 29000 9046 29052 9052
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 29380 7954 29408 8366
rect 29472 8362 29500 9318
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29368 7948 29420 7954
rect 29368 7890 29420 7896
rect 29472 7750 29500 8298
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 29472 7206 29500 7686
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28828 6322 28856 6598
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 28540 5908 28592 5914
rect 28540 5850 28592 5856
rect 28552 5574 28580 5850
rect 29012 5574 29040 6802
rect 29276 5636 29328 5642
rect 29276 5578 29328 5584
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28080 4548 28132 4554
rect 28080 4490 28132 4496
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 27264 3194 27292 4082
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27356 3369 27384 3878
rect 27342 3360 27398 3369
rect 27342 3295 27398 3304
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27448 2650 27476 4014
rect 27540 3194 27568 4082
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27632 3058 27660 4218
rect 27804 3936 27856 3942
rect 27804 3878 27856 3884
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27816 2961 27844 3878
rect 27802 2952 27858 2961
rect 27802 2887 27858 2896
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 27632 1442 27660 2450
rect 27724 2446 27752 2790
rect 28092 2774 28120 4490
rect 28276 3398 28304 4558
rect 28736 4486 28764 4966
rect 28828 4758 28856 4966
rect 28816 4752 28868 4758
rect 28816 4694 28868 4700
rect 29012 4706 29040 5510
rect 29288 5370 29316 5578
rect 29368 5568 29420 5574
rect 29368 5510 29420 5516
rect 29276 5364 29328 5370
rect 29276 5306 29328 5312
rect 29380 5234 29408 5510
rect 29368 5228 29420 5234
rect 29368 5170 29420 5176
rect 29012 4678 29408 4706
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 28632 4480 28684 4486
rect 28632 4422 28684 4428
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28276 3126 28304 3334
rect 28264 3120 28316 3126
rect 28264 3062 28316 3068
rect 28000 2746 28120 2774
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27448 1414 27660 1442
rect 26804 870 26924 898
rect 26804 762 26832 870
rect 26896 800 26924 870
rect 27448 800 27476 1414
rect 28000 800 28028 2746
rect 28552 800 28580 3402
rect 28644 2650 28672 4422
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 28736 3738 28764 4082
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28828 2310 28856 4082
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 29104 3194 29132 3402
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29196 3058 29224 4490
rect 29380 3398 29408 4678
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29472 3738 29500 4082
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 29564 3505 29592 12106
rect 29656 7546 29684 12786
rect 29838 11996 30146 12005
rect 29838 11994 29844 11996
rect 29900 11994 29924 11996
rect 29980 11994 30004 11996
rect 30060 11994 30084 11996
rect 30140 11994 30146 11996
rect 29900 11942 29902 11994
rect 30082 11942 30084 11994
rect 29838 11940 29844 11942
rect 29900 11940 29924 11942
rect 29980 11940 30004 11942
rect 30060 11940 30084 11942
rect 30140 11940 30146 11942
rect 29838 11931 30146 11940
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29748 10810 29776 10950
rect 29838 10908 30146 10917
rect 29838 10906 29844 10908
rect 29900 10906 29924 10908
rect 29980 10906 30004 10908
rect 30060 10906 30084 10908
rect 30140 10906 30146 10908
rect 29900 10854 29902 10906
rect 30082 10854 30084 10906
rect 29838 10852 29844 10854
rect 29900 10852 29924 10854
rect 29980 10852 30004 10854
rect 30060 10852 30084 10854
rect 30140 10852 30146 10854
rect 29838 10843 30146 10852
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29838 9820 30146 9829
rect 29838 9818 29844 9820
rect 29900 9818 29924 9820
rect 29980 9818 30004 9820
rect 30060 9818 30084 9820
rect 30140 9818 30146 9820
rect 29900 9766 29902 9818
rect 30082 9766 30084 9818
rect 29838 9764 29844 9766
rect 29900 9764 29924 9766
rect 29980 9764 30004 9766
rect 30060 9764 30084 9766
rect 30140 9764 30146 9766
rect 29838 9755 30146 9764
rect 30208 8906 30236 14010
rect 30300 12918 30328 14214
rect 30288 12912 30340 12918
rect 30288 12854 30340 12860
rect 30576 11694 30604 15438
rect 30852 15366 30880 16050
rect 30944 16028 30972 18838
rect 31116 18624 31168 18630
rect 31168 18584 31248 18612
rect 31116 18566 31168 18572
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31036 17338 31064 17546
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 31220 16454 31248 18584
rect 31208 16448 31260 16454
rect 31208 16390 31260 16396
rect 31024 16040 31076 16046
rect 30944 16000 31024 16028
rect 31024 15982 31076 15988
rect 30840 15360 30892 15366
rect 30892 15320 30972 15348
rect 30840 15302 30892 15308
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30852 14074 30880 14350
rect 30944 14074 30972 15320
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30944 13326 30972 14010
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31036 12238 31064 15982
rect 31220 15502 31248 16390
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31300 15428 31352 15434
rect 31300 15370 31352 15376
rect 31312 15162 31340 15370
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31128 13870 31156 14282
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 31208 13864 31260 13870
rect 31208 13806 31260 13812
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 31128 13025 31156 13126
rect 31114 13016 31170 13025
rect 31114 12951 31170 12960
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30576 10606 30604 11018
rect 30668 10810 30696 12038
rect 30932 11688 30984 11694
rect 30932 11630 30984 11636
rect 30944 11354 30972 11630
rect 31036 11626 31064 12174
rect 31128 11898 31156 12951
rect 31220 12714 31248 13806
rect 31404 13734 31432 20454
rect 31484 20460 31536 20466
rect 31484 20402 31536 20408
rect 31496 18698 31524 20402
rect 31588 20330 31616 21422
rect 31668 21412 31720 21418
rect 31668 21354 31720 21360
rect 31680 20466 31708 21354
rect 32968 21350 32996 21422
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31864 20602 31892 20878
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 31852 20596 31904 20602
rect 31852 20538 31904 20544
rect 32140 20534 32168 20742
rect 32128 20528 32180 20534
rect 32128 20470 32180 20476
rect 32968 20466 32996 21286
rect 33428 20806 33456 21422
rect 36912 21412 36964 21418
rect 36912 21354 36964 21360
rect 37648 21412 37700 21418
rect 37648 21354 37700 21360
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 36728 21344 36780 21350
rect 36728 21286 36780 21292
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 33416 20800 33468 20806
rect 33416 20742 33468 20748
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 32956 20460 33008 20466
rect 32956 20402 33008 20408
rect 31576 20324 31628 20330
rect 31576 20266 31628 20272
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 31576 19168 31628 19174
rect 31576 19110 31628 19116
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31588 18902 31616 19110
rect 31576 18896 31628 18902
rect 31576 18838 31628 18844
rect 31956 18766 31984 19110
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 31588 17202 31616 18566
rect 31944 18080 31996 18086
rect 31944 18022 31996 18028
rect 31956 17610 31984 18022
rect 31944 17604 31996 17610
rect 31944 17546 31996 17552
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31956 16794 31984 17546
rect 32048 17338 32076 18702
rect 32140 18086 32168 19654
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32128 18080 32180 18086
rect 32128 18022 32180 18028
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32416 16726 32444 18362
rect 32784 18222 32812 19110
rect 32968 18630 32996 20402
rect 33520 20398 33548 20810
rect 33784 20800 33836 20806
rect 33784 20742 33836 20748
rect 33796 20466 33824 20742
rect 33784 20460 33836 20466
rect 33784 20402 33836 20408
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33876 20392 33928 20398
rect 33876 20334 33928 20340
rect 33244 20058 33272 20334
rect 33600 20324 33652 20330
rect 33600 20266 33652 20272
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33508 19780 33560 19786
rect 33508 19722 33560 19728
rect 33520 19514 33548 19722
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33612 19310 33640 20266
rect 33600 19304 33652 19310
rect 33600 19246 33652 19252
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 33152 18834 33180 19110
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33612 18766 33640 19246
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 32968 18272 32996 18566
rect 33140 18284 33192 18290
rect 32968 18244 33140 18272
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32968 17610 32996 18244
rect 33140 18226 33192 18232
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32956 17604 33008 17610
rect 32956 17546 33008 17552
rect 32876 17338 32904 17546
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 32864 16788 32916 16794
rect 32864 16730 32916 16736
rect 32404 16720 32456 16726
rect 32404 16662 32456 16668
rect 31852 16040 31904 16046
rect 31852 15982 31904 15988
rect 31864 15638 31892 15982
rect 31760 15632 31812 15638
rect 31760 15574 31812 15580
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 31772 14958 31800 15574
rect 31760 14952 31812 14958
rect 31760 14894 31812 14900
rect 31864 14890 31892 15574
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 31944 15360 31996 15366
rect 31944 15302 31996 15308
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 31956 15162 31984 15302
rect 31944 15156 31996 15162
rect 31944 15098 31996 15104
rect 32048 15026 32076 15302
rect 32036 15020 32088 15026
rect 32036 14962 32088 14968
rect 31852 14884 31904 14890
rect 31852 14826 31904 14832
rect 32232 14278 32260 15438
rect 32416 14618 32444 16662
rect 32876 15910 32904 16730
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32876 14958 32904 15846
rect 32968 15570 32996 17546
rect 33428 17542 33456 18158
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 33428 17202 33456 17478
rect 33612 17202 33640 18566
rect 33888 18426 33916 20334
rect 33980 19514 34008 21286
rect 34532 20942 34560 21286
rect 36740 21078 36768 21286
rect 36728 21072 36780 21078
rect 36728 21014 36780 21020
rect 36924 21026 36952 21354
rect 37060 21244 37368 21253
rect 37060 21242 37066 21244
rect 37122 21242 37146 21244
rect 37202 21242 37226 21244
rect 37282 21242 37306 21244
rect 37362 21242 37368 21244
rect 37122 21190 37124 21242
rect 37304 21190 37306 21242
rect 37060 21188 37066 21190
rect 37122 21188 37146 21190
rect 37202 21188 37226 21190
rect 37282 21188 37306 21190
rect 37362 21188 37368 21190
rect 37060 21179 37368 21188
rect 36924 21010 37044 21026
rect 36924 21004 37056 21010
rect 36924 20998 37004 21004
rect 37004 20946 37056 20952
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 34532 20534 34560 20878
rect 34612 20868 34664 20874
rect 34612 20810 34664 20816
rect 34520 20528 34572 20534
rect 34520 20470 34572 20476
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34164 20058 34192 20402
rect 34624 20058 34652 20810
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34716 20466 34744 20742
rect 35268 20602 35296 20878
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 37556 20800 37608 20806
rect 37556 20742 37608 20748
rect 35256 20596 35308 20602
rect 35256 20538 35308 20544
rect 36004 20466 36032 20742
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 35716 20460 35768 20466
rect 35716 20402 35768 20408
rect 35992 20460 36044 20466
rect 35992 20402 36044 20408
rect 35532 20324 35584 20330
rect 35532 20266 35584 20272
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34980 20256 35032 20262
rect 34980 20198 35032 20204
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 34612 20052 34664 20058
rect 34612 19994 34664 20000
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 34348 19310 34376 19654
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34244 18760 34296 18766
rect 34244 18702 34296 18708
rect 33876 18420 33928 18426
rect 33876 18362 33928 18368
rect 33888 18154 33916 18362
rect 34256 18222 34284 18702
rect 34244 18216 34296 18222
rect 34244 18158 34296 18164
rect 33876 18148 33928 18154
rect 33876 18090 33928 18096
rect 33784 18080 33836 18086
rect 33784 18022 33836 18028
rect 33796 17746 33824 18022
rect 34256 17882 34284 18158
rect 34244 17876 34296 17882
rect 34244 17818 34296 17824
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 34428 17740 34480 17746
rect 34428 17682 34480 17688
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33520 15638 33548 16526
rect 34244 16516 34296 16522
rect 34244 16458 34296 16464
rect 34256 16182 34284 16458
rect 34244 16176 34296 16182
rect 34244 16118 34296 16124
rect 33508 15632 33560 15638
rect 33508 15574 33560 15580
rect 32956 15564 33008 15570
rect 32956 15506 33008 15512
rect 33140 15496 33192 15502
rect 33060 15444 33140 15450
rect 33060 15438 33192 15444
rect 33060 15422 33180 15438
rect 33060 15026 33088 15422
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32404 14612 32456 14618
rect 32404 14554 32456 14560
rect 32220 14272 32272 14278
rect 32220 14214 32272 14220
rect 31392 13728 31444 13734
rect 31392 13670 31444 13676
rect 32128 13728 32180 13734
rect 32128 13670 32180 13676
rect 31404 13394 31432 13670
rect 32140 13394 32168 13670
rect 31392 13388 31444 13394
rect 31392 13330 31444 13336
rect 32128 13388 32180 13394
rect 32128 13330 32180 13336
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31312 12918 31340 13194
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31208 12708 31260 12714
rect 31208 12650 31260 12656
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31024 11620 31076 11626
rect 31024 11562 31076 11568
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 30944 11098 30972 11290
rect 31128 11150 31156 11834
rect 31116 11144 31168 11150
rect 30944 11070 31064 11098
rect 31116 11086 31168 11092
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30668 10713 30696 10746
rect 30654 10704 30710 10713
rect 31036 10674 31064 11070
rect 30654 10639 30710 10648
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 30564 10600 30616 10606
rect 30564 10542 30616 10548
rect 30576 9926 30604 10542
rect 30944 10130 30972 10610
rect 31300 10600 31352 10606
rect 31300 10542 31352 10548
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 30564 9920 30616 9926
rect 30564 9862 30616 9868
rect 30196 8900 30248 8906
rect 30196 8842 30248 8848
rect 29838 8732 30146 8741
rect 29838 8730 29844 8732
rect 29900 8730 29924 8732
rect 29980 8730 30004 8732
rect 30060 8730 30084 8732
rect 30140 8730 30146 8732
rect 29900 8678 29902 8730
rect 30082 8678 30084 8730
rect 29838 8676 29844 8678
rect 29900 8676 29924 8678
rect 29980 8676 30004 8678
rect 30060 8676 30084 8678
rect 30140 8676 30146 8678
rect 29838 8667 30146 8676
rect 29838 7644 30146 7653
rect 29838 7642 29844 7644
rect 29900 7642 29924 7644
rect 29980 7642 30004 7644
rect 30060 7642 30084 7644
rect 30140 7642 30146 7644
rect 29900 7590 29902 7642
rect 30082 7590 30084 7642
rect 29838 7588 29844 7590
rect 29900 7588 29924 7590
rect 29980 7588 30004 7590
rect 30060 7588 30084 7590
rect 30140 7588 30146 7590
rect 29838 7579 30146 7588
rect 29644 7540 29696 7546
rect 29644 7482 29696 7488
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29656 5370 29684 5646
rect 29644 5364 29696 5370
rect 29644 5306 29696 5312
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29550 3496 29606 3505
rect 29550 3431 29606 3440
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 29012 2650 29040 2994
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 29104 800 29132 2926
rect 29288 2446 29316 3334
rect 29276 2440 29328 2446
rect 29276 2382 29328 2388
rect 29656 800 29684 4082
rect 29748 4078 29776 7346
rect 30208 7274 30236 8842
rect 30576 8498 30604 9862
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30760 9489 30788 9522
rect 30746 9480 30802 9489
rect 30746 9415 30802 9424
rect 30760 8838 30788 9415
rect 30852 9178 30880 9590
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30932 9172 30984 9178
rect 30932 9114 30984 9120
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30852 8498 30880 9114
rect 30564 8492 30616 8498
rect 30564 8434 30616 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30196 7268 30248 7274
rect 30196 7210 30248 7216
rect 30208 6934 30236 7210
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30392 7002 30420 7142
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30196 6928 30248 6934
rect 30194 6896 30196 6905
rect 30248 6896 30250 6905
rect 30194 6831 30250 6840
rect 29838 6556 30146 6565
rect 29838 6554 29844 6556
rect 29900 6554 29924 6556
rect 29980 6554 30004 6556
rect 30060 6554 30084 6556
rect 30140 6554 30146 6556
rect 29900 6502 29902 6554
rect 30082 6502 30084 6554
rect 29838 6500 29844 6502
rect 29900 6500 29924 6502
rect 29980 6500 30004 6502
rect 30060 6500 30084 6502
rect 30140 6500 30146 6502
rect 29838 6491 30146 6500
rect 30196 6112 30248 6118
rect 30196 6054 30248 6060
rect 30208 5778 30236 6054
rect 30392 5914 30420 6938
rect 30484 6866 30512 7754
rect 30576 7546 30604 8434
rect 30564 7540 30616 7546
rect 30564 7482 30616 7488
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6866 30604 7142
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 29838 5468 30146 5477
rect 29838 5466 29844 5468
rect 29900 5466 29924 5468
rect 29980 5466 30004 5468
rect 30060 5466 30084 5468
rect 30140 5466 30146 5468
rect 29900 5414 29902 5466
rect 30082 5414 30084 5466
rect 29838 5412 29844 5414
rect 29900 5412 29924 5414
rect 29980 5412 30004 5414
rect 30060 5412 30084 5414
rect 30140 5412 30146 5414
rect 29838 5403 30146 5412
rect 30208 5166 30236 5714
rect 30944 5710 30972 9114
rect 31220 9042 31248 10406
rect 31312 9654 31340 10542
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 31208 9036 31260 9042
rect 31208 8978 31260 8984
rect 31312 8922 31340 9590
rect 31404 9178 31432 13330
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31496 12782 31524 13262
rect 32128 13252 32180 13258
rect 32232 13240 32260 14214
rect 32324 13870 32352 14554
rect 32876 14278 32904 14894
rect 32864 14272 32916 14278
rect 32864 14214 32916 14220
rect 32876 13938 32904 14214
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32180 13212 32260 13240
rect 32128 13194 32180 13200
rect 32036 13184 32088 13190
rect 32036 13126 32088 13132
rect 31668 12980 31720 12986
rect 31668 12922 31720 12928
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 31680 12442 31708 12922
rect 32048 12918 32076 13126
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 31668 12436 31720 12442
rect 31668 12378 31720 12384
rect 32036 12096 32088 12102
rect 32140 12084 32168 13194
rect 32324 12986 32352 13806
rect 32692 13530 32720 13806
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32680 13524 32732 13530
rect 32680 13466 32732 13472
rect 32968 13394 32996 13670
rect 33520 13462 33548 15574
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34348 14822 34376 15438
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34336 14408 34388 14414
rect 34336 14350 34388 14356
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33796 13938 33824 14214
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33508 13456 33560 13462
rect 33508 13398 33560 13404
rect 33600 13456 33652 13462
rect 33600 13398 33652 13404
rect 32956 13388 33008 13394
rect 32956 13330 33008 13336
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32404 12640 32456 12646
rect 32404 12582 32456 12588
rect 32088 12056 32168 12084
rect 32036 12038 32088 12044
rect 32048 11082 32076 12038
rect 32416 11626 32444 12582
rect 33324 12164 33376 12170
rect 33324 12106 33376 12112
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32416 11150 32444 11562
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32036 11076 32088 11082
rect 32036 11018 32088 11024
rect 32784 10674 32812 11834
rect 33140 11688 33192 11694
rect 33140 11630 33192 11636
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 33152 10470 33180 11630
rect 33336 11354 33364 12106
rect 33520 11898 33548 13398
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31392 9172 31444 9178
rect 31392 9114 31444 9120
rect 31772 8974 31800 10066
rect 31956 9926 31984 10406
rect 33428 10062 33456 10610
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31944 9920 31996 9926
rect 31944 9862 31996 9868
rect 33232 9920 33284 9926
rect 33232 9862 33284 9868
rect 31864 9586 31892 9862
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 31852 9580 31904 9586
rect 31852 9522 31904 9528
rect 31864 9382 31892 9522
rect 31852 9376 31904 9382
rect 31852 9318 31904 9324
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 31760 8968 31812 8974
rect 31312 8894 31432 8922
rect 31760 8910 31812 8916
rect 31300 8832 31352 8838
rect 31300 8774 31352 8780
rect 31312 8634 31340 8774
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31404 8362 31432 8894
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31392 8356 31444 8362
rect 31392 8298 31444 8304
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 31128 7002 31156 7278
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 31298 6896 31354 6905
rect 31298 6831 31354 6840
rect 31024 6656 31076 6662
rect 31024 6598 31076 6604
rect 31036 6390 31064 6598
rect 31024 6384 31076 6390
rect 31024 6326 31076 6332
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 30932 5704 30984 5710
rect 30932 5646 30984 5652
rect 31128 5370 31156 6258
rect 31312 5370 31340 6831
rect 31392 6248 31444 6254
rect 31392 6190 31444 6196
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 31300 5364 31352 5370
rect 31300 5306 31352 5312
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30196 4548 30248 4554
rect 30300 4536 30328 5306
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 30748 4752 30800 4758
rect 30748 4694 30800 4700
rect 30248 4508 30328 4536
rect 30196 4490 30248 4496
rect 29838 4380 30146 4389
rect 29838 4378 29844 4380
rect 29900 4378 29924 4380
rect 29980 4378 30004 4380
rect 30060 4378 30084 4380
rect 30140 4378 30146 4380
rect 29900 4326 29902 4378
rect 30082 4326 30084 4378
rect 29838 4324 29844 4326
rect 29900 4324 29924 4326
rect 29980 4324 30004 4326
rect 30060 4324 30084 4326
rect 30140 4324 30146 4326
rect 29838 4315 30146 4324
rect 30208 4162 30236 4490
rect 30116 4134 30236 4162
rect 30378 4176 30434 4185
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 30116 3602 30144 4134
rect 30760 4146 30788 4694
rect 31312 4690 31340 5170
rect 31404 5166 31432 6190
rect 31588 5710 31616 7482
rect 31576 5704 31628 5710
rect 31496 5664 31576 5692
rect 31496 5273 31524 5664
rect 31576 5646 31628 5652
rect 31482 5264 31538 5273
rect 31482 5199 31538 5208
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31496 4758 31524 5199
rect 31484 4752 31536 4758
rect 31484 4694 31536 4700
rect 31300 4684 31352 4690
rect 31300 4626 31352 4632
rect 30378 4111 30434 4120
rect 30748 4140 30800 4146
rect 30392 4078 30420 4111
rect 30748 4082 30800 4088
rect 31312 4078 31340 4626
rect 30380 4072 30432 4078
rect 30286 4040 30342 4049
rect 30208 3998 30286 4026
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 29748 2514 29776 3334
rect 29838 3292 30146 3301
rect 29838 3290 29844 3292
rect 29900 3290 29924 3292
rect 29980 3290 30004 3292
rect 30060 3290 30084 3292
rect 30140 3290 30146 3292
rect 29900 3238 29902 3290
rect 30082 3238 30084 3290
rect 29838 3236 29844 3238
rect 29900 3236 29924 3238
rect 29980 3236 30004 3238
rect 30060 3236 30084 3238
rect 30140 3236 30146 3238
rect 29838 3227 30146 3236
rect 30208 3176 30236 3998
rect 30380 4014 30432 4020
rect 30840 4072 30892 4078
rect 30840 4014 30892 4020
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 30286 3975 30342 3984
rect 30852 3194 30880 4014
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 30944 3738 30972 3878
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 30116 3148 30236 3176
rect 30840 3188 30892 3194
rect 30116 2514 30144 3148
rect 30840 3130 30892 3136
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 29838 2204 30146 2213
rect 29838 2202 29844 2204
rect 29900 2202 29924 2204
rect 29980 2202 30004 2204
rect 30060 2202 30084 2204
rect 30140 2202 30146 2204
rect 29900 2150 29902 2202
rect 30082 2150 30084 2202
rect 29838 2148 29844 2150
rect 29900 2148 29924 2150
rect 29980 2148 30004 2150
rect 30060 2148 30084 2150
rect 30140 2148 30146 2150
rect 29838 2139 30146 2148
rect 30208 800 30236 2926
rect 31128 2514 31156 3334
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 30748 2372 30800 2378
rect 30748 2314 30800 2320
rect 30760 800 30788 2314
rect 31312 800 31340 3470
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 31404 2650 31432 3334
rect 31680 3058 31708 8774
rect 31772 7954 31800 8910
rect 32416 8430 32444 9318
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31864 7818 31892 8366
rect 32128 8356 32180 8362
rect 32128 8298 32180 8304
rect 31852 7812 31904 7818
rect 31852 7754 31904 7760
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 31772 5710 31800 6598
rect 32140 5846 32168 8298
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32232 6390 32260 7890
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32324 7274 32352 7686
rect 32416 7546 32444 8366
rect 32508 7954 32536 9590
rect 33244 9586 33272 9862
rect 33520 9722 33548 9998
rect 33508 9716 33560 9722
rect 33508 9658 33560 9664
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 32496 7948 32548 7954
rect 32496 7890 32548 7896
rect 32680 7948 32732 7954
rect 32680 7890 32732 7896
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32312 7268 32364 7274
rect 32312 7210 32364 7216
rect 32508 7206 32536 7890
rect 32692 7274 32720 7890
rect 32876 7886 32904 8910
rect 33428 8634 33456 8910
rect 33612 8820 33640 13398
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33796 10742 33824 11494
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33888 10674 33916 11494
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 33692 10600 33744 10606
rect 33692 10542 33744 10548
rect 33704 9722 33732 10542
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33784 8832 33836 8838
rect 33612 8792 33784 8820
rect 33784 8774 33836 8780
rect 33416 8628 33468 8634
rect 33416 8570 33468 8576
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33428 8090 33456 8434
rect 33416 8084 33468 8090
rect 33416 8026 33468 8032
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 33416 7336 33468 7342
rect 33416 7278 33468 7284
rect 32680 7268 32732 7274
rect 32680 7210 32732 7216
rect 33428 7206 33456 7278
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 32508 6798 32536 7142
rect 33428 6882 33456 7142
rect 33336 6854 33456 6882
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32220 6384 32272 6390
rect 32220 6326 32272 6332
rect 33232 6316 33284 6322
rect 33232 6258 33284 6264
rect 32772 6112 32824 6118
rect 32772 6054 32824 6060
rect 32128 5840 32180 5846
rect 32128 5782 32180 5788
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 32140 5370 32168 5782
rect 32784 5710 32812 6054
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32864 5568 32916 5574
rect 32864 5510 32916 5516
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 32140 5234 32168 5306
rect 32588 5296 32640 5302
rect 32588 5238 32640 5244
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32404 5160 32456 5166
rect 32404 5102 32456 5108
rect 32324 5001 32352 5102
rect 32310 4992 32366 5001
rect 32310 4927 32366 4936
rect 32036 4548 32088 4554
rect 32036 4490 32088 4496
rect 31944 4480 31996 4486
rect 31944 4422 31996 4428
rect 31956 4078 31984 4422
rect 31760 4072 31812 4078
rect 31760 4014 31812 4020
rect 31944 4072 31996 4078
rect 31944 4014 31996 4020
rect 31772 3670 31800 4014
rect 31760 3664 31812 3670
rect 31760 3606 31812 3612
rect 31772 3194 31800 3606
rect 32048 3602 32076 4490
rect 32416 4128 32444 5102
rect 32600 4758 32628 5238
rect 32588 4752 32640 4758
rect 32588 4694 32640 4700
rect 32588 4480 32640 4486
rect 32588 4422 32640 4428
rect 32600 4282 32628 4422
rect 32692 4282 32720 5510
rect 32876 5234 32904 5510
rect 33244 5234 33272 6258
rect 33336 5778 33364 6854
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 33416 6724 33468 6730
rect 33416 6666 33468 6672
rect 33428 5914 33456 6666
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 33520 5846 33548 6598
rect 33612 6186 33640 6734
rect 33692 6724 33744 6730
rect 33692 6666 33744 6672
rect 33600 6180 33652 6186
rect 33600 6122 33652 6128
rect 33508 5840 33560 5846
rect 33508 5782 33560 5788
rect 33324 5772 33376 5778
rect 33324 5714 33376 5720
rect 33508 5704 33560 5710
rect 33508 5646 33560 5652
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 33520 5098 33548 5646
rect 33600 5568 33652 5574
rect 33600 5510 33652 5516
rect 33612 5234 33640 5510
rect 33600 5228 33652 5234
rect 33600 5170 33652 5176
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 33600 5092 33652 5098
rect 33600 5034 33652 5040
rect 32770 4992 32826 5001
rect 32770 4927 32826 4936
rect 32784 4554 32812 4927
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 32772 4548 32824 4554
rect 32772 4490 32824 4496
rect 32588 4276 32640 4282
rect 32588 4218 32640 4224
rect 32680 4276 32732 4282
rect 32680 4218 32732 4224
rect 32876 4146 32904 4558
rect 33230 4176 33286 4185
rect 32496 4140 32548 4146
rect 32416 4100 32496 4128
rect 32496 4082 32548 4088
rect 32864 4140 32916 4146
rect 33230 4111 33232 4120
rect 32864 4082 32916 4088
rect 33284 4111 33286 4120
rect 33232 4082 33284 4088
rect 32508 3602 32536 4082
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 32496 3596 32548 3602
rect 33520 3584 33548 4558
rect 33612 4078 33640 5034
rect 33600 4072 33652 4078
rect 33600 4014 33652 4020
rect 33600 3596 33652 3602
rect 33520 3556 33600 3584
rect 32496 3538 32548 3544
rect 33600 3538 33652 3544
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31760 3188 31812 3194
rect 31760 3130 31812 3136
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 31772 2446 31800 2790
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 31956 1850 31984 3470
rect 33232 3460 33284 3466
rect 33232 3402 33284 3408
rect 32036 2916 32088 2922
rect 32036 2858 32088 2864
rect 32048 2446 32076 2858
rect 33244 2446 33272 3402
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 33520 3194 33548 3334
rect 33508 3188 33560 3194
rect 33508 3130 33560 3136
rect 33508 3052 33560 3058
rect 33612 3040 33640 3538
rect 33560 3012 33640 3040
rect 33508 2994 33560 3000
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 31864 1822 31984 1850
rect 31864 800 31892 1822
rect 32416 800 32444 2314
rect 33048 1420 33100 1426
rect 33048 1362 33100 1368
rect 33060 898 33088 1362
rect 32968 870 33088 898
rect 32968 800 32996 870
rect 33520 800 33548 2858
rect 33704 2774 33732 6666
rect 33796 5098 33824 8774
rect 33876 5840 33928 5846
rect 33876 5782 33928 5788
rect 33888 5234 33916 5782
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 33784 4684 33836 4690
rect 33784 4626 33836 4632
rect 33796 4146 33824 4626
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33888 4078 33916 4558
rect 33980 4146 34008 14010
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 34164 13258 34192 13874
rect 34244 13796 34296 13802
rect 34244 13738 34296 13744
rect 34256 13394 34284 13738
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34152 13252 34204 13258
rect 34152 13194 34204 13200
rect 34348 12986 34376 14350
rect 34440 13462 34468 17682
rect 34716 17610 34744 20198
rect 34992 19378 35020 20198
rect 35544 19854 35572 20266
rect 35728 19922 35756 20402
rect 37060 20156 37368 20165
rect 37060 20154 37066 20156
rect 37122 20154 37146 20156
rect 37202 20154 37226 20156
rect 37282 20154 37306 20156
rect 37362 20154 37368 20156
rect 37122 20102 37124 20154
rect 37304 20102 37306 20154
rect 37060 20100 37066 20102
rect 37122 20100 37146 20102
rect 37202 20100 37226 20102
rect 37282 20100 37306 20102
rect 37362 20100 37368 20102
rect 37060 20091 37368 20100
rect 35716 19916 35768 19922
rect 35716 19858 35768 19864
rect 35256 19848 35308 19854
rect 35256 19790 35308 19796
rect 35532 19848 35584 19854
rect 35532 19790 35584 19796
rect 35268 19514 35296 19790
rect 37280 19780 37332 19786
rect 37280 19722 37332 19728
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35256 19508 35308 19514
rect 35256 19450 35308 19456
rect 34980 19372 35032 19378
rect 34980 19314 35032 19320
rect 34888 19168 34940 19174
rect 34888 19110 34940 19116
rect 34900 18834 34928 19110
rect 34888 18828 34940 18834
rect 34888 18770 34940 18776
rect 35164 18828 35216 18834
rect 35164 18770 35216 18776
rect 34704 17604 34756 17610
rect 34704 17546 34756 17552
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34532 16998 34560 17478
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34532 16794 34560 16934
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 34704 16448 34756 16454
rect 34704 16390 34756 16396
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34532 15570 34560 16186
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34716 15162 34744 16390
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 15156 34756 15162
rect 34704 15098 34756 15104
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 34428 13456 34480 13462
rect 34428 13398 34480 13404
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 34336 12980 34388 12986
rect 34336 12922 34388 12928
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34152 11076 34204 11082
rect 34152 11018 34204 11024
rect 34164 9586 34192 11018
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 34244 9376 34296 9382
rect 34244 9318 34296 9324
rect 34256 8838 34284 9318
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34256 8498 34284 8774
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34244 7540 34296 7546
rect 34348 7528 34376 12786
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 34532 12442 34560 12718
rect 34624 12646 34652 13262
rect 34716 12918 34744 14214
rect 34808 13870 34836 15370
rect 34900 15366 34928 18770
rect 35176 15570 35204 18770
rect 35360 18358 35388 19654
rect 37292 19514 37320 19722
rect 37280 19508 37332 19514
rect 37280 19450 37332 19456
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 36924 18970 36952 19110
rect 37060 19068 37368 19077
rect 37060 19066 37066 19068
rect 37122 19066 37146 19068
rect 37202 19066 37226 19068
rect 37282 19066 37306 19068
rect 37362 19066 37368 19068
rect 37122 19014 37124 19066
rect 37304 19014 37306 19066
rect 37060 19012 37066 19014
rect 37122 19012 37146 19014
rect 37202 19012 37226 19014
rect 37282 19012 37306 19014
rect 37362 19012 37368 19014
rect 37060 19003 37368 19012
rect 36912 18964 36964 18970
rect 36912 18906 36964 18912
rect 35900 18760 35952 18766
rect 35900 18702 35952 18708
rect 36820 18760 36872 18766
rect 36820 18702 36872 18708
rect 35532 18624 35584 18630
rect 35532 18566 35584 18572
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 35360 16998 35388 18294
rect 35544 18290 35572 18566
rect 35532 18284 35584 18290
rect 35532 18226 35584 18232
rect 35440 17536 35492 17542
rect 35440 17478 35492 17484
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35256 16584 35308 16590
rect 35256 16526 35308 16532
rect 35268 16250 35296 16526
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35360 16114 35388 16934
rect 35452 16697 35480 17478
rect 35438 16688 35494 16697
rect 35438 16623 35494 16632
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 35440 16448 35492 16454
rect 35440 16390 35492 16396
rect 35452 16250 35480 16390
rect 35440 16244 35492 16250
rect 35440 16186 35492 16192
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 35164 15564 35216 15570
rect 35164 15506 35216 15512
rect 34888 15360 34940 15366
rect 34888 15302 34940 15308
rect 34980 15360 35032 15366
rect 34980 15302 35032 15308
rect 35072 15360 35124 15366
rect 35072 15302 35124 15308
rect 34900 14890 34928 15302
rect 34992 15162 35020 15302
rect 34980 15156 35032 15162
rect 34980 15098 35032 15104
rect 35084 14958 35112 15302
rect 35072 14952 35124 14958
rect 35072 14894 35124 14900
rect 34888 14884 34940 14890
rect 34888 14826 34940 14832
rect 34796 13864 34848 13870
rect 34796 13806 34848 13812
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34520 12436 34572 12442
rect 34624 12434 34652 12582
rect 34624 12406 34744 12434
rect 34520 12378 34572 12384
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 34440 10538 34468 11630
rect 34532 11218 34560 12378
rect 34716 12306 34744 12406
rect 34704 12300 34756 12306
rect 34704 12242 34756 12248
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34532 10674 34560 11154
rect 34612 11008 34664 11014
rect 34808 10996 34836 13262
rect 34900 11082 34928 14826
rect 34980 14408 35032 14414
rect 34980 14350 35032 14356
rect 34992 13530 35020 14350
rect 34980 13524 35032 13530
rect 34980 13466 35032 13472
rect 35084 13190 35112 14894
rect 35176 13326 35204 15506
rect 35532 15360 35584 15366
rect 35532 15302 35584 15308
rect 35544 15094 35572 15302
rect 35532 15088 35584 15094
rect 35532 15030 35584 15036
rect 35636 14958 35664 16594
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35256 13728 35308 13734
rect 35256 13670 35308 13676
rect 35164 13320 35216 13326
rect 35164 13262 35216 13268
rect 35072 13184 35124 13190
rect 35072 13126 35124 13132
rect 35164 13184 35216 13190
rect 35164 13126 35216 13132
rect 35084 12850 35112 13126
rect 35072 12844 35124 12850
rect 35072 12786 35124 12792
rect 35176 12442 35204 13126
rect 35268 12986 35296 13670
rect 35360 13530 35388 13806
rect 35348 13524 35400 13530
rect 35348 13466 35400 13472
rect 35808 13456 35860 13462
rect 35806 13424 35808 13433
rect 35860 13424 35862 13433
rect 35636 13382 35806 13410
rect 35256 12980 35308 12986
rect 35256 12922 35308 12928
rect 35532 12776 35584 12782
rect 35530 12744 35532 12753
rect 35584 12744 35586 12753
rect 35530 12679 35586 12688
rect 35164 12436 35216 12442
rect 35164 12378 35216 12384
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34888 11076 34940 11082
rect 34888 11018 34940 11024
rect 34664 10968 34836 10996
rect 34612 10950 34664 10956
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34624 10606 34652 10950
rect 34612 10600 34664 10606
rect 34612 10542 34664 10548
rect 34428 10532 34480 10538
rect 34428 10474 34480 10480
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34532 7546 34560 8434
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 34296 7500 34376 7528
rect 34520 7540 34572 7546
rect 34244 7482 34296 7488
rect 34520 7482 34572 7488
rect 34900 7410 34928 7686
rect 35268 7546 35296 7686
rect 35256 7540 35308 7546
rect 35256 7482 35308 7488
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 34980 6928 35032 6934
rect 34978 6896 34980 6905
rect 35032 6896 35034 6905
rect 34978 6831 35034 6840
rect 35256 6724 35308 6730
rect 35256 6666 35308 6672
rect 35268 6390 35296 6666
rect 35256 6384 35308 6390
rect 35256 6326 35308 6332
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34440 5166 34468 6190
rect 34888 5296 34940 5302
rect 34886 5264 34888 5273
rect 34940 5264 34942 5273
rect 34886 5199 34942 5208
rect 34428 5160 34480 5166
rect 34428 5102 34480 5108
rect 34612 5024 34664 5030
rect 34612 4966 34664 4972
rect 34152 4548 34204 4554
rect 34152 4490 34204 4496
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 34060 3936 34112 3942
rect 34060 3878 34112 3884
rect 33704 2746 33824 2774
rect 33796 2650 33824 2746
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 34072 2446 34100 3878
rect 34164 2854 34192 4490
rect 34520 3936 34572 3942
rect 34520 3878 34572 3884
rect 34532 3534 34560 3878
rect 34520 3528 34572 3534
rect 34520 3470 34572 3476
rect 34624 3194 34652 4966
rect 35162 4584 35218 4593
rect 35162 4519 35164 4528
rect 35216 4519 35218 4528
rect 35164 4490 35216 4496
rect 35360 4078 35388 11698
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 35452 6390 35480 6598
rect 35544 6390 35572 12679
rect 35636 7410 35664 13382
rect 35806 13359 35862 13368
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35820 12850 35848 13262
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35716 12096 35768 12102
rect 35716 12038 35768 12044
rect 35728 10742 35756 12038
rect 35808 11076 35860 11082
rect 35808 11018 35860 11024
rect 35716 10736 35768 10742
rect 35716 10678 35768 10684
rect 35820 10266 35848 11018
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35912 9654 35940 18702
rect 36832 18426 36860 18702
rect 37568 18630 37596 20742
rect 37660 20602 37688 21354
rect 38016 21344 38068 21350
rect 38016 21286 38068 21292
rect 38028 21146 38056 21286
rect 38016 21140 38068 21146
rect 38016 21082 38068 21088
rect 38108 20800 38160 20806
rect 38108 20742 38160 20748
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 37924 20596 37976 20602
rect 37924 20538 37976 20544
rect 37740 18760 37792 18766
rect 37740 18702 37792 18708
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 36820 18420 36872 18426
rect 36820 18362 36872 18368
rect 37568 18086 37596 18566
rect 35992 18080 36044 18086
rect 35992 18022 36044 18028
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 36004 17814 36032 18022
rect 37060 17980 37368 17989
rect 37060 17978 37066 17980
rect 37122 17978 37146 17980
rect 37202 17978 37226 17980
rect 37282 17978 37306 17980
rect 37362 17978 37368 17980
rect 37122 17926 37124 17978
rect 37304 17926 37306 17978
rect 37060 17924 37066 17926
rect 37122 17924 37146 17926
rect 37202 17924 37226 17926
rect 37282 17924 37306 17926
rect 37362 17924 37368 17926
rect 37060 17915 37368 17924
rect 35992 17808 36044 17814
rect 35992 17750 36044 17756
rect 36728 17604 36780 17610
rect 36728 17546 36780 17552
rect 36452 16448 36504 16454
rect 36452 16390 36504 16396
rect 36464 16250 36492 16390
rect 36452 16244 36504 16250
rect 36452 16186 36504 16192
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 36556 14822 36584 15302
rect 36740 15162 36768 17546
rect 37060 16892 37368 16901
rect 37060 16890 37066 16892
rect 37122 16890 37146 16892
rect 37202 16890 37226 16892
rect 37282 16890 37306 16892
rect 37362 16890 37368 16892
rect 37122 16838 37124 16890
rect 37304 16838 37306 16890
rect 37060 16836 37066 16838
rect 37122 16836 37146 16838
rect 37202 16836 37226 16838
rect 37282 16836 37306 16838
rect 37362 16836 37368 16838
rect 37060 16827 37368 16836
rect 36820 16584 36872 16590
rect 36820 16526 36872 16532
rect 36832 15706 36860 16526
rect 36912 16448 36964 16454
rect 36912 16390 36964 16396
rect 36820 15700 36872 15706
rect 36820 15642 36872 15648
rect 36924 15570 36952 16390
rect 37060 15804 37368 15813
rect 37060 15802 37066 15804
rect 37122 15802 37146 15804
rect 37202 15802 37226 15804
rect 37282 15802 37306 15804
rect 37362 15802 37368 15804
rect 37122 15750 37124 15802
rect 37304 15750 37306 15802
rect 37060 15748 37066 15750
rect 37122 15748 37146 15750
rect 37202 15748 37226 15750
rect 37282 15748 37306 15750
rect 37362 15748 37368 15750
rect 37060 15739 37368 15748
rect 36912 15564 36964 15570
rect 36912 15506 36964 15512
rect 37464 15564 37516 15570
rect 37464 15506 37516 15512
rect 36728 15156 36780 15162
rect 36728 15098 36780 15104
rect 37476 15026 37504 15506
rect 37568 15366 37596 18022
rect 37752 17746 37780 18702
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 37844 18426 37872 18566
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37936 17814 37964 20538
rect 38120 19310 38148 20742
rect 38396 20466 38424 21490
rect 38660 21480 38712 21486
rect 38660 21422 38712 21428
rect 39856 21480 39908 21486
rect 39856 21422 39908 21428
rect 43260 21480 43312 21486
rect 43260 21422 43312 21428
rect 43996 21480 44048 21486
rect 43996 21422 44048 21428
rect 44088 21480 44140 21486
rect 44088 21422 44140 21428
rect 46112 21480 46164 21486
rect 46112 21422 46164 21428
rect 48228 21480 48280 21486
rect 48228 21422 48280 21428
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 53380 21480 53432 21486
rect 53380 21422 53432 21428
rect 56600 21480 56652 21486
rect 56600 21422 56652 21428
rect 38476 20800 38528 20806
rect 38476 20742 38528 20748
rect 38568 20800 38620 20806
rect 38568 20742 38620 20748
rect 38488 20602 38516 20742
rect 38476 20596 38528 20602
rect 38476 20538 38528 20544
rect 38384 20460 38436 20466
rect 38384 20402 38436 20408
rect 38580 19310 38608 20742
rect 38672 20398 38700 21422
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 39224 21010 39252 21286
rect 39868 21146 39896 21422
rect 40040 21344 40092 21350
rect 40040 21286 40092 21292
rect 42708 21344 42760 21350
rect 42708 21286 42760 21292
rect 39856 21140 39908 21146
rect 39856 21082 39908 21088
rect 39212 21004 39264 21010
rect 39212 20946 39264 20952
rect 39028 20800 39080 20806
rect 39028 20742 39080 20748
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38856 20398 38884 20538
rect 38660 20392 38712 20398
rect 38660 20334 38712 20340
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38672 20058 38700 20334
rect 38844 20256 38896 20262
rect 38844 20198 38896 20204
rect 38660 20052 38712 20058
rect 38660 19994 38712 20000
rect 38752 19780 38804 19786
rect 38752 19722 38804 19728
rect 38764 19514 38792 19722
rect 38752 19508 38804 19514
rect 38752 19450 38804 19456
rect 38108 19304 38160 19310
rect 38108 19246 38160 19252
rect 38568 19304 38620 19310
rect 38568 19246 38620 19252
rect 38660 19304 38712 19310
rect 38660 19246 38712 19252
rect 38016 19168 38068 19174
rect 38016 19110 38068 19116
rect 38028 18834 38056 19110
rect 38016 18828 38068 18834
rect 38016 18770 38068 18776
rect 38672 18426 38700 19246
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38672 17882 38700 18362
rect 38752 18216 38804 18222
rect 38752 18158 38804 18164
rect 38660 17876 38712 17882
rect 38660 17818 38712 17824
rect 37924 17808 37976 17814
rect 37924 17750 37976 17756
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37648 17672 37700 17678
rect 37648 17614 37700 17620
rect 37660 15910 37688 17614
rect 37752 17338 37780 17682
rect 37740 17332 37792 17338
rect 37740 17274 37792 17280
rect 37936 16810 37964 17750
rect 38476 17672 38528 17678
rect 38476 17614 38528 17620
rect 37752 16782 37964 16810
rect 38292 16788 38344 16794
rect 37648 15904 37700 15910
rect 37648 15846 37700 15852
rect 37556 15360 37608 15366
rect 37556 15302 37608 15308
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 36452 13728 36504 13734
rect 36452 13670 36504 13676
rect 36464 12918 36492 13670
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36176 12232 36228 12238
rect 36176 12174 36228 12180
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36188 11218 36216 12174
rect 36280 11898 36308 12174
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36268 11892 36320 11898
rect 36268 11834 36320 11840
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 35900 9648 35952 9654
rect 35900 9590 35952 9596
rect 36084 9512 36136 9518
rect 36084 9454 36136 9460
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35912 8634 35940 9318
rect 36096 8838 36124 9454
rect 36084 8832 36136 8838
rect 36084 8774 36136 8780
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 36004 7954 36032 8434
rect 36084 8288 36136 8294
rect 36084 8230 36136 8236
rect 35716 7948 35768 7954
rect 35716 7890 35768 7896
rect 35992 7948 36044 7954
rect 35992 7890 36044 7896
rect 35728 7449 35756 7890
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35714 7440 35770 7449
rect 35624 7404 35676 7410
rect 35714 7375 35770 7384
rect 35624 7346 35676 7352
rect 35636 7206 35664 7346
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35728 6934 35756 7375
rect 35716 6928 35768 6934
rect 35716 6870 35768 6876
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 35440 6384 35492 6390
rect 35440 6326 35492 6332
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35636 5846 35664 6802
rect 35624 5840 35676 5846
rect 35624 5782 35676 5788
rect 35636 4690 35664 5782
rect 35820 5234 35848 7482
rect 36096 7342 36124 8230
rect 35900 7336 35952 7342
rect 35900 7278 35952 7284
rect 36084 7336 36136 7342
rect 36084 7278 36136 7284
rect 35912 6934 35940 7278
rect 35900 6928 35952 6934
rect 35900 6870 35952 6876
rect 35992 6792 36044 6798
rect 35992 6734 36044 6740
rect 36004 5370 36032 6734
rect 36084 6656 36136 6662
rect 36084 6598 36136 6604
rect 36096 5370 36124 6598
rect 36188 6254 36216 11154
rect 36360 11008 36412 11014
rect 36360 10950 36412 10956
rect 36372 10130 36400 10950
rect 36360 10124 36412 10130
rect 36360 10066 36412 10072
rect 36464 9178 36492 12038
rect 36556 11694 36584 14758
rect 37060 14716 37368 14725
rect 37060 14714 37066 14716
rect 37122 14714 37146 14716
rect 37202 14714 37226 14716
rect 37282 14714 37306 14716
rect 37362 14714 37368 14716
rect 37122 14662 37124 14714
rect 37304 14662 37306 14714
rect 37060 14660 37066 14662
rect 37122 14660 37146 14662
rect 37202 14660 37226 14662
rect 37282 14660 37306 14662
rect 37362 14660 37368 14662
rect 37060 14651 37368 14660
rect 37464 14272 37516 14278
rect 37464 14214 37516 14220
rect 37476 14074 37504 14214
rect 37464 14068 37516 14074
rect 37752 14056 37780 16782
rect 38292 16730 38344 16736
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37844 16250 37872 16594
rect 37924 16584 37976 16590
rect 37924 16526 37976 16532
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37936 15706 37964 16526
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 37832 14340 37884 14346
rect 37832 14282 37884 14288
rect 37464 14010 37516 14016
rect 37660 14028 37780 14056
rect 37060 13628 37368 13637
rect 37060 13626 37066 13628
rect 37122 13626 37146 13628
rect 37202 13626 37226 13628
rect 37282 13626 37306 13628
rect 37362 13626 37368 13628
rect 37122 13574 37124 13626
rect 37304 13574 37306 13626
rect 37060 13572 37066 13574
rect 37122 13572 37146 13574
rect 37202 13572 37226 13574
rect 37282 13572 37306 13574
rect 37362 13572 37368 13574
rect 37060 13563 37368 13572
rect 36820 13252 36872 13258
rect 36820 13194 36872 13200
rect 36728 12708 36780 12714
rect 36728 12650 36780 12656
rect 36740 12434 36768 12650
rect 36832 12442 36860 13194
rect 37556 12912 37608 12918
rect 37556 12854 37608 12860
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37060 12540 37368 12549
rect 37060 12538 37066 12540
rect 37122 12538 37146 12540
rect 37202 12538 37226 12540
rect 37282 12538 37306 12540
rect 37362 12538 37368 12540
rect 37122 12486 37124 12538
rect 37304 12486 37306 12538
rect 37060 12484 37066 12486
rect 37122 12484 37146 12486
rect 37202 12484 37226 12486
rect 37282 12484 37306 12486
rect 37362 12484 37368 12486
rect 37060 12475 37368 12484
rect 36648 12406 36768 12434
rect 36820 12436 36872 12442
rect 36648 12102 36676 12406
rect 36820 12378 36872 12384
rect 37476 12306 37504 12582
rect 37568 12374 37596 12854
rect 37660 12646 37688 14028
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37752 12918 37780 13874
rect 37844 13870 37872 14282
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 37844 12918 37872 13806
rect 38028 12918 38056 15098
rect 38200 14952 38252 14958
rect 38200 14894 38252 14900
rect 38212 14618 38240 14894
rect 38200 14612 38252 14618
rect 38200 14554 38252 14560
rect 38108 13796 38160 13802
rect 38108 13738 38160 13744
rect 38120 13462 38148 13738
rect 38108 13456 38160 13462
rect 38108 13398 38160 13404
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 37832 12912 37884 12918
rect 37832 12854 37884 12860
rect 38016 12912 38068 12918
rect 38016 12854 38068 12860
rect 37740 12776 37792 12782
rect 37740 12718 37792 12724
rect 37648 12640 37700 12646
rect 37648 12582 37700 12588
rect 37556 12368 37608 12374
rect 37556 12310 37608 12316
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36740 11830 36768 12174
rect 36728 11824 36780 11830
rect 37568 11778 37596 12310
rect 37660 11898 37688 12582
rect 37752 12442 37780 12718
rect 37740 12436 37792 12442
rect 37740 12378 37792 12384
rect 38028 11898 38056 12854
rect 38120 12442 38148 13398
rect 38212 13190 38240 14554
rect 38304 13734 38332 16730
rect 38488 16658 38516 17614
rect 38476 16652 38528 16658
rect 38476 16594 38528 16600
rect 38568 16448 38620 16454
rect 38568 16390 38620 16396
rect 38580 16250 38608 16390
rect 38568 16244 38620 16250
rect 38568 16186 38620 16192
rect 38764 15994 38792 18158
rect 38856 17338 38884 20198
rect 39040 20058 39068 20742
rect 39028 20052 39080 20058
rect 39028 19994 39080 20000
rect 39224 19718 39252 20946
rect 39764 20800 39816 20806
rect 39764 20742 39816 20748
rect 39776 20398 39804 20742
rect 39868 20466 39896 21082
rect 39948 20868 40000 20874
rect 39948 20810 40000 20816
rect 39960 20602 39988 20810
rect 40052 20602 40080 21286
rect 41880 20936 41932 20942
rect 41880 20878 41932 20884
rect 42432 20936 42484 20942
rect 42432 20878 42484 20884
rect 41892 20602 41920 20878
rect 39948 20596 40000 20602
rect 39948 20538 40000 20544
rect 40040 20596 40092 20602
rect 40040 20538 40092 20544
rect 41880 20596 41932 20602
rect 41880 20538 41932 20544
rect 39856 20460 39908 20466
rect 39856 20402 39908 20408
rect 42444 20398 42472 20878
rect 42720 20534 42748 21286
rect 42708 20528 42760 20534
rect 42708 20470 42760 20476
rect 43076 20528 43128 20534
rect 43076 20470 43128 20476
rect 39764 20392 39816 20398
rect 39764 20334 39816 20340
rect 40040 20392 40092 20398
rect 40040 20334 40092 20340
rect 42432 20392 42484 20398
rect 42432 20334 42484 20340
rect 39580 20256 39632 20262
rect 39580 20198 39632 20204
rect 39592 19922 39620 20198
rect 39580 19916 39632 19922
rect 39580 19858 39632 19864
rect 39672 19848 39724 19854
rect 40052 19825 40080 20334
rect 40500 19916 40552 19922
rect 40500 19858 40552 19864
rect 39672 19790 39724 19796
rect 40038 19816 40094 19825
rect 39212 19712 39264 19718
rect 39212 19654 39264 19660
rect 39684 19514 39712 19790
rect 40038 19751 40094 19760
rect 39672 19508 39724 19514
rect 39672 19450 39724 19456
rect 39684 18970 39712 19450
rect 40052 19378 40080 19751
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 39672 18964 39724 18970
rect 39672 18906 39724 18912
rect 39212 18624 39264 18630
rect 39212 18566 39264 18572
rect 39580 18624 39632 18630
rect 39580 18566 39632 18572
rect 39224 18426 39252 18566
rect 39212 18420 39264 18426
rect 39212 18362 39264 18368
rect 39592 18222 39620 18566
rect 39580 18216 39632 18222
rect 39580 18158 39632 18164
rect 39580 18080 39632 18086
rect 39580 18022 39632 18028
rect 39304 17536 39356 17542
rect 39304 17478 39356 17484
rect 39316 17338 39344 17478
rect 38844 17332 38896 17338
rect 38844 17274 38896 17280
rect 39304 17332 39356 17338
rect 39304 17274 39356 17280
rect 39592 17270 39620 18022
rect 39580 17264 39632 17270
rect 39580 17206 39632 17212
rect 38844 16992 38896 16998
rect 38844 16934 38896 16940
rect 39304 16992 39356 16998
rect 39856 16992 39908 16998
rect 39356 16952 39528 16980
rect 39304 16934 39356 16940
rect 38856 16590 38884 16934
rect 38844 16584 38896 16590
rect 38844 16526 38896 16532
rect 38856 16114 38884 16526
rect 38844 16108 38896 16114
rect 38844 16050 38896 16056
rect 38672 15966 38792 15994
rect 38672 15638 38700 15966
rect 38752 15904 38804 15910
rect 38752 15846 38804 15852
rect 38764 15706 38792 15846
rect 38856 15706 38884 16050
rect 38752 15700 38804 15706
rect 38752 15642 38804 15648
rect 38844 15700 38896 15706
rect 38844 15642 38896 15648
rect 38660 15632 38712 15638
rect 38660 15574 38712 15580
rect 38660 15360 38712 15366
rect 38660 15302 38712 15308
rect 38568 14408 38620 14414
rect 38568 14350 38620 14356
rect 38292 13728 38344 13734
rect 38292 13670 38344 13676
rect 38292 13524 38344 13530
rect 38292 13466 38344 13472
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38108 12436 38160 12442
rect 38108 12378 38160 12384
rect 38120 12170 38148 12378
rect 38304 12306 38332 13466
rect 38476 13388 38528 13394
rect 38476 13330 38528 13336
rect 38488 12646 38516 13330
rect 38580 13190 38608 14350
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38580 12986 38608 13126
rect 38568 12980 38620 12986
rect 38568 12922 38620 12928
rect 38476 12640 38528 12646
rect 38476 12582 38528 12588
rect 38292 12300 38344 12306
rect 38292 12242 38344 12248
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 37648 11892 37700 11898
rect 37648 11834 37700 11840
rect 38016 11892 38068 11898
rect 38016 11834 38068 11840
rect 36728 11766 36780 11772
rect 37476 11750 37596 11778
rect 37476 11694 37504 11750
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 37464 11688 37516 11694
rect 37464 11630 37516 11636
rect 37648 11688 37700 11694
rect 37648 11630 37700 11636
rect 37060 11452 37368 11461
rect 37060 11450 37066 11452
rect 37122 11450 37146 11452
rect 37202 11450 37226 11452
rect 37282 11450 37306 11452
rect 37362 11450 37368 11452
rect 37122 11398 37124 11450
rect 37304 11398 37306 11450
rect 37060 11396 37066 11398
rect 37122 11396 37146 11398
rect 37202 11396 37226 11398
rect 37282 11396 37306 11398
rect 37362 11396 37368 11398
rect 37060 11387 37368 11396
rect 37372 11348 37424 11354
rect 37372 11290 37424 11296
rect 36728 11280 36780 11286
rect 36728 11222 36780 11228
rect 36740 10130 36768 11222
rect 36912 11212 36964 11218
rect 36912 11154 36964 11160
rect 36820 11008 36872 11014
rect 36820 10950 36872 10956
rect 36832 10266 36860 10950
rect 36924 10742 36952 11154
rect 37384 11150 37412 11290
rect 37476 11150 37504 11630
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37568 11286 37596 11562
rect 37556 11280 37608 11286
rect 37556 11222 37608 11228
rect 37372 11144 37424 11150
rect 37372 11086 37424 11092
rect 37464 11144 37516 11150
rect 37660 11098 37688 11630
rect 38028 11218 38056 11834
rect 38120 11354 38148 12106
rect 38292 11688 38344 11694
rect 38292 11630 38344 11636
rect 38108 11348 38160 11354
rect 38108 11290 38160 11296
rect 38016 11212 38068 11218
rect 38304 11200 38332 11630
rect 38488 11354 38516 12582
rect 38476 11348 38528 11354
rect 38476 11290 38528 11296
rect 38384 11212 38436 11218
rect 38304 11172 38384 11200
rect 38016 11154 38068 11160
rect 38384 11154 38436 11160
rect 37464 11086 37516 11092
rect 36912 10736 36964 10742
rect 36912 10678 36964 10684
rect 37384 10674 37412 11086
rect 37568 11070 37688 11098
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 37372 10668 37424 10674
rect 37424 10628 37504 10656
rect 37372 10610 37424 10616
rect 37060 10364 37368 10373
rect 37060 10362 37066 10364
rect 37122 10362 37146 10364
rect 37202 10362 37226 10364
rect 37282 10362 37306 10364
rect 37362 10362 37368 10364
rect 37122 10310 37124 10362
rect 37304 10310 37306 10362
rect 37060 10308 37066 10310
rect 37122 10308 37146 10310
rect 37202 10308 37226 10310
rect 37282 10308 37306 10310
rect 37362 10308 37368 10310
rect 37060 10299 37368 10308
rect 37476 10266 37504 10628
rect 37568 10538 37596 11070
rect 38488 11014 38516 11086
rect 38476 11008 38528 11014
rect 38476 10950 38528 10956
rect 37648 10668 37700 10674
rect 37648 10610 37700 10616
rect 37556 10532 37608 10538
rect 37556 10474 37608 10480
rect 36820 10260 36872 10266
rect 36820 10202 36872 10208
rect 37464 10260 37516 10266
rect 37464 10202 37516 10208
rect 37660 10198 37688 10610
rect 37740 10464 37792 10470
rect 37740 10406 37792 10412
rect 37648 10192 37700 10198
rect 37648 10134 37700 10140
rect 36728 10124 36780 10130
rect 36728 10066 36780 10072
rect 36636 9580 36688 9586
rect 36636 9522 36688 9528
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36464 8498 36492 9114
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36452 7948 36504 7954
rect 36452 7890 36504 7896
rect 36464 7546 36492 7890
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36544 7404 36596 7410
rect 36464 7364 36544 7392
rect 36464 7206 36492 7364
rect 36544 7346 36596 7352
rect 36452 7200 36504 7206
rect 36452 7142 36504 7148
rect 36360 6928 36412 6934
rect 36360 6870 36412 6876
rect 36268 6860 36320 6866
rect 36268 6802 36320 6808
rect 36280 6390 36308 6802
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 36176 6248 36228 6254
rect 36176 6190 36228 6196
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35808 5228 35860 5234
rect 35808 5170 35860 5176
rect 35820 5030 35848 5170
rect 35808 5024 35860 5030
rect 35808 4966 35860 4972
rect 35624 4684 35676 4690
rect 35624 4626 35676 4632
rect 35716 4616 35768 4622
rect 35716 4558 35768 4564
rect 34704 4072 34756 4078
rect 35348 4072 35400 4078
rect 34704 4014 34756 4020
rect 35346 4040 35348 4049
rect 35400 4040 35402 4049
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 34152 2848 34204 2854
rect 34152 2790 34204 2796
rect 34348 2514 34468 2530
rect 34348 2508 34480 2514
rect 34348 2502 34428 2508
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 870 34192 898
rect 34072 800 34100 870
rect 26620 734 26832 762
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34164 762 34192 870
rect 34348 762 34376 2502
rect 34428 2450 34480 2456
rect 34716 2446 34744 4014
rect 35346 3975 35402 3984
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 35636 3058 35664 3946
rect 35440 3052 35492 3058
rect 35624 3052 35676 3058
rect 35492 3012 35572 3040
rect 35440 2994 35492 3000
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 35360 2774 35388 2926
rect 35544 2774 35572 3012
rect 35624 2994 35676 3000
rect 35728 2990 35756 4558
rect 35900 4548 35952 4554
rect 35900 4490 35952 4496
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 35360 2746 35480 2774
rect 35544 2746 35664 2774
rect 35452 2582 35480 2746
rect 35440 2576 35492 2582
rect 35440 2518 35492 2524
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 34612 2100 34664 2106
rect 34612 2042 34664 2048
rect 34624 800 34652 2042
rect 35268 1306 35296 2382
rect 35636 2378 35664 2746
rect 35728 2650 35756 2926
rect 35716 2644 35768 2650
rect 35716 2586 35768 2592
rect 35716 2508 35768 2514
rect 35716 2450 35768 2456
rect 35624 2372 35676 2378
rect 35624 2314 35676 2320
rect 35176 1278 35296 1306
rect 35176 800 35204 1278
rect 35728 800 35756 2450
rect 35912 2310 35940 4490
rect 36096 4162 36124 5306
rect 36188 5234 36216 6190
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36188 4758 36216 5170
rect 36176 4752 36228 4758
rect 36176 4694 36228 4700
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 36004 4146 36124 4162
rect 35992 4140 36124 4146
rect 36044 4134 36124 4140
rect 35992 4082 36044 4088
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 36096 3738 36124 4014
rect 36188 3738 36216 4558
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 36176 3732 36228 3738
rect 36176 3674 36228 3680
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 3058 36032 3334
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 2650 36032 2790
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 35900 2304 35952 2310
rect 35900 2246 35952 2252
rect 36280 800 36308 4082
rect 36372 3194 36400 6870
rect 36464 6322 36492 7142
rect 36452 6316 36504 6322
rect 36452 6258 36504 6264
rect 36464 5302 36492 6258
rect 36544 6112 36596 6118
rect 36544 6054 36596 6060
rect 36556 5642 36584 6054
rect 36544 5636 36596 5642
rect 36544 5578 36596 5584
rect 36452 5296 36504 5302
rect 36452 5238 36504 5244
rect 36464 4758 36492 5238
rect 36452 4752 36504 4758
rect 36452 4694 36504 4700
rect 36556 4690 36584 5578
rect 36544 4684 36596 4690
rect 36544 4626 36596 4632
rect 36648 3942 36676 9522
rect 37752 9518 37780 10406
rect 38200 9580 38252 9586
rect 38200 9522 38252 9528
rect 37740 9512 37792 9518
rect 37740 9454 37792 9460
rect 38212 9382 38240 9522
rect 38290 9480 38346 9489
rect 38672 9450 38700 15302
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 39316 14074 39344 14758
rect 39304 14068 39356 14074
rect 39304 14010 39356 14016
rect 38844 13864 38896 13870
rect 38844 13806 38896 13812
rect 38752 13524 38804 13530
rect 38752 13466 38804 13472
rect 38764 13326 38792 13466
rect 38856 13433 38884 13806
rect 39120 13728 39172 13734
rect 39120 13670 39172 13676
rect 38842 13424 38898 13433
rect 38842 13359 38898 13368
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 38844 13320 38896 13326
rect 38844 13262 38896 13268
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 38856 13190 38884 13262
rect 38844 13184 38896 13190
rect 38844 13126 38896 13132
rect 38936 13184 38988 13190
rect 38936 13126 38988 13132
rect 38948 12374 38976 13126
rect 39040 12918 39068 13262
rect 39028 12912 39080 12918
rect 39028 12854 39080 12860
rect 38936 12368 38988 12374
rect 38936 12310 38988 12316
rect 38752 11008 38804 11014
rect 38752 10950 38804 10956
rect 38764 10062 38792 10950
rect 38844 10124 38896 10130
rect 38844 10066 38896 10072
rect 38752 10056 38804 10062
rect 38752 9998 38804 10004
rect 38856 9908 38884 10066
rect 38948 9926 38976 12310
rect 39132 11898 39160 13670
rect 39500 12434 39528 16952
rect 39856 16934 39908 16940
rect 39868 16794 39896 16934
rect 39856 16788 39908 16794
rect 39856 16730 39908 16736
rect 39764 14884 39816 14890
rect 39764 14826 39816 14832
rect 39776 14618 39804 14826
rect 39764 14612 39816 14618
rect 39764 14554 39816 14560
rect 39580 13864 39632 13870
rect 39580 13806 39632 13812
rect 39592 13394 39620 13806
rect 40052 13394 40080 19314
rect 40408 14408 40460 14414
rect 40408 14350 40460 14356
rect 40420 14074 40448 14350
rect 40408 14068 40460 14074
rect 40408 14010 40460 14016
rect 40512 13938 40540 19858
rect 43088 19854 43116 20470
rect 43272 20058 43300 21422
rect 43444 21344 43496 21350
rect 43444 21286 43496 21292
rect 43456 21146 43484 21286
rect 43444 21140 43496 21146
rect 43444 21082 43496 21088
rect 43812 20800 43864 20806
rect 43812 20742 43864 20748
rect 43260 20052 43312 20058
rect 43260 19994 43312 20000
rect 43720 19984 43772 19990
rect 43720 19926 43772 19932
rect 43352 19916 43404 19922
rect 43352 19858 43404 19864
rect 43628 19916 43680 19922
rect 43628 19858 43680 19864
rect 43076 19848 43128 19854
rect 43076 19790 43128 19796
rect 42984 19712 43036 19718
rect 42984 19654 43036 19660
rect 42248 19304 42300 19310
rect 42248 19246 42300 19252
rect 42708 19304 42760 19310
rect 42760 19252 42840 19258
rect 42708 19246 42840 19252
rect 41604 19168 41656 19174
rect 41604 19110 41656 19116
rect 41420 18964 41472 18970
rect 41420 18906 41472 18912
rect 41144 18692 41196 18698
rect 41144 18634 41196 18640
rect 41156 18290 41184 18634
rect 41432 18358 41460 18906
rect 41616 18698 41644 19110
rect 42260 18970 42288 19246
rect 42720 19230 42840 19246
rect 42248 18964 42300 18970
rect 42248 18906 42300 18912
rect 41604 18692 41656 18698
rect 41604 18634 41656 18640
rect 42064 18624 42116 18630
rect 42064 18566 42116 18572
rect 41420 18352 41472 18358
rect 41420 18294 41472 18300
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 41604 16992 41656 16998
rect 41604 16934 41656 16940
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 41248 16250 41276 16458
rect 41236 16244 41288 16250
rect 41236 16186 41288 16192
rect 41328 16040 41380 16046
rect 41064 16000 41328 16028
rect 41064 15910 41092 16000
rect 41328 15982 41380 15988
rect 41052 15904 41104 15910
rect 41052 15846 41104 15852
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 40224 13728 40276 13734
rect 40224 13670 40276 13676
rect 39580 13388 39632 13394
rect 39580 13330 39632 13336
rect 40040 13388 40092 13394
rect 40040 13330 40092 13336
rect 39592 12986 39620 13330
rect 39672 13184 39724 13190
rect 39672 13126 39724 13132
rect 39580 12980 39632 12986
rect 39580 12922 39632 12928
rect 39580 12844 39632 12850
rect 39580 12786 39632 12792
rect 39408 12406 39528 12434
rect 39120 11892 39172 11898
rect 39120 11834 39172 11840
rect 39212 11212 39264 11218
rect 39212 11154 39264 11160
rect 39224 10606 39252 11154
rect 39212 10600 39264 10606
rect 39212 10542 39264 10548
rect 38764 9880 38884 9908
rect 38936 9920 38988 9926
rect 38764 9586 38792 9880
rect 38936 9862 38988 9868
rect 39304 9920 39356 9926
rect 39304 9862 39356 9868
rect 39316 9654 39344 9862
rect 39304 9648 39356 9654
rect 39304 9590 39356 9596
rect 38752 9580 38804 9586
rect 38752 9522 38804 9528
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 38290 9415 38346 9424
rect 38660 9444 38712 9450
rect 38304 9382 38332 9415
rect 38660 9386 38712 9392
rect 37464 9376 37516 9382
rect 37464 9318 37516 9324
rect 38200 9376 38252 9382
rect 38200 9318 38252 9324
rect 38292 9376 38344 9382
rect 38292 9318 38344 9324
rect 37060 9276 37368 9285
rect 37060 9274 37066 9276
rect 37122 9274 37146 9276
rect 37202 9274 37226 9276
rect 37282 9274 37306 9276
rect 37362 9274 37368 9276
rect 37122 9222 37124 9274
rect 37304 9222 37306 9274
rect 37060 9220 37066 9222
rect 37122 9220 37146 9222
rect 37202 9220 37226 9222
rect 37282 9220 37306 9222
rect 37362 9220 37368 9222
rect 37060 9211 37368 9220
rect 36728 8968 36780 8974
rect 36728 8910 36780 8916
rect 36740 8634 36768 8910
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 36728 8628 36780 8634
rect 36728 8570 36780 8576
rect 36728 8288 36780 8294
rect 36728 8230 36780 8236
rect 36740 7886 36768 8230
rect 36924 7954 36952 8774
rect 37060 8188 37368 8197
rect 37060 8186 37066 8188
rect 37122 8186 37146 8188
rect 37202 8186 37226 8188
rect 37282 8186 37306 8188
rect 37362 8186 37368 8188
rect 37122 8134 37124 8186
rect 37304 8134 37306 8186
rect 37060 8132 37066 8134
rect 37122 8132 37146 8134
rect 37202 8132 37226 8134
rect 37282 8132 37306 8134
rect 37362 8132 37368 8134
rect 37060 8123 37368 8132
rect 36912 7948 36964 7954
rect 36912 7890 36964 7896
rect 37188 7948 37240 7954
rect 37188 7890 37240 7896
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36820 7540 36872 7546
rect 36820 7482 36872 7488
rect 36728 7336 36780 7342
rect 36728 7278 36780 7284
rect 36740 5302 36768 7278
rect 36832 6934 36860 7482
rect 37200 7410 37228 7890
rect 37188 7404 37240 7410
rect 37188 7346 37240 7352
rect 37060 7100 37368 7109
rect 37060 7098 37066 7100
rect 37122 7098 37146 7100
rect 37202 7098 37226 7100
rect 37282 7098 37306 7100
rect 37362 7098 37368 7100
rect 37122 7046 37124 7098
rect 37304 7046 37306 7098
rect 37060 7044 37066 7046
rect 37122 7044 37146 7046
rect 37202 7044 37226 7046
rect 37282 7044 37306 7046
rect 37362 7044 37368 7046
rect 37060 7035 37368 7044
rect 36820 6928 36872 6934
rect 36820 6870 36872 6876
rect 37188 6928 37240 6934
rect 37188 6870 37240 6876
rect 37200 6458 37228 6870
rect 37188 6452 37240 6458
rect 37188 6394 37240 6400
rect 37476 6322 37504 9318
rect 37648 9172 37700 9178
rect 37648 9114 37700 9120
rect 37660 7954 37688 9114
rect 37740 8288 37792 8294
rect 37740 8230 37792 8236
rect 37752 7954 37780 8230
rect 37648 7948 37700 7954
rect 37648 7890 37700 7896
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 38016 7948 38068 7954
rect 38016 7890 38068 7896
rect 37648 7744 37700 7750
rect 37648 7686 37700 7692
rect 37924 7744 37976 7750
rect 37924 7686 37976 7692
rect 37556 6724 37608 6730
rect 37556 6666 37608 6672
rect 37464 6316 37516 6322
rect 37464 6258 37516 6264
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 36924 5710 36952 6054
rect 37060 6012 37368 6021
rect 37060 6010 37066 6012
rect 37122 6010 37146 6012
rect 37202 6010 37226 6012
rect 37282 6010 37306 6012
rect 37362 6010 37368 6012
rect 37122 5958 37124 6010
rect 37304 5958 37306 6010
rect 37060 5956 37066 5958
rect 37122 5956 37146 5958
rect 37202 5956 37226 5958
rect 37282 5956 37306 5958
rect 37362 5956 37368 5958
rect 37060 5947 37368 5956
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 37108 5370 37136 5510
rect 37096 5364 37148 5370
rect 37096 5306 37148 5312
rect 36728 5296 36780 5302
rect 36728 5238 36780 5244
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 36924 4672 36952 4966
rect 37060 4924 37368 4933
rect 37060 4922 37066 4924
rect 37122 4922 37146 4924
rect 37202 4922 37226 4924
rect 37282 4922 37306 4924
rect 37362 4922 37368 4924
rect 37122 4870 37124 4922
rect 37304 4870 37306 4922
rect 37060 4868 37066 4870
rect 37122 4868 37146 4870
rect 37202 4868 37226 4870
rect 37282 4868 37306 4870
rect 37362 4868 37368 4870
rect 37060 4859 37368 4868
rect 37004 4684 37056 4690
rect 36924 4644 37004 4672
rect 37004 4626 37056 4632
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 36832 4078 36860 4558
rect 37476 4282 37504 6258
rect 37568 5710 37596 6666
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 37568 5250 37596 5646
rect 37660 5370 37688 7686
rect 37740 7472 37792 7478
rect 37740 7414 37792 7420
rect 37752 7188 37780 7414
rect 37936 7410 37964 7686
rect 37924 7404 37976 7410
rect 37924 7346 37976 7352
rect 38028 7342 38056 7890
rect 38108 7472 38160 7478
rect 38108 7414 38160 7420
rect 38016 7336 38068 7342
rect 38016 7278 38068 7284
rect 38120 7188 38148 7414
rect 38212 7342 38240 9318
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 38292 8288 38344 8294
rect 38292 8230 38344 8236
rect 38304 7818 38332 8230
rect 38292 7812 38344 7818
rect 38292 7754 38344 7760
rect 38200 7336 38252 7342
rect 38200 7278 38252 7284
rect 37752 7160 38148 7188
rect 38304 6662 38332 7754
rect 38396 7546 38424 8434
rect 38476 8084 38528 8090
rect 38476 8026 38528 8032
rect 38488 7546 38516 8026
rect 38384 7540 38436 7546
rect 38384 7482 38436 7488
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38474 7440 38530 7449
rect 38474 7375 38476 7384
rect 38528 7375 38530 7384
rect 38476 7346 38528 7352
rect 38384 7336 38436 7342
rect 38384 7278 38436 7284
rect 38292 6656 38344 6662
rect 38292 6598 38344 6604
rect 38304 5914 38332 6598
rect 38108 5908 38160 5914
rect 38108 5850 38160 5856
rect 38292 5908 38344 5914
rect 38292 5850 38344 5856
rect 37924 5636 37976 5642
rect 37924 5578 37976 5584
rect 37648 5364 37700 5370
rect 37648 5306 37700 5312
rect 37568 5222 37688 5250
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37096 4140 37148 4146
rect 36924 4100 37096 4128
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 36636 3936 36688 3942
rect 36636 3878 36688 3884
rect 36818 3904 36874 3913
rect 36818 3839 36874 3848
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36832 3058 36860 3839
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 36372 2854 36400 2994
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36924 2632 36952 4100
rect 37096 4082 37148 4088
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37060 3836 37368 3845
rect 37060 3834 37066 3836
rect 37122 3834 37146 3836
rect 37202 3834 37226 3836
rect 37282 3834 37306 3836
rect 37362 3834 37368 3836
rect 37122 3782 37124 3834
rect 37304 3782 37306 3834
rect 37060 3780 37066 3782
rect 37122 3780 37146 3782
rect 37202 3780 37226 3782
rect 37282 3780 37306 3782
rect 37362 3780 37368 3782
rect 37060 3771 37368 3780
rect 37476 3466 37504 3878
rect 37464 3460 37516 3466
rect 37464 3402 37516 3408
rect 37568 3398 37596 4966
rect 37660 3534 37688 5222
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 37752 4826 37780 5102
rect 37936 4826 37964 5578
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 38028 4826 38056 4966
rect 37740 4820 37792 4826
rect 37740 4762 37792 4768
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 37832 4072 37884 4078
rect 37832 4014 37884 4020
rect 37844 3738 37872 4014
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37924 3732 37976 3738
rect 37924 3674 37976 3680
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37060 2748 37368 2757
rect 37060 2746 37066 2748
rect 37122 2746 37146 2748
rect 37202 2746 37226 2748
rect 37282 2746 37306 2748
rect 37362 2746 37368 2748
rect 37122 2694 37124 2746
rect 37304 2694 37306 2746
rect 37060 2692 37066 2694
rect 37122 2692 37146 2694
rect 37202 2692 37226 2694
rect 37282 2692 37306 2694
rect 37362 2692 37368 2694
rect 37060 2683 37368 2692
rect 37004 2644 37056 2650
rect 36924 2604 37004 2632
rect 37004 2586 37056 2592
rect 37476 2446 37504 2790
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 36820 2304 36872 2310
rect 36820 2246 36872 2252
rect 36832 800 36860 2246
rect 37108 1426 37136 2382
rect 37096 1420 37148 1426
rect 37096 1362 37148 1368
rect 37384 870 37504 898
rect 37384 800 37412 870
rect 34164 734 34376 762
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37476 762 37504 870
rect 37660 762 37688 2926
rect 37936 800 37964 3674
rect 38120 3602 38148 5850
rect 38292 4480 38344 4486
rect 38292 4422 38344 4428
rect 38304 4282 38332 4422
rect 38292 4276 38344 4282
rect 38292 4218 38344 4224
rect 38396 3602 38424 7278
rect 38476 7200 38528 7206
rect 38476 7142 38528 7148
rect 38752 7200 38804 7206
rect 38752 7142 38804 7148
rect 38488 5914 38516 7142
rect 38660 6724 38712 6730
rect 38660 6666 38712 6672
rect 38568 6656 38620 6662
rect 38568 6598 38620 6604
rect 38476 5908 38528 5914
rect 38476 5850 38528 5856
rect 38488 3602 38516 5850
rect 38580 5846 38608 6598
rect 38672 6254 38700 6666
rect 38660 6248 38712 6254
rect 38660 6190 38712 6196
rect 38672 5914 38700 6190
rect 38764 6186 38792 7142
rect 38752 6180 38804 6186
rect 38752 6122 38804 6128
rect 38660 5908 38712 5914
rect 38660 5850 38712 5856
rect 38568 5840 38620 5846
rect 38568 5782 38620 5788
rect 38672 5234 38700 5850
rect 38764 5778 38792 6122
rect 38752 5772 38804 5778
rect 38752 5714 38804 5720
rect 38752 5568 38804 5574
rect 38752 5510 38804 5516
rect 38660 5228 38712 5234
rect 38660 5170 38712 5176
rect 38764 5166 38792 5510
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 38856 4826 38884 9522
rect 39120 9376 39172 9382
rect 39120 9318 39172 9324
rect 39132 9110 39160 9318
rect 39120 9104 39172 9110
rect 39120 9046 39172 9052
rect 38936 8968 38988 8974
rect 38936 8910 38988 8916
rect 38948 8634 38976 8910
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 39028 7744 39080 7750
rect 39028 7686 39080 7692
rect 39040 7206 39068 7686
rect 39028 7200 39080 7206
rect 39028 7142 39080 7148
rect 39120 6656 39172 6662
rect 39120 6598 39172 6604
rect 39132 6322 39160 6598
rect 39120 6316 39172 6322
rect 39120 6258 39172 6264
rect 38844 4820 38896 4826
rect 38844 4762 38896 4768
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 38384 3596 38436 3602
rect 38384 3538 38436 3544
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 38488 3194 38516 3538
rect 38672 3534 38700 4082
rect 39408 3534 39436 12406
rect 39592 11898 39620 12786
rect 39684 11898 39712 13126
rect 40052 12753 40080 13330
rect 40236 13326 40264 13670
rect 40512 13530 40540 13874
rect 40500 13524 40552 13530
rect 40500 13466 40552 13472
rect 40224 13320 40276 13326
rect 40224 13262 40276 13268
rect 40316 13320 40368 13326
rect 40316 13262 40368 13268
rect 40328 12782 40356 13262
rect 40592 13184 40644 13190
rect 40592 13126 40644 13132
rect 40604 12782 40632 13126
rect 41064 13025 41092 15846
rect 41236 15428 41288 15434
rect 41236 15370 41288 15376
rect 41248 15162 41276 15370
rect 41236 15156 41288 15162
rect 41236 15098 41288 15104
rect 41616 14006 41644 16934
rect 41788 16448 41840 16454
rect 41788 16390 41840 16396
rect 41800 16250 41828 16390
rect 41788 16244 41840 16250
rect 41788 16186 41840 16192
rect 42076 15910 42104 18566
rect 42616 18352 42668 18358
rect 42616 18294 42668 18300
rect 42248 18284 42300 18290
rect 42248 18226 42300 18232
rect 42260 16454 42288 18226
rect 42524 18216 42576 18222
rect 42524 18158 42576 18164
rect 42536 18086 42564 18158
rect 42524 18080 42576 18086
rect 42524 18022 42576 18028
rect 42536 17542 42564 18022
rect 42628 17814 42656 18294
rect 42616 17808 42668 17814
rect 42616 17750 42668 17756
rect 42524 17536 42576 17542
rect 42524 17478 42576 17484
rect 42708 17536 42760 17542
rect 42708 17478 42760 17484
rect 42340 16992 42392 16998
rect 42340 16934 42392 16940
rect 42432 16992 42484 16998
rect 42432 16934 42484 16940
rect 42352 16658 42380 16934
rect 42444 16794 42472 16934
rect 42432 16788 42484 16794
rect 42432 16730 42484 16736
rect 42340 16652 42392 16658
rect 42340 16594 42392 16600
rect 42248 16448 42300 16454
rect 42248 16390 42300 16396
rect 42064 15904 42116 15910
rect 42064 15846 42116 15852
rect 42156 15564 42208 15570
rect 42156 15506 42208 15512
rect 41788 15360 41840 15366
rect 41788 15302 41840 15308
rect 41800 15026 41828 15302
rect 41788 15020 41840 15026
rect 41788 14962 41840 14968
rect 42168 14822 42196 15506
rect 42260 15502 42288 16390
rect 42616 15972 42668 15978
rect 42616 15914 42668 15920
rect 42628 15706 42656 15914
rect 42616 15700 42668 15706
rect 42616 15642 42668 15648
rect 42248 15496 42300 15502
rect 42248 15438 42300 15444
rect 42156 14816 42208 14822
rect 42156 14758 42208 14764
rect 41604 14000 41656 14006
rect 41604 13942 41656 13948
rect 41604 13252 41656 13258
rect 41604 13194 41656 13200
rect 41050 13016 41106 13025
rect 41616 12986 41644 13194
rect 41050 12951 41106 12960
rect 41604 12980 41656 12986
rect 41604 12922 41656 12928
rect 40316 12776 40368 12782
rect 40038 12744 40094 12753
rect 40316 12718 40368 12724
rect 40592 12776 40644 12782
rect 40592 12718 40644 12724
rect 41236 12776 41288 12782
rect 41236 12718 41288 12724
rect 40038 12679 40094 12688
rect 40052 12434 40080 12679
rect 40052 12406 40264 12434
rect 40236 12102 40264 12406
rect 40328 12170 40356 12718
rect 41248 12238 41276 12718
rect 42168 12442 42196 14758
rect 42524 14272 42576 14278
rect 42524 14214 42576 14220
rect 42248 13728 42300 13734
rect 42248 13670 42300 13676
rect 42260 12714 42288 13670
rect 42536 13394 42564 14214
rect 42616 13864 42668 13870
rect 42616 13806 42668 13812
rect 42524 13388 42576 13394
rect 42524 13330 42576 13336
rect 42340 13184 42392 13190
rect 42340 13126 42392 13132
rect 42352 12986 42380 13126
rect 42340 12980 42392 12986
rect 42340 12922 42392 12928
rect 42628 12782 42656 13806
rect 42616 12776 42668 12782
rect 42616 12718 42668 12724
rect 42248 12708 42300 12714
rect 42248 12650 42300 12656
rect 42156 12436 42208 12442
rect 42156 12378 42208 12384
rect 42720 12306 42748 17478
rect 42812 16028 42840 19230
rect 42996 18630 43024 19654
rect 43088 18834 43116 19790
rect 43364 19514 43392 19858
rect 43352 19508 43404 19514
rect 43352 19450 43404 19456
rect 43260 19304 43312 19310
rect 43260 19246 43312 19252
rect 43076 18828 43128 18834
rect 43128 18788 43208 18816
rect 43076 18770 43128 18776
rect 42984 18624 43036 18630
rect 42984 18566 43036 18572
rect 42996 18358 43024 18566
rect 42984 18352 43036 18358
rect 42984 18294 43036 18300
rect 42984 17128 43036 17134
rect 42984 17070 43036 17076
rect 42996 16590 43024 17070
rect 42984 16584 43036 16590
rect 42984 16526 43036 16532
rect 42892 16040 42944 16046
rect 42812 16000 42892 16028
rect 42892 15982 42944 15988
rect 43076 16040 43128 16046
rect 43076 15982 43128 15988
rect 43088 15434 43116 15982
rect 43076 15428 43128 15434
rect 43076 15370 43128 15376
rect 43076 14408 43128 14414
rect 43076 14350 43128 14356
rect 43088 13258 43116 14350
rect 43180 13734 43208 18788
rect 43272 18154 43300 19246
rect 43640 19242 43668 19858
rect 43732 19825 43760 19926
rect 43824 19922 43852 20742
rect 44008 20058 44036 21422
rect 44100 21010 44128 21422
rect 44824 21344 44876 21350
rect 44824 21286 44876 21292
rect 45836 21344 45888 21350
rect 45836 21286 45888 21292
rect 44088 21004 44140 21010
rect 44088 20946 44140 20952
rect 43996 20052 44048 20058
rect 43996 19994 44048 20000
rect 43812 19916 43864 19922
rect 43812 19858 43864 19864
rect 43718 19816 43774 19825
rect 43718 19751 43774 19760
rect 44100 19378 44128 20946
rect 44180 20936 44232 20942
rect 44180 20878 44232 20884
rect 44192 20602 44220 20878
rect 44282 20700 44590 20709
rect 44282 20698 44288 20700
rect 44344 20698 44368 20700
rect 44424 20698 44448 20700
rect 44504 20698 44528 20700
rect 44584 20698 44590 20700
rect 44344 20646 44346 20698
rect 44526 20646 44528 20698
rect 44282 20644 44288 20646
rect 44344 20644 44368 20646
rect 44424 20644 44448 20646
rect 44504 20644 44528 20646
rect 44584 20644 44590 20646
rect 44282 20635 44590 20644
rect 44180 20596 44232 20602
rect 44180 20538 44232 20544
rect 44192 19378 44220 20538
rect 44640 19916 44692 19922
rect 44640 19858 44692 19864
rect 44282 19612 44590 19621
rect 44282 19610 44288 19612
rect 44344 19610 44368 19612
rect 44424 19610 44448 19612
rect 44504 19610 44528 19612
rect 44584 19610 44590 19612
rect 44344 19558 44346 19610
rect 44526 19558 44528 19610
rect 44282 19556 44288 19558
rect 44344 19556 44368 19558
rect 44424 19556 44448 19558
rect 44504 19556 44528 19558
rect 44584 19556 44590 19558
rect 44282 19547 44590 19556
rect 44652 19446 44680 19858
rect 44836 19854 44864 21286
rect 45008 20800 45060 20806
rect 45008 20742 45060 20748
rect 45020 20262 45048 20742
rect 45744 20460 45796 20466
rect 45744 20402 45796 20408
rect 45008 20256 45060 20262
rect 45008 20198 45060 20204
rect 45020 19854 45048 20198
rect 44824 19848 44876 19854
rect 44824 19790 44876 19796
rect 45008 19848 45060 19854
rect 45008 19790 45060 19796
rect 44640 19440 44692 19446
rect 44640 19382 44692 19388
rect 44088 19372 44140 19378
rect 44088 19314 44140 19320
rect 44180 19372 44232 19378
rect 44180 19314 44232 19320
rect 43628 19236 43680 19242
rect 43628 19178 43680 19184
rect 43640 18970 43668 19178
rect 43720 19168 43772 19174
rect 43720 19110 43772 19116
rect 43812 19168 43864 19174
rect 43812 19110 43864 19116
rect 44180 19168 44232 19174
rect 44180 19110 44232 19116
rect 44916 19168 44968 19174
rect 44916 19110 44968 19116
rect 43628 18964 43680 18970
rect 43628 18906 43680 18912
rect 43260 18148 43312 18154
rect 43260 18090 43312 18096
rect 43444 17536 43496 17542
rect 43444 17478 43496 17484
rect 43456 17134 43484 17478
rect 43640 17218 43668 18906
rect 43732 17338 43760 19110
rect 43824 18834 43852 19110
rect 43812 18828 43864 18834
rect 43812 18770 43864 18776
rect 43996 18760 44048 18766
rect 43996 18702 44048 18708
rect 44008 18426 44036 18702
rect 43996 18420 44048 18426
rect 43996 18362 44048 18368
rect 43720 17332 43772 17338
rect 43720 17274 43772 17280
rect 43548 17190 43668 17218
rect 43444 17128 43496 17134
rect 43444 17070 43496 17076
rect 43352 16516 43404 16522
rect 43352 16458 43404 16464
rect 43364 16114 43392 16458
rect 43352 16108 43404 16114
rect 43352 16050 43404 16056
rect 43548 16046 43576 17190
rect 43628 17128 43680 17134
rect 43628 17070 43680 17076
rect 43640 16250 43668 17070
rect 43996 17060 44048 17066
rect 43996 17002 44048 17008
rect 44008 16590 44036 17002
rect 44088 16992 44140 16998
rect 44088 16934 44140 16940
rect 43996 16584 44048 16590
rect 43996 16526 44048 16532
rect 43628 16244 43680 16250
rect 43628 16186 43680 16192
rect 43260 16040 43312 16046
rect 43536 16040 43588 16046
rect 43260 15982 43312 15988
rect 43456 16000 43536 16028
rect 43272 15638 43300 15982
rect 43456 15706 43484 16000
rect 43536 15982 43588 15988
rect 43536 15904 43588 15910
rect 43536 15846 43588 15852
rect 43444 15700 43496 15706
rect 43444 15642 43496 15648
rect 43260 15632 43312 15638
rect 43260 15574 43312 15580
rect 43168 13728 43220 13734
rect 43168 13670 43220 13676
rect 43180 13394 43208 13670
rect 43168 13388 43220 13394
rect 43168 13330 43220 13336
rect 43076 13252 43128 13258
rect 43076 13194 43128 13200
rect 43088 12986 43116 13194
rect 43076 12980 43128 12986
rect 43076 12922 43128 12928
rect 43456 12434 43484 15642
rect 43548 15570 43576 15846
rect 43536 15564 43588 15570
rect 43536 15506 43588 15512
rect 43548 15162 43576 15506
rect 43536 15156 43588 15162
rect 43536 15098 43588 15104
rect 43812 14272 43864 14278
rect 43812 14214 43864 14220
rect 43824 13394 43852 14214
rect 43812 13388 43864 13394
rect 43812 13330 43864 13336
rect 43812 13184 43864 13190
rect 43812 13126 43864 13132
rect 43364 12406 43484 12434
rect 42524 12300 42576 12306
rect 42524 12242 42576 12248
rect 42708 12300 42760 12306
rect 42708 12242 42760 12248
rect 41236 12232 41288 12238
rect 41236 12174 41288 12180
rect 40316 12164 40368 12170
rect 40316 12106 40368 12112
rect 40224 12096 40276 12102
rect 40224 12038 40276 12044
rect 39580 11892 39632 11898
rect 39580 11834 39632 11840
rect 39672 11892 39724 11898
rect 39672 11834 39724 11840
rect 39856 11144 39908 11150
rect 39856 11086 39908 11092
rect 39868 10198 39896 11086
rect 39856 10192 39908 10198
rect 39856 10134 39908 10140
rect 39764 9648 39816 9654
rect 39764 9590 39816 9596
rect 39672 8832 39724 8838
rect 39672 8774 39724 8780
rect 39684 8634 39712 8774
rect 39776 8634 39804 9590
rect 39868 9586 39896 10134
rect 39856 9580 39908 9586
rect 39856 9522 39908 9528
rect 39672 8628 39724 8634
rect 39672 8570 39724 8576
rect 39764 8628 39816 8634
rect 39764 8570 39816 8576
rect 39672 8492 39724 8498
rect 39672 8434 39724 8440
rect 39684 4826 39712 8434
rect 40236 8430 40264 12038
rect 40776 11348 40828 11354
rect 40776 11290 40828 11296
rect 40788 10810 40816 11290
rect 41248 10810 41276 12174
rect 42432 12164 42484 12170
rect 42432 12106 42484 12112
rect 42444 11898 42472 12106
rect 42432 11892 42484 11898
rect 42432 11834 42484 11840
rect 42536 11830 42564 12242
rect 42708 12096 42760 12102
rect 42708 12038 42760 12044
rect 42892 12096 42944 12102
rect 42892 12038 42944 12044
rect 42720 11898 42748 12038
rect 42708 11892 42760 11898
rect 42708 11834 42760 11840
rect 42524 11824 42576 11830
rect 42524 11766 42576 11772
rect 41512 11552 41564 11558
rect 41512 11494 41564 11500
rect 40776 10804 40828 10810
rect 40776 10746 40828 10752
rect 41236 10804 41288 10810
rect 41236 10746 41288 10752
rect 40408 8968 40460 8974
rect 40408 8910 40460 8916
rect 40316 8900 40368 8906
rect 40316 8842 40368 8848
rect 40224 8424 40276 8430
rect 40224 8366 40276 8372
rect 40132 7336 40184 7342
rect 40132 7278 40184 7284
rect 39856 7268 39908 7274
rect 39856 7210 39908 7216
rect 39868 7041 39896 7210
rect 40144 7177 40172 7278
rect 40130 7168 40186 7177
rect 40130 7103 40186 7112
rect 39854 7032 39910 7041
rect 39854 6967 39910 6976
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 39764 6112 39816 6118
rect 39764 6054 39816 6060
rect 39776 5642 39804 6054
rect 40144 5778 40172 6734
rect 40236 5778 40264 8366
rect 40328 7818 40356 8842
rect 40420 8498 40448 8910
rect 40500 8832 40552 8838
rect 40500 8774 40552 8780
rect 40512 8566 40540 8774
rect 40500 8560 40552 8566
rect 40500 8502 40552 8508
rect 40408 8492 40460 8498
rect 40408 8434 40460 8440
rect 40512 7886 40540 8502
rect 40500 7880 40552 7886
rect 40500 7822 40552 7828
rect 40316 7812 40368 7818
rect 40316 7754 40368 7760
rect 40132 5772 40184 5778
rect 40132 5714 40184 5720
rect 40224 5772 40276 5778
rect 40224 5714 40276 5720
rect 39764 5636 39816 5642
rect 39764 5578 39816 5584
rect 39672 4820 39724 4826
rect 39672 4762 39724 4768
rect 39856 4480 39908 4486
rect 39856 4422 39908 4428
rect 39868 4214 39896 4422
rect 40144 4214 40172 5714
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 39856 4208 39908 4214
rect 39856 4150 39908 4156
rect 40132 4208 40184 4214
rect 40132 4150 40184 4156
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39946 4040 40002 4049
rect 38660 3528 38712 3534
rect 38660 3470 38712 3476
rect 39396 3528 39448 3534
rect 39396 3470 39448 3476
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38672 3058 38700 3470
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38476 2984 38528 2990
rect 38476 2926 38528 2932
rect 38488 800 38516 2926
rect 39120 2372 39172 2378
rect 39120 2314 39172 2320
rect 39132 1170 39160 2314
rect 39040 1142 39160 1170
rect 39040 800 39068 1142
rect 39592 800 39620 4014
rect 39946 3975 40002 3984
rect 39960 3602 39988 3975
rect 40144 3602 40172 4150
rect 40236 4010 40264 4626
rect 40224 4004 40276 4010
rect 40224 3946 40276 3952
rect 40328 3942 40356 7754
rect 40684 7472 40736 7478
rect 40682 7440 40684 7449
rect 40736 7440 40738 7449
rect 40408 7404 40460 7410
rect 40682 7375 40738 7384
rect 40408 7346 40460 7352
rect 40420 6866 40448 7346
rect 40500 7336 40552 7342
rect 40500 7278 40552 7284
rect 40408 6860 40460 6866
rect 40408 6802 40460 6808
rect 40420 6322 40448 6802
rect 40512 6390 40540 7278
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40408 6316 40460 6322
rect 40408 6258 40460 6264
rect 40512 5370 40540 6326
rect 40788 5710 40816 10746
rect 41248 10130 41276 10746
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 41144 9988 41196 9994
rect 41144 9930 41196 9936
rect 41156 9722 41184 9930
rect 41144 9716 41196 9722
rect 41144 9658 41196 9664
rect 41524 9602 41552 11494
rect 42904 11014 42932 12038
rect 43260 11552 43312 11558
rect 43260 11494 43312 11500
rect 43272 11286 43300 11494
rect 43260 11280 43312 11286
rect 43260 11222 43312 11228
rect 42524 11008 42576 11014
rect 42524 10950 42576 10956
rect 42892 11008 42944 11014
rect 42892 10950 42944 10956
rect 42536 10674 42564 10950
rect 42432 10668 42484 10674
rect 42432 10610 42484 10616
rect 42524 10668 42576 10674
rect 42524 10610 42576 10616
rect 41604 9988 41656 9994
rect 41604 9930 41656 9936
rect 41616 9722 41644 9930
rect 42444 9722 42472 10610
rect 41604 9716 41656 9722
rect 41604 9658 41656 9664
rect 42432 9716 42484 9722
rect 42432 9658 42484 9664
rect 41524 9574 41644 9602
rect 42904 9586 42932 10950
rect 43364 9586 43392 12406
rect 43824 12102 43852 13126
rect 43996 12980 44048 12986
rect 43996 12922 44048 12928
rect 44008 12850 44036 12922
rect 43904 12844 43956 12850
rect 43904 12786 43956 12792
rect 43996 12844 44048 12850
rect 43996 12786 44048 12792
rect 43916 12374 43944 12786
rect 43904 12368 43956 12374
rect 43904 12310 43956 12316
rect 43996 12300 44048 12306
rect 43996 12242 44048 12248
rect 43812 12096 43864 12102
rect 43812 12038 43864 12044
rect 44008 11898 44036 12242
rect 43996 11892 44048 11898
rect 43996 11834 44048 11840
rect 43628 11620 43680 11626
rect 43628 11562 43680 11568
rect 43720 11620 43772 11626
rect 43720 11562 43772 11568
rect 43640 11286 43668 11562
rect 43628 11280 43680 11286
rect 43628 11222 43680 11228
rect 43732 10742 43760 11562
rect 44100 11234 44128 16934
rect 44192 16454 44220 19110
rect 44282 18524 44590 18533
rect 44282 18522 44288 18524
rect 44344 18522 44368 18524
rect 44424 18522 44448 18524
rect 44504 18522 44528 18524
rect 44584 18522 44590 18524
rect 44344 18470 44346 18522
rect 44526 18470 44528 18522
rect 44282 18468 44288 18470
rect 44344 18468 44368 18470
rect 44424 18468 44448 18470
rect 44504 18468 44528 18470
rect 44584 18468 44590 18470
rect 44282 18459 44590 18468
rect 44282 17436 44590 17445
rect 44282 17434 44288 17436
rect 44344 17434 44368 17436
rect 44424 17434 44448 17436
rect 44504 17434 44528 17436
rect 44584 17434 44590 17436
rect 44344 17382 44346 17434
rect 44526 17382 44528 17434
rect 44282 17380 44288 17382
rect 44344 17380 44368 17382
rect 44424 17380 44448 17382
rect 44504 17380 44528 17382
rect 44584 17380 44590 17382
rect 44282 17371 44590 17380
rect 44272 17128 44324 17134
rect 44272 17070 44324 17076
rect 44284 16726 44312 17070
rect 44824 16992 44876 16998
rect 44824 16934 44876 16940
rect 44272 16720 44324 16726
rect 44272 16662 44324 16668
rect 44640 16720 44692 16726
rect 44640 16662 44692 16668
rect 44180 16448 44232 16454
rect 44180 16390 44232 16396
rect 44192 11830 44220 16390
rect 44282 16348 44590 16357
rect 44282 16346 44288 16348
rect 44344 16346 44368 16348
rect 44424 16346 44448 16348
rect 44504 16346 44528 16348
rect 44584 16346 44590 16348
rect 44344 16294 44346 16346
rect 44526 16294 44528 16346
rect 44282 16292 44288 16294
rect 44344 16292 44368 16294
rect 44424 16292 44448 16294
rect 44504 16292 44528 16294
rect 44584 16292 44590 16294
rect 44282 16283 44590 16292
rect 44652 16114 44680 16662
rect 44836 16590 44864 16934
rect 44824 16584 44876 16590
rect 44824 16526 44876 16532
rect 44928 16436 44956 19110
rect 45020 18426 45048 19790
rect 45284 19372 45336 19378
rect 45284 19314 45336 19320
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 45020 17882 45048 18362
rect 45008 17876 45060 17882
rect 45008 17818 45060 17824
rect 45296 17678 45324 19314
rect 45756 19242 45784 20402
rect 45744 19236 45796 19242
rect 45744 19178 45796 19184
rect 45848 18086 45876 21286
rect 46124 21146 46152 21422
rect 46940 21412 46992 21418
rect 46940 21354 46992 21360
rect 46480 21344 46532 21350
rect 46480 21286 46532 21292
rect 46756 21344 46808 21350
rect 46756 21286 46808 21292
rect 46112 21140 46164 21146
rect 46112 21082 46164 21088
rect 46492 21010 46520 21286
rect 46480 21004 46532 21010
rect 46480 20946 46532 20952
rect 46768 20534 46796 21286
rect 46952 21010 46980 21354
rect 47584 21344 47636 21350
rect 47584 21286 47636 21292
rect 47596 21146 47624 21286
rect 47584 21140 47636 21146
rect 47584 21082 47636 21088
rect 46940 21004 46992 21010
rect 46940 20946 46992 20952
rect 46952 20534 46980 20946
rect 47768 20936 47820 20942
rect 47768 20878 47820 20884
rect 47492 20800 47544 20806
rect 47492 20742 47544 20748
rect 46756 20528 46808 20534
rect 46756 20470 46808 20476
rect 46940 20528 46992 20534
rect 46940 20470 46992 20476
rect 45928 20392 45980 20398
rect 45928 20334 45980 20340
rect 45940 19854 45968 20334
rect 47504 19922 47532 20742
rect 47780 20262 47808 20878
rect 48240 20602 48268 21422
rect 48504 21344 48556 21350
rect 48504 21286 48556 21292
rect 48228 20596 48280 20602
rect 48228 20538 48280 20544
rect 48240 20482 48268 20538
rect 48240 20466 48360 20482
rect 48240 20460 48372 20466
rect 48240 20454 48320 20460
rect 48320 20402 48372 20408
rect 47584 20256 47636 20262
rect 47584 20198 47636 20204
rect 47676 20256 47728 20262
rect 47676 20198 47728 20204
rect 47768 20256 47820 20262
rect 47768 20198 47820 20204
rect 47596 19990 47624 20198
rect 47584 19984 47636 19990
rect 47584 19926 47636 19932
rect 47492 19916 47544 19922
rect 47492 19858 47544 19864
rect 45928 19848 45980 19854
rect 45928 19790 45980 19796
rect 47400 19848 47452 19854
rect 47400 19790 47452 19796
rect 46020 19304 46072 19310
rect 46020 19246 46072 19252
rect 46032 18970 46060 19246
rect 46020 18964 46072 18970
rect 46020 18906 46072 18912
rect 46756 18828 46808 18834
rect 46756 18770 46808 18776
rect 46020 18624 46072 18630
rect 46020 18566 46072 18572
rect 46204 18624 46256 18630
rect 46204 18566 46256 18572
rect 46388 18624 46440 18630
rect 46388 18566 46440 18572
rect 46664 18624 46716 18630
rect 46664 18566 46716 18572
rect 45836 18080 45888 18086
rect 45836 18022 45888 18028
rect 46032 17882 46060 18566
rect 46216 18426 46244 18566
rect 46400 18426 46428 18566
rect 46676 18426 46704 18566
rect 46204 18420 46256 18426
rect 46204 18362 46256 18368
rect 46388 18420 46440 18426
rect 46388 18362 46440 18368
rect 46664 18420 46716 18426
rect 46664 18362 46716 18368
rect 46768 18154 46796 18770
rect 47032 18760 47084 18766
rect 47032 18702 47084 18708
rect 47044 18426 47072 18702
rect 47032 18420 47084 18426
rect 47032 18362 47084 18368
rect 46756 18148 46808 18154
rect 46756 18090 46808 18096
rect 47124 18148 47176 18154
rect 47124 18090 47176 18096
rect 46572 18080 46624 18086
rect 46572 18022 46624 18028
rect 46020 17876 46072 17882
rect 46020 17818 46072 17824
rect 45284 17672 45336 17678
rect 45284 17614 45336 17620
rect 45652 17128 45704 17134
rect 45652 17070 45704 17076
rect 45560 16788 45612 16794
rect 45560 16730 45612 16736
rect 45100 16652 45152 16658
rect 45100 16594 45152 16600
rect 44836 16408 44956 16436
rect 44640 16108 44692 16114
rect 44640 16050 44692 16056
rect 44732 16040 44784 16046
rect 44732 15982 44784 15988
rect 44364 15904 44416 15910
rect 44364 15846 44416 15852
rect 44376 15706 44404 15846
rect 44364 15700 44416 15706
rect 44364 15642 44416 15648
rect 44640 15360 44692 15366
rect 44640 15302 44692 15308
rect 44282 15260 44590 15269
rect 44282 15258 44288 15260
rect 44344 15258 44368 15260
rect 44424 15258 44448 15260
rect 44504 15258 44528 15260
rect 44584 15258 44590 15260
rect 44344 15206 44346 15258
rect 44526 15206 44528 15258
rect 44282 15204 44288 15206
rect 44344 15204 44368 15206
rect 44424 15204 44448 15206
rect 44504 15204 44528 15206
rect 44584 15204 44590 15206
rect 44282 15195 44590 15204
rect 44652 14958 44680 15302
rect 44640 14952 44692 14958
rect 44640 14894 44692 14900
rect 44744 14822 44772 15982
rect 44732 14816 44784 14822
rect 44732 14758 44784 14764
rect 44640 14272 44692 14278
rect 44640 14214 44692 14220
rect 44282 14172 44590 14181
rect 44282 14170 44288 14172
rect 44344 14170 44368 14172
rect 44424 14170 44448 14172
rect 44504 14170 44528 14172
rect 44584 14170 44590 14172
rect 44344 14118 44346 14170
rect 44526 14118 44528 14170
rect 44282 14116 44288 14118
rect 44344 14116 44368 14118
rect 44424 14116 44448 14118
rect 44504 14116 44528 14118
rect 44584 14116 44590 14118
rect 44282 14107 44590 14116
rect 44272 13864 44324 13870
rect 44272 13806 44324 13812
rect 44284 13530 44312 13806
rect 44272 13524 44324 13530
rect 44272 13466 44324 13472
rect 44282 13084 44590 13093
rect 44282 13082 44288 13084
rect 44344 13082 44368 13084
rect 44424 13082 44448 13084
rect 44504 13082 44528 13084
rect 44584 13082 44590 13084
rect 44344 13030 44346 13082
rect 44526 13030 44528 13082
rect 44282 13028 44288 13030
rect 44344 13028 44368 13030
rect 44424 13028 44448 13030
rect 44504 13028 44528 13030
rect 44584 13028 44590 13030
rect 44282 13019 44590 13028
rect 44652 12170 44680 14214
rect 44836 13190 44864 16408
rect 45112 15910 45140 16594
rect 45376 16448 45428 16454
rect 45376 16390 45428 16396
rect 45100 15904 45152 15910
rect 45100 15846 45152 15852
rect 44916 14408 44968 14414
rect 44916 14350 44968 14356
rect 44928 13734 44956 14350
rect 44916 13728 44968 13734
rect 44916 13670 44968 13676
rect 44824 13184 44876 13190
rect 44824 13126 44876 13132
rect 44836 12782 44864 13126
rect 44928 12782 44956 13670
rect 44824 12776 44876 12782
rect 44824 12718 44876 12724
rect 44916 12776 44968 12782
rect 44916 12718 44968 12724
rect 44732 12640 44784 12646
rect 44732 12582 44784 12588
rect 44640 12164 44692 12170
rect 44640 12106 44692 12112
rect 44282 11996 44590 12005
rect 44282 11994 44288 11996
rect 44344 11994 44368 11996
rect 44424 11994 44448 11996
rect 44504 11994 44528 11996
rect 44584 11994 44590 11996
rect 44344 11942 44346 11994
rect 44526 11942 44528 11994
rect 44282 11940 44288 11942
rect 44344 11940 44368 11942
rect 44424 11940 44448 11942
rect 44504 11940 44528 11942
rect 44584 11940 44590 11942
rect 44282 11931 44590 11940
rect 44180 11824 44232 11830
rect 44180 11766 44232 11772
rect 44192 11354 44220 11766
rect 44652 11626 44680 12106
rect 44640 11620 44692 11626
rect 44640 11562 44692 11568
rect 44180 11348 44232 11354
rect 44180 11290 44232 11296
rect 43824 11206 44128 11234
rect 43720 10736 43772 10742
rect 43720 10678 43772 10684
rect 43444 10124 43496 10130
rect 43444 10066 43496 10072
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 40868 8288 40920 8294
rect 40868 8230 40920 8236
rect 40880 7818 40908 8230
rect 40868 7812 40920 7818
rect 40868 7754 40920 7760
rect 41432 7546 41460 8366
rect 41512 8356 41564 8362
rect 41512 8298 41564 8304
rect 41524 7546 41552 8298
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 41512 7540 41564 7546
rect 41512 7482 41564 7488
rect 41420 7404 41472 7410
rect 41420 7346 41472 7352
rect 41432 7002 41460 7346
rect 41420 6996 41472 7002
rect 41420 6938 41472 6944
rect 41236 6656 41288 6662
rect 41236 6598 41288 6604
rect 41248 6458 41276 6598
rect 41236 6452 41288 6458
rect 41236 6394 41288 6400
rect 40868 6248 40920 6254
rect 40868 6190 40920 6196
rect 40776 5704 40828 5710
rect 40776 5646 40828 5652
rect 40500 5364 40552 5370
rect 40500 5306 40552 5312
rect 40880 5098 40908 6190
rect 41144 6112 41196 6118
rect 41144 6054 41196 6060
rect 41156 5914 41184 6054
rect 41144 5908 41196 5914
rect 41144 5850 41196 5856
rect 41156 5574 41184 5850
rect 41144 5568 41196 5574
rect 41144 5510 41196 5516
rect 41236 5228 41288 5234
rect 41236 5170 41288 5176
rect 41052 5160 41104 5166
rect 41052 5102 41104 5108
rect 40868 5092 40920 5098
rect 40868 5034 40920 5040
rect 40500 5024 40552 5030
rect 40500 4966 40552 4972
rect 40408 4616 40460 4622
rect 40408 4558 40460 4564
rect 40420 4282 40448 4558
rect 40512 4282 40540 4966
rect 41064 4758 41092 5102
rect 41248 4758 41276 5170
rect 41328 5024 41380 5030
rect 41328 4966 41380 4972
rect 41052 4752 41104 4758
rect 41052 4694 41104 4700
rect 41236 4752 41288 4758
rect 41236 4694 41288 4700
rect 41340 4690 41368 4966
rect 41328 4684 41380 4690
rect 41328 4626 41380 4632
rect 40592 4548 40644 4554
rect 40592 4490 40644 4496
rect 40408 4276 40460 4282
rect 40408 4218 40460 4224
rect 40500 4276 40552 4282
rect 40500 4218 40552 4224
rect 40316 3936 40368 3942
rect 40316 3878 40368 3884
rect 39948 3596 40000 3602
rect 39948 3538 40000 3544
rect 40132 3596 40184 3602
rect 40132 3538 40184 3544
rect 39856 3392 39908 3398
rect 39856 3334 39908 3340
rect 39868 2446 39896 3334
rect 40132 2916 40184 2922
rect 40132 2858 40184 2864
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39684 2106 39712 2382
rect 39672 2100 39724 2106
rect 39672 2042 39724 2048
rect 40144 800 40172 2858
rect 40408 2848 40460 2854
rect 40408 2790 40460 2796
rect 40420 2446 40448 2790
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 40604 2378 40632 4490
rect 41236 4208 41288 4214
rect 41236 4150 41288 4156
rect 41052 4072 41104 4078
rect 41050 4040 41052 4049
rect 41104 4040 41106 4049
rect 41050 3975 41106 3984
rect 41248 3942 41276 4150
rect 41616 4146 41644 9574
rect 42800 9580 42852 9586
rect 42800 9522 42852 9528
rect 42892 9580 42944 9586
rect 42892 9522 42944 9528
rect 43352 9580 43404 9586
rect 43352 9522 43404 9528
rect 42340 9376 42392 9382
rect 42340 9318 42392 9324
rect 42352 8838 42380 9318
rect 42812 9178 42840 9522
rect 43364 9178 43392 9522
rect 42800 9172 42852 9178
rect 42800 9114 42852 9120
rect 43352 9172 43404 9178
rect 43352 9114 43404 9120
rect 43456 9042 43484 10066
rect 43628 10056 43680 10062
rect 43628 9998 43680 10004
rect 43536 9716 43588 9722
rect 43536 9658 43588 9664
rect 43444 9036 43496 9042
rect 43444 8978 43496 8984
rect 42340 8832 42392 8838
rect 42340 8774 42392 8780
rect 42248 8424 42300 8430
rect 42248 8366 42300 8372
rect 42156 8288 42208 8294
rect 42156 8230 42208 8236
rect 41696 8084 41748 8090
rect 41696 8026 41748 8032
rect 41708 7342 41736 8026
rect 42168 7886 42196 8230
rect 41972 7880 42024 7886
rect 41972 7822 42024 7828
rect 42156 7880 42208 7886
rect 42156 7822 42208 7828
rect 41984 7478 42012 7822
rect 42260 7546 42288 8366
rect 42352 8294 42380 8774
rect 43548 8498 43576 9658
rect 43640 9654 43668 9998
rect 43628 9648 43680 9654
rect 43628 9590 43680 9596
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 42340 8288 42392 8294
rect 42340 8230 42392 8236
rect 42536 8090 42564 8366
rect 42524 8084 42576 8090
rect 42524 8026 42576 8032
rect 42248 7540 42300 7546
rect 42248 7482 42300 7488
rect 41972 7472 42024 7478
rect 41972 7414 42024 7420
rect 41696 7336 41748 7342
rect 41696 7278 41748 7284
rect 42536 6866 42564 8026
rect 43260 7744 43312 7750
rect 43260 7686 43312 7692
rect 42708 7404 42760 7410
rect 42708 7346 42760 7352
rect 42720 7002 42748 7346
rect 43272 7290 43300 7686
rect 43548 7546 43576 8434
rect 43536 7540 43588 7546
rect 43536 7482 43588 7488
rect 43444 7336 43496 7342
rect 43272 7284 43444 7290
rect 43272 7278 43496 7284
rect 43272 7262 43484 7278
rect 42708 6996 42760 7002
rect 42708 6938 42760 6944
rect 42524 6860 42576 6866
rect 42524 6802 42576 6808
rect 42616 6860 42668 6866
rect 42616 6802 42668 6808
rect 42064 6792 42116 6798
rect 42064 6734 42116 6740
rect 42076 6458 42104 6734
rect 42064 6452 42116 6458
rect 42064 6394 42116 6400
rect 41696 6248 41748 6254
rect 41696 6190 41748 6196
rect 41708 5914 41736 6190
rect 41696 5908 41748 5914
rect 41696 5850 41748 5856
rect 42076 5846 42104 6394
rect 41880 5840 41932 5846
rect 41880 5782 41932 5788
rect 42064 5840 42116 5846
rect 42064 5782 42116 5788
rect 41788 5568 41840 5574
rect 41788 5510 41840 5516
rect 41800 5370 41828 5510
rect 41788 5364 41840 5370
rect 41788 5306 41840 5312
rect 41892 5250 41920 5782
rect 42156 5568 42208 5574
rect 42156 5510 42208 5516
rect 41800 5222 41920 5250
rect 41800 4622 41828 5222
rect 42168 5030 42196 5510
rect 42628 5234 42656 6802
rect 42720 5574 42748 6938
rect 43272 6866 43300 7262
rect 43260 6860 43312 6866
rect 43260 6802 43312 6808
rect 43076 6792 43128 6798
rect 43076 6734 43128 6740
rect 42800 6656 42852 6662
rect 42800 6598 42852 6604
rect 42708 5568 42760 5574
rect 42708 5510 42760 5516
rect 42812 5302 42840 6598
rect 43088 6458 43116 6734
rect 43628 6656 43680 6662
rect 43628 6598 43680 6604
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 43640 6390 43668 6598
rect 43628 6384 43680 6390
rect 43628 6326 43680 6332
rect 43352 6112 43404 6118
rect 43352 6054 43404 6060
rect 43364 5710 43392 6054
rect 43640 5914 43668 6326
rect 43628 5908 43680 5914
rect 43628 5850 43680 5856
rect 43824 5794 43852 11206
rect 44282 10908 44590 10917
rect 44282 10906 44288 10908
rect 44344 10906 44368 10908
rect 44424 10906 44448 10908
rect 44504 10906 44528 10908
rect 44584 10906 44590 10908
rect 44344 10854 44346 10906
rect 44526 10854 44528 10906
rect 44282 10852 44288 10854
rect 44344 10852 44368 10854
rect 44424 10852 44448 10854
rect 44504 10852 44528 10854
rect 44584 10852 44590 10854
rect 44282 10843 44590 10852
rect 44456 10668 44508 10674
rect 44456 10610 44508 10616
rect 43904 10464 43956 10470
rect 43904 10406 43956 10412
rect 43916 10130 43944 10406
rect 44468 10266 44496 10610
rect 44456 10260 44508 10266
rect 44456 10202 44508 10208
rect 43904 10124 43956 10130
rect 43904 10066 43956 10072
rect 44180 10124 44232 10130
rect 44180 10066 44232 10072
rect 44192 9654 44220 10066
rect 44640 10056 44692 10062
rect 44640 9998 44692 10004
rect 44282 9820 44590 9829
rect 44282 9818 44288 9820
rect 44344 9818 44368 9820
rect 44424 9818 44448 9820
rect 44504 9818 44528 9820
rect 44584 9818 44590 9820
rect 44344 9766 44346 9818
rect 44526 9766 44528 9818
rect 44282 9764 44288 9766
rect 44344 9764 44368 9766
rect 44424 9764 44448 9766
rect 44504 9764 44528 9766
rect 44584 9764 44590 9766
rect 44282 9755 44590 9764
rect 44180 9648 44232 9654
rect 44180 9590 44232 9596
rect 44364 9648 44416 9654
rect 44364 9590 44416 9596
rect 44180 9512 44232 9518
rect 44180 9454 44232 9460
rect 44192 7750 44220 9454
rect 44376 9178 44404 9590
rect 44364 9172 44416 9178
rect 44364 9114 44416 9120
rect 44282 8732 44590 8741
rect 44282 8730 44288 8732
rect 44344 8730 44368 8732
rect 44424 8730 44448 8732
rect 44504 8730 44528 8732
rect 44584 8730 44590 8732
rect 44344 8678 44346 8730
rect 44526 8678 44528 8730
rect 44282 8676 44288 8678
rect 44344 8676 44368 8678
rect 44424 8676 44448 8678
rect 44504 8676 44528 8678
rect 44584 8676 44590 8678
rect 44282 8667 44590 8676
rect 44652 8634 44680 9998
rect 44744 9654 44772 12582
rect 44836 9994 44864 12718
rect 45112 11914 45140 15846
rect 45388 15502 45416 16390
rect 45572 15502 45600 16730
rect 45664 16590 45692 17070
rect 45652 16584 45704 16590
rect 45652 16526 45704 16532
rect 45744 16516 45796 16522
rect 45744 16458 45796 16464
rect 45376 15496 45428 15502
rect 45376 15438 45428 15444
rect 45560 15496 45612 15502
rect 45560 15438 45612 15444
rect 45284 13864 45336 13870
rect 45284 13806 45336 13812
rect 45192 13184 45244 13190
rect 45192 13126 45244 13132
rect 45204 12238 45232 13126
rect 45192 12232 45244 12238
rect 45192 12174 45244 12180
rect 45112 11886 45232 11914
rect 45100 11688 45152 11694
rect 45100 11630 45152 11636
rect 45112 11354 45140 11630
rect 45100 11348 45152 11354
rect 45100 11290 45152 11296
rect 44916 11144 44968 11150
rect 44916 11086 44968 11092
rect 44928 10606 44956 11086
rect 44916 10600 44968 10606
rect 44916 10542 44968 10548
rect 44824 9988 44876 9994
rect 44824 9930 44876 9936
rect 44732 9648 44784 9654
rect 44732 9590 44784 9596
rect 44836 9586 44864 9930
rect 44824 9580 44876 9586
rect 44824 9522 44876 9528
rect 44836 9042 44864 9522
rect 45008 9512 45060 9518
rect 45008 9454 45060 9460
rect 44824 9036 44876 9042
rect 44824 8978 44876 8984
rect 44732 8900 44784 8906
rect 44732 8842 44784 8848
rect 44640 8628 44692 8634
rect 44640 8570 44692 8576
rect 44652 7954 44680 8570
rect 44640 7948 44692 7954
rect 44640 7890 44692 7896
rect 43996 7744 44048 7750
rect 43996 7686 44048 7692
rect 44180 7744 44232 7750
rect 44180 7686 44232 7692
rect 44008 7478 44036 7686
rect 44282 7644 44590 7653
rect 44282 7642 44288 7644
rect 44344 7642 44368 7644
rect 44424 7642 44448 7644
rect 44504 7642 44528 7644
rect 44584 7642 44590 7644
rect 44344 7590 44346 7642
rect 44526 7590 44528 7642
rect 44282 7588 44288 7590
rect 44344 7588 44368 7590
rect 44424 7588 44448 7590
rect 44504 7588 44528 7590
rect 44584 7588 44590 7590
rect 44282 7579 44590 7588
rect 43996 7472 44048 7478
rect 44088 7472 44140 7478
rect 43996 7414 44048 7420
rect 44086 7440 44088 7449
rect 44140 7440 44142 7449
rect 44008 6934 44036 7414
rect 44086 7375 44142 7384
rect 43996 6928 44048 6934
rect 43996 6870 44048 6876
rect 44282 6556 44590 6565
rect 44282 6554 44288 6556
rect 44344 6554 44368 6556
rect 44424 6554 44448 6556
rect 44504 6554 44528 6556
rect 44584 6554 44590 6556
rect 44344 6502 44346 6554
rect 44526 6502 44528 6554
rect 44282 6500 44288 6502
rect 44344 6500 44368 6502
rect 44424 6500 44448 6502
rect 44504 6500 44528 6502
rect 44584 6500 44590 6502
rect 44282 6491 44590 6500
rect 44088 6384 44140 6390
rect 44088 6326 44140 6332
rect 43824 5766 43944 5794
rect 43352 5704 43404 5710
rect 43352 5646 43404 5652
rect 42800 5296 42852 5302
rect 42800 5238 42852 5244
rect 42616 5228 42668 5234
rect 42616 5170 42668 5176
rect 42708 5160 42760 5166
rect 42708 5102 42760 5108
rect 42156 5024 42208 5030
rect 42156 4966 42208 4972
rect 41880 4820 41932 4826
rect 41880 4762 41932 4768
rect 41788 4616 41840 4622
rect 41788 4558 41840 4564
rect 41604 4140 41656 4146
rect 41604 4082 41656 4088
rect 41236 3936 41288 3942
rect 41236 3878 41288 3884
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 40696 3194 40724 3334
rect 41616 3194 41644 3878
rect 41788 3460 41840 3466
rect 41788 3402 41840 3408
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 41604 3188 41656 3194
rect 41604 3130 41656 3136
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40696 800 40724 2926
rect 41328 2508 41380 2514
rect 41248 2468 41328 2496
rect 41248 800 41276 2468
rect 41328 2450 41380 2456
rect 41800 800 41828 3402
rect 41892 3194 41920 4762
rect 41972 4684 42024 4690
rect 41972 4626 42024 4632
rect 41984 3534 42012 4626
rect 42168 4078 42196 4966
rect 42720 4826 42748 5102
rect 43536 5024 43588 5030
rect 43536 4966 43588 4972
rect 42708 4820 42760 4826
rect 42708 4762 42760 4768
rect 42616 4616 42668 4622
rect 42616 4558 42668 4564
rect 42890 4584 42946 4593
rect 42628 4078 42656 4558
rect 42890 4519 42946 4528
rect 42156 4072 42208 4078
rect 42076 4032 42156 4060
rect 42076 3670 42104 4032
rect 42156 4014 42208 4020
rect 42616 4072 42668 4078
rect 42616 4014 42668 4020
rect 42248 3936 42300 3942
rect 42248 3878 42300 3884
rect 42156 3732 42208 3738
rect 42156 3674 42208 3680
rect 42064 3664 42116 3670
rect 42064 3606 42116 3612
rect 41972 3528 42024 3534
rect 41972 3470 42024 3476
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41984 2854 42012 3470
rect 41972 2848 42024 2854
rect 41972 2790 42024 2796
rect 42168 2774 42196 3674
rect 42260 2922 42288 3878
rect 42904 3738 42932 4519
rect 42984 4208 43036 4214
rect 42984 4150 43036 4156
rect 42996 3738 43024 4150
rect 42892 3732 42944 3738
rect 42892 3674 42944 3680
rect 42984 3732 43036 3738
rect 42984 3674 43036 3680
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 42892 3460 42944 3466
rect 42892 3402 42944 3408
rect 42904 2961 42932 3402
rect 43088 3194 43116 3538
rect 43168 3392 43220 3398
rect 43168 3334 43220 3340
rect 43076 3188 43128 3194
rect 43076 3130 43128 3136
rect 42890 2952 42946 2961
rect 42248 2916 42300 2922
rect 42890 2887 42946 2896
rect 42248 2858 42300 2864
rect 42168 2746 42288 2774
rect 42260 2446 42288 2746
rect 42248 2440 42300 2446
rect 42248 2382 42300 2388
rect 42352 2378 42564 2394
rect 42352 2372 42576 2378
rect 42352 2366 42524 2372
rect 42352 800 42380 2366
rect 42524 2314 42576 2320
rect 42904 870 43024 898
rect 42904 800 42932 870
rect 37476 734 37688 762
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 42996 762 43024 870
rect 43180 762 43208 3334
rect 43548 3194 43576 4966
rect 43812 4480 43864 4486
rect 43812 4422 43864 4428
rect 43824 4146 43852 4422
rect 43812 4140 43864 4146
rect 43812 4082 43864 4088
rect 43916 3534 43944 5766
rect 44100 4622 44128 6326
rect 44178 5672 44234 5681
rect 44178 5607 44180 5616
rect 44232 5607 44234 5616
rect 44180 5578 44232 5584
rect 44282 5468 44590 5477
rect 44282 5466 44288 5468
rect 44344 5466 44368 5468
rect 44424 5466 44448 5468
rect 44504 5466 44528 5468
rect 44584 5466 44590 5468
rect 44344 5414 44346 5466
rect 44526 5414 44528 5466
rect 44282 5412 44288 5414
rect 44344 5412 44368 5414
rect 44424 5412 44448 5414
rect 44504 5412 44528 5414
rect 44584 5412 44590 5414
rect 44282 5403 44590 5412
rect 44180 5364 44232 5370
rect 44180 5306 44232 5312
rect 44192 4690 44220 5306
rect 44180 4684 44232 4690
rect 44180 4626 44232 4632
rect 44088 4616 44140 4622
rect 44088 4558 44140 4564
rect 44192 4282 44220 4626
rect 44640 4616 44692 4622
rect 44640 4558 44692 4564
rect 44282 4380 44590 4389
rect 44282 4378 44288 4380
rect 44344 4378 44368 4380
rect 44424 4378 44448 4380
rect 44504 4378 44528 4380
rect 44584 4378 44590 4380
rect 44344 4326 44346 4378
rect 44526 4326 44528 4378
rect 44282 4324 44288 4326
rect 44344 4324 44368 4326
rect 44424 4324 44448 4326
rect 44504 4324 44528 4326
rect 44584 4324 44590 4326
rect 44282 4315 44590 4324
rect 44180 4276 44232 4282
rect 44180 4218 44232 4224
rect 44272 4276 44324 4282
rect 44652 4264 44680 4558
rect 44272 4218 44324 4224
rect 44560 4236 44680 4264
rect 44284 4146 44312 4218
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 43996 3528 44048 3534
rect 44192 3482 44220 3538
rect 44284 3482 44312 4082
rect 44560 4026 44588 4236
rect 44640 4140 44692 4146
rect 44640 4082 44692 4088
rect 44468 4010 44588 4026
rect 44456 4004 44588 4010
rect 44508 3998 44588 4004
rect 44456 3946 44508 3952
rect 43996 3470 44048 3476
rect 43812 3460 43864 3466
rect 43812 3402 43864 3408
rect 43536 3188 43588 3194
rect 43536 3130 43588 3136
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43364 2650 43392 2994
rect 43720 2848 43772 2854
rect 43720 2790 43772 2796
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 43732 2446 43760 2790
rect 43720 2440 43772 2446
rect 43720 2382 43772 2388
rect 43444 2372 43496 2378
rect 43444 2314 43496 2320
rect 43456 800 43484 2314
rect 43824 2310 43852 3402
rect 44008 3058 44036 3470
rect 44100 3454 44312 3482
rect 44100 3058 44128 3454
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44192 3108 44220 3334
rect 44282 3292 44590 3301
rect 44282 3290 44288 3292
rect 44344 3290 44368 3292
rect 44424 3290 44448 3292
rect 44504 3290 44528 3292
rect 44584 3290 44590 3292
rect 44344 3238 44346 3290
rect 44526 3238 44528 3290
rect 44282 3236 44288 3238
rect 44344 3236 44368 3238
rect 44424 3236 44448 3238
rect 44504 3236 44528 3238
rect 44584 3236 44590 3238
rect 44282 3227 44590 3236
rect 44192 3080 44312 3108
rect 43996 3052 44048 3058
rect 43996 2994 44048 3000
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 43996 2848 44048 2854
rect 43996 2790 44048 2796
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 44008 800 44036 2790
rect 44284 2446 44312 3080
rect 44652 3058 44680 4082
rect 44744 3194 44772 8842
rect 45020 8838 45048 9454
rect 45100 9376 45152 9382
rect 45100 9318 45152 9324
rect 45008 8832 45060 8838
rect 45008 8774 45060 8780
rect 44824 8016 44876 8022
rect 44824 7958 44876 7964
rect 44836 7206 44864 7958
rect 44916 7268 44968 7274
rect 44916 7210 44968 7216
rect 44824 7200 44876 7206
rect 44822 7168 44824 7177
rect 44876 7168 44878 7177
rect 44822 7103 44878 7112
rect 44836 6662 44864 7103
rect 44928 7041 44956 7210
rect 44914 7032 44970 7041
rect 44914 6967 44970 6976
rect 44824 6656 44876 6662
rect 44824 6598 44876 6604
rect 44836 6390 44864 6598
rect 44824 6384 44876 6390
rect 44824 6326 44876 6332
rect 44824 6112 44876 6118
rect 44824 6054 44876 6060
rect 44836 5574 44864 6054
rect 44824 5568 44876 5574
rect 44824 5510 44876 5516
rect 44836 4690 44864 5510
rect 45020 5098 45048 8774
rect 45008 5092 45060 5098
rect 45008 5034 45060 5040
rect 44824 4684 44876 4690
rect 44824 4626 44876 4632
rect 44836 4282 44864 4626
rect 44916 4616 44968 4622
rect 44916 4558 44968 4564
rect 44824 4276 44876 4282
rect 44824 4218 44876 4224
rect 44824 3392 44876 3398
rect 44824 3334 44876 3340
rect 44732 3188 44784 3194
rect 44732 3130 44784 3136
rect 44836 3126 44864 3334
rect 44824 3120 44876 3126
rect 44824 3062 44876 3068
rect 44456 3052 44508 3058
rect 44456 2994 44508 3000
rect 44640 3052 44692 3058
rect 44640 2994 44692 3000
rect 44468 2650 44496 2994
rect 44456 2644 44508 2650
rect 44456 2586 44508 2592
rect 44272 2440 44324 2446
rect 44272 2382 44324 2388
rect 44282 2204 44590 2213
rect 44282 2202 44288 2204
rect 44344 2202 44368 2204
rect 44424 2202 44448 2204
rect 44504 2202 44528 2204
rect 44584 2202 44590 2204
rect 44344 2150 44346 2202
rect 44526 2150 44528 2202
rect 44282 2148 44288 2150
rect 44344 2148 44368 2150
rect 44424 2148 44448 2150
rect 44504 2148 44528 2150
rect 44584 2148 44590 2150
rect 44282 2139 44590 2148
rect 44560 870 44680 898
rect 44560 800 44588 870
rect 42996 734 43208 762
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 44652 762 44680 870
rect 44928 762 44956 4558
rect 45008 4480 45060 4486
rect 45008 4422 45060 4428
rect 45020 3602 45048 4422
rect 45112 4128 45140 9318
rect 45204 8022 45232 11886
rect 45296 8276 45324 13806
rect 45388 9178 45416 15438
rect 45572 15162 45600 15438
rect 45756 15434 45784 16458
rect 46296 15496 46348 15502
rect 46296 15438 46348 15444
rect 45744 15428 45796 15434
rect 45744 15370 45796 15376
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 45560 15156 45612 15162
rect 45560 15098 45612 15104
rect 45560 13320 45612 13326
rect 45560 13262 45612 13268
rect 45744 13320 45796 13326
rect 45744 13262 45796 13268
rect 45468 12640 45520 12646
rect 45468 12582 45520 12588
rect 45480 12306 45508 12582
rect 45468 12300 45520 12306
rect 45468 12242 45520 12248
rect 45572 12238 45600 13262
rect 45756 12986 45784 13262
rect 45744 12980 45796 12986
rect 45744 12922 45796 12928
rect 45560 12232 45612 12238
rect 45560 12174 45612 12180
rect 45652 11688 45704 11694
rect 45652 11630 45704 11636
rect 45664 10810 45692 11630
rect 45836 11212 45888 11218
rect 45836 11154 45888 11160
rect 45744 11008 45796 11014
rect 45744 10950 45796 10956
rect 45652 10804 45704 10810
rect 45652 10746 45704 10752
rect 45664 10130 45692 10746
rect 45756 10742 45784 10950
rect 45744 10736 45796 10742
rect 45744 10678 45796 10684
rect 45848 10606 45876 11154
rect 46020 11008 46072 11014
rect 46020 10950 46072 10956
rect 46032 10606 46060 10950
rect 45836 10600 45888 10606
rect 45836 10542 45888 10548
rect 46020 10600 46072 10606
rect 46020 10542 46072 10548
rect 45836 10464 45888 10470
rect 45836 10406 45888 10412
rect 45652 10124 45704 10130
rect 45652 10066 45704 10072
rect 45848 9994 45876 10406
rect 46216 10266 46244 15302
rect 46308 13394 46336 15438
rect 46584 14822 46612 18022
rect 47136 16046 47164 18090
rect 47412 17678 47440 19790
rect 47688 19174 47716 20198
rect 47780 20058 47808 20198
rect 47768 20052 47820 20058
rect 47768 19994 47820 20000
rect 48516 19786 48544 21286
rect 49160 21146 49188 21422
rect 52000 21412 52052 21418
rect 52000 21354 52052 21360
rect 51504 21244 51812 21253
rect 51504 21242 51510 21244
rect 51566 21242 51590 21244
rect 51646 21242 51670 21244
rect 51726 21242 51750 21244
rect 51806 21242 51812 21244
rect 51566 21190 51568 21242
rect 51748 21190 51750 21242
rect 51504 21188 51510 21190
rect 51566 21188 51590 21190
rect 51646 21188 51670 21190
rect 51726 21188 51750 21190
rect 51806 21188 51812 21190
rect 51504 21179 51812 21188
rect 52012 21146 52040 21354
rect 52828 21344 52880 21350
rect 52828 21286 52880 21292
rect 52840 21146 52868 21286
rect 49148 21140 49200 21146
rect 49148 21082 49200 21088
rect 52000 21140 52052 21146
rect 52000 21082 52052 21088
rect 52828 21140 52880 21146
rect 52828 21082 52880 21088
rect 48780 21004 48832 21010
rect 48780 20946 48832 20952
rect 48504 19780 48556 19786
rect 48504 19722 48556 19728
rect 48320 19712 48372 19718
rect 48320 19654 48372 19660
rect 48332 19310 48360 19654
rect 48792 19514 48820 20946
rect 49424 20936 49476 20942
rect 49424 20878 49476 20884
rect 51264 20936 51316 20942
rect 51264 20878 51316 20884
rect 49332 20800 49384 20806
rect 49332 20742 49384 20748
rect 48872 20324 48924 20330
rect 48872 20266 48924 20272
rect 48780 19508 48832 19514
rect 48780 19450 48832 19456
rect 48884 19394 48912 20266
rect 49056 20052 49108 20058
rect 49056 19994 49108 20000
rect 48964 19848 49016 19854
rect 48964 19790 49016 19796
rect 48976 19514 49004 19790
rect 48964 19508 49016 19514
rect 48964 19450 49016 19456
rect 48792 19366 48912 19394
rect 48792 19310 48820 19366
rect 48320 19304 48372 19310
rect 48320 19246 48372 19252
rect 48780 19304 48832 19310
rect 48780 19246 48832 19252
rect 47676 19168 47728 19174
rect 47676 19110 47728 19116
rect 48228 19168 48280 19174
rect 48228 19110 48280 19116
rect 48596 19168 48648 19174
rect 48596 19110 48648 19116
rect 47584 18896 47636 18902
rect 47584 18838 47636 18844
rect 47492 18828 47544 18834
rect 47492 18770 47544 18776
rect 47504 18426 47532 18770
rect 47492 18420 47544 18426
rect 47492 18362 47544 18368
rect 47400 17672 47452 17678
rect 47400 17614 47452 17620
rect 47412 17338 47440 17614
rect 47400 17332 47452 17338
rect 47400 17274 47452 17280
rect 47596 16114 47624 18838
rect 47688 18358 47716 19110
rect 48240 18902 48268 19110
rect 48228 18896 48280 18902
rect 48228 18838 48280 18844
rect 48608 18834 48636 19110
rect 48596 18828 48648 18834
rect 48596 18770 48648 18776
rect 48136 18692 48188 18698
rect 48136 18634 48188 18640
rect 47676 18352 47728 18358
rect 47676 18294 47728 18300
rect 48148 18272 48176 18634
rect 48412 18624 48464 18630
rect 48412 18566 48464 18572
rect 48320 18284 48372 18290
rect 48148 18244 48320 18272
rect 48320 18226 48372 18232
rect 47768 17604 47820 17610
rect 47768 17546 47820 17552
rect 47780 17338 47808 17546
rect 47768 17332 47820 17338
rect 47768 17274 47820 17280
rect 48424 17202 48452 18566
rect 48504 18216 48556 18222
rect 48504 18158 48556 18164
rect 48516 17882 48544 18158
rect 48504 17876 48556 17882
rect 48504 17818 48556 17824
rect 48608 17678 48636 18770
rect 48792 18222 48820 19246
rect 49068 18766 49096 19994
rect 49344 19378 49372 20742
rect 49436 20466 49464 20878
rect 50896 20800 50948 20806
rect 50896 20742 50948 20748
rect 50908 20534 50936 20742
rect 50896 20528 50948 20534
rect 50896 20470 50948 20476
rect 49424 20460 49476 20466
rect 49424 20402 49476 20408
rect 49436 20058 49464 20402
rect 50712 20256 50764 20262
rect 50712 20198 50764 20204
rect 49424 20052 49476 20058
rect 49424 19994 49476 20000
rect 50724 19922 50752 20198
rect 50712 19916 50764 19922
rect 50712 19858 50764 19864
rect 50160 19712 50212 19718
rect 50160 19654 50212 19660
rect 50172 19514 50200 19654
rect 50160 19508 50212 19514
rect 50160 19450 50212 19456
rect 51276 19446 51304 20878
rect 51908 20800 51960 20806
rect 51908 20742 51960 20748
rect 52552 20800 52604 20806
rect 52552 20742 52604 20748
rect 52920 20800 52972 20806
rect 52920 20742 52972 20748
rect 53012 20800 53064 20806
rect 53012 20742 53064 20748
rect 51920 20602 51948 20742
rect 51908 20596 51960 20602
rect 51908 20538 51960 20544
rect 51504 20156 51812 20165
rect 51504 20154 51510 20156
rect 51566 20154 51590 20156
rect 51646 20154 51670 20156
rect 51726 20154 51750 20156
rect 51806 20154 51812 20156
rect 51566 20102 51568 20154
rect 51748 20102 51750 20154
rect 51504 20100 51510 20102
rect 51566 20100 51590 20102
rect 51646 20100 51670 20102
rect 51726 20100 51750 20102
rect 51806 20100 51812 20102
rect 51504 20091 51812 20100
rect 51920 20058 51948 20538
rect 52564 20466 52592 20742
rect 52826 20496 52882 20505
rect 52552 20460 52604 20466
rect 52826 20431 52882 20440
rect 52552 20402 52604 20408
rect 52840 20398 52868 20431
rect 52828 20392 52880 20398
rect 52828 20334 52880 20340
rect 52840 20058 52868 20334
rect 51908 20052 51960 20058
rect 51908 19994 51960 20000
rect 52828 20052 52880 20058
rect 52828 19994 52880 20000
rect 52932 19922 52960 20742
rect 53024 20534 53052 20742
rect 53012 20528 53064 20534
rect 53012 20470 53064 20476
rect 53012 20392 53064 20398
rect 53012 20334 53064 20340
rect 52920 19916 52972 19922
rect 52920 19858 52972 19864
rect 51264 19440 51316 19446
rect 51264 19382 51316 19388
rect 49332 19372 49384 19378
rect 49332 19314 49384 19320
rect 49344 18766 49372 19314
rect 49700 19236 49752 19242
rect 49700 19178 49752 19184
rect 49056 18760 49108 18766
rect 49056 18702 49108 18708
rect 49332 18760 49384 18766
rect 49332 18702 49384 18708
rect 48872 18624 48924 18630
rect 48872 18566 48924 18572
rect 48964 18624 49016 18630
rect 48964 18566 49016 18572
rect 49148 18624 49200 18630
rect 49148 18566 49200 18572
rect 48780 18216 48832 18222
rect 48700 18176 48780 18204
rect 48596 17672 48648 17678
rect 48596 17614 48648 17620
rect 48412 17196 48464 17202
rect 48412 17138 48464 17144
rect 47768 16584 47820 16590
rect 47768 16526 47820 16532
rect 47780 16250 47808 16526
rect 48228 16448 48280 16454
rect 48228 16390 48280 16396
rect 48596 16448 48648 16454
rect 48596 16390 48648 16396
rect 47768 16244 47820 16250
rect 47768 16186 47820 16192
rect 47584 16108 47636 16114
rect 47584 16050 47636 16056
rect 48044 16108 48096 16114
rect 48044 16050 48096 16056
rect 47124 16040 47176 16046
rect 47124 15982 47176 15988
rect 47136 15910 47164 15982
rect 46848 15904 46900 15910
rect 46848 15846 46900 15852
rect 47124 15904 47176 15910
rect 47124 15846 47176 15852
rect 46860 15502 46888 15846
rect 46848 15496 46900 15502
rect 46848 15438 46900 15444
rect 46756 15428 46808 15434
rect 46756 15370 46808 15376
rect 46768 15162 46796 15370
rect 46756 15156 46808 15162
rect 46756 15098 46808 15104
rect 46572 14816 46624 14822
rect 46572 14758 46624 14764
rect 46584 13870 46612 14758
rect 47032 14272 47084 14278
rect 47032 14214 47084 14220
rect 46572 13864 46624 13870
rect 46572 13806 46624 13812
rect 47044 13734 47072 14214
rect 46756 13728 46808 13734
rect 47032 13728 47084 13734
rect 46756 13670 46808 13676
rect 46952 13676 47032 13682
rect 46952 13670 47084 13676
rect 46296 13388 46348 13394
rect 46296 13330 46348 13336
rect 46308 12850 46336 13330
rect 46768 13258 46796 13670
rect 46952 13654 47072 13670
rect 46756 13252 46808 13258
rect 46756 13194 46808 13200
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46848 12844 46900 12850
rect 46848 12786 46900 12792
rect 46860 12442 46888 12786
rect 46848 12436 46900 12442
rect 46848 12378 46900 12384
rect 46952 11898 46980 13654
rect 47032 12776 47084 12782
rect 47032 12718 47084 12724
rect 47044 12442 47072 12718
rect 47032 12436 47084 12442
rect 47032 12378 47084 12384
rect 46940 11892 46992 11898
rect 46940 11834 46992 11840
rect 46952 11218 46980 11834
rect 47136 11558 47164 15846
rect 48056 15434 48084 16050
rect 48240 15502 48268 16390
rect 48608 16250 48636 16390
rect 48596 16244 48648 16250
rect 48596 16186 48648 16192
rect 48412 15904 48464 15910
rect 48412 15846 48464 15852
rect 48228 15496 48280 15502
rect 48228 15438 48280 15444
rect 48044 15428 48096 15434
rect 48044 15370 48096 15376
rect 48056 14958 48084 15370
rect 48424 15162 48452 15846
rect 48412 15156 48464 15162
rect 48412 15098 48464 15104
rect 48700 15094 48728 18176
rect 48780 18158 48832 18164
rect 48780 17536 48832 17542
rect 48780 17478 48832 17484
rect 48792 16658 48820 17478
rect 48884 17338 48912 18566
rect 48976 18426 49004 18566
rect 48964 18420 49016 18426
rect 48964 18362 49016 18368
rect 48872 17332 48924 17338
rect 48872 17274 48924 17280
rect 49160 16674 49188 18566
rect 49344 17542 49372 18702
rect 49424 18216 49476 18222
rect 49424 18158 49476 18164
rect 49436 17882 49464 18158
rect 49424 17876 49476 17882
rect 49424 17818 49476 17824
rect 49332 17536 49384 17542
rect 49332 17478 49384 17484
rect 49436 17202 49464 17818
rect 49424 17196 49476 17202
rect 49424 17138 49476 17144
rect 49712 16794 49740 19178
rect 51356 19168 51408 19174
rect 51356 19110 51408 19116
rect 52184 19168 52236 19174
rect 52184 19110 52236 19116
rect 52552 19168 52604 19174
rect 52552 19110 52604 19116
rect 52920 19168 52972 19174
rect 52920 19110 52972 19116
rect 50344 18760 50396 18766
rect 50344 18702 50396 18708
rect 50356 17882 50384 18702
rect 50988 18624 51040 18630
rect 50988 18566 51040 18572
rect 51000 18426 51028 18566
rect 50988 18420 51040 18426
rect 50988 18362 51040 18368
rect 51172 18216 51224 18222
rect 51172 18158 51224 18164
rect 50712 18080 50764 18086
rect 50712 18022 50764 18028
rect 50344 17876 50396 17882
rect 50344 17818 50396 17824
rect 50724 17746 50752 18022
rect 50712 17740 50764 17746
rect 50712 17682 50764 17688
rect 51184 17678 51212 18158
rect 51172 17672 51224 17678
rect 51172 17614 51224 17620
rect 49884 17536 49936 17542
rect 49884 17478 49936 17484
rect 49700 16788 49752 16794
rect 49700 16730 49752 16736
rect 48780 16652 48832 16658
rect 48780 16594 48832 16600
rect 48976 16646 49188 16674
rect 49424 16652 49476 16658
rect 48688 15088 48740 15094
rect 48688 15030 48740 15036
rect 48044 14952 48096 14958
rect 48044 14894 48096 14900
rect 47952 14340 48004 14346
rect 47952 14282 48004 14288
rect 47964 14074 47992 14282
rect 47952 14068 48004 14074
rect 47952 14010 48004 14016
rect 47400 13864 47452 13870
rect 47400 13806 47452 13812
rect 47952 13864 48004 13870
rect 48056 13852 48084 14894
rect 48004 13824 48084 13852
rect 47952 13806 48004 13812
rect 47412 12986 47440 13806
rect 47964 12986 47992 13806
rect 48412 13728 48464 13734
rect 48412 13670 48464 13676
rect 48424 13258 48452 13670
rect 48596 13320 48648 13326
rect 48596 13262 48648 13268
rect 48412 13252 48464 13258
rect 48412 13194 48464 13200
rect 48608 12986 48636 13262
rect 47400 12980 47452 12986
rect 47400 12922 47452 12928
rect 47952 12980 48004 12986
rect 47952 12922 48004 12928
rect 48596 12980 48648 12986
rect 48596 12922 48648 12928
rect 47400 12776 47452 12782
rect 47400 12718 47452 12724
rect 47216 12640 47268 12646
rect 47216 12582 47268 12588
rect 47228 12306 47256 12582
rect 47216 12300 47268 12306
rect 47216 12242 47268 12248
rect 47412 12238 47440 12718
rect 48504 12640 48556 12646
rect 48504 12582 48556 12588
rect 48516 12442 48544 12582
rect 48608 12442 48636 12922
rect 48504 12436 48556 12442
rect 48504 12378 48556 12384
rect 48596 12436 48648 12442
rect 48976 12434 49004 16646
rect 49424 16594 49476 16600
rect 49148 16584 49200 16590
rect 49148 16526 49200 16532
rect 49056 16040 49108 16046
rect 49056 15982 49108 15988
rect 49068 15910 49096 15982
rect 49056 15904 49108 15910
rect 49056 15846 49108 15852
rect 49068 15366 49096 15846
rect 49160 15706 49188 16526
rect 49148 15700 49200 15706
rect 49148 15642 49200 15648
rect 49056 15360 49108 15366
rect 49056 15302 49108 15308
rect 49436 15026 49464 16594
rect 49516 15904 49568 15910
rect 49516 15846 49568 15852
rect 49528 15026 49556 15846
rect 49608 15700 49660 15706
rect 49608 15642 49660 15648
rect 49620 15042 49648 15642
rect 49712 15502 49740 16730
rect 49700 15496 49752 15502
rect 49700 15438 49752 15444
rect 49620 15026 49740 15042
rect 49424 15020 49476 15026
rect 49424 14962 49476 14968
rect 49516 15020 49568 15026
rect 49620 15020 49752 15026
rect 49620 15014 49700 15020
rect 49516 14962 49568 14968
rect 49700 14962 49752 14968
rect 49436 14550 49464 14962
rect 49424 14544 49476 14550
rect 49424 14486 49476 14492
rect 49148 14408 49200 14414
rect 49148 14350 49200 14356
rect 49160 13530 49188 14350
rect 49148 13524 49200 13530
rect 49148 13466 49200 13472
rect 49240 13252 49292 13258
rect 49240 13194 49292 13200
rect 49252 12782 49280 13194
rect 49332 13184 49384 13190
rect 49332 13126 49384 13132
rect 49344 12986 49372 13126
rect 49332 12980 49384 12986
rect 49332 12922 49384 12928
rect 49436 12850 49464 14486
rect 49516 13524 49568 13530
rect 49516 13466 49568 13472
rect 49528 12850 49556 13466
rect 49700 13320 49752 13326
rect 49700 13262 49752 13268
rect 49712 12850 49740 13262
rect 49424 12844 49476 12850
rect 49424 12786 49476 12792
rect 49516 12844 49568 12850
rect 49516 12786 49568 12792
rect 49700 12844 49752 12850
rect 49700 12786 49752 12792
rect 49240 12776 49292 12782
rect 49240 12718 49292 12724
rect 48596 12378 48648 12384
rect 48884 12406 49004 12434
rect 47400 12232 47452 12238
rect 47400 12174 47452 12180
rect 47124 11552 47176 11558
rect 47124 11494 47176 11500
rect 46940 11212 46992 11218
rect 46940 11154 46992 11160
rect 46204 10260 46256 10266
rect 46204 10202 46256 10208
rect 45836 9988 45888 9994
rect 45836 9930 45888 9936
rect 45468 9920 45520 9926
rect 45468 9862 45520 9868
rect 45480 9722 45508 9862
rect 45468 9716 45520 9722
rect 45468 9658 45520 9664
rect 45848 9382 45876 9930
rect 46756 9580 46808 9586
rect 46756 9522 46808 9528
rect 45836 9376 45888 9382
rect 45836 9318 45888 9324
rect 46204 9376 46256 9382
rect 46204 9318 46256 9324
rect 45376 9172 45428 9178
rect 45376 9114 45428 9120
rect 45848 8838 45876 9318
rect 45376 8832 45428 8838
rect 45376 8774 45428 8780
rect 45836 8832 45888 8838
rect 45836 8774 45888 8780
rect 45388 8566 45416 8774
rect 46216 8634 46244 9318
rect 46664 9104 46716 9110
rect 46664 9046 46716 9052
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 45376 8560 45428 8566
rect 45376 8502 45428 8508
rect 45560 8424 45612 8430
rect 45560 8366 45612 8372
rect 45376 8288 45428 8294
rect 45296 8248 45376 8276
rect 45376 8230 45428 8236
rect 45192 8016 45244 8022
rect 45192 7958 45244 7964
rect 45388 7410 45416 8230
rect 45572 8090 45600 8366
rect 45560 8084 45612 8090
rect 45560 8026 45612 8032
rect 46480 7812 46532 7818
rect 46480 7754 46532 7760
rect 45468 7744 45520 7750
rect 45468 7686 45520 7692
rect 45376 7404 45428 7410
rect 45376 7346 45428 7352
rect 45192 7200 45244 7206
rect 45192 7142 45244 7148
rect 45204 6934 45232 7142
rect 45192 6928 45244 6934
rect 45192 6870 45244 6876
rect 45204 6322 45232 6870
rect 45192 6316 45244 6322
rect 45192 6258 45244 6264
rect 45204 5778 45232 6258
rect 45192 5772 45244 5778
rect 45192 5714 45244 5720
rect 45204 5370 45232 5714
rect 45192 5364 45244 5370
rect 45192 5306 45244 5312
rect 45388 5030 45416 7346
rect 45480 7002 45508 7686
rect 46492 7206 46520 7754
rect 46480 7200 46532 7206
rect 46480 7142 46532 7148
rect 45468 6996 45520 7002
rect 45468 6938 45520 6944
rect 45652 6792 45704 6798
rect 45652 6734 45704 6740
rect 45664 5370 45692 6734
rect 46492 6730 46520 7142
rect 46676 6866 46704 9046
rect 46768 9042 46796 9522
rect 46940 9512 46992 9518
rect 46940 9454 46992 9460
rect 46952 9178 46980 9454
rect 47136 9382 47164 11494
rect 47308 10600 47360 10606
rect 47412 10588 47440 12174
rect 48780 12096 48832 12102
rect 48780 12038 48832 12044
rect 48412 11688 48464 11694
rect 48412 11630 48464 11636
rect 47768 11552 47820 11558
rect 47768 11494 47820 11500
rect 47492 11076 47544 11082
rect 47492 11018 47544 11024
rect 47360 10560 47440 10588
rect 47308 10542 47360 10548
rect 47504 9654 47532 11018
rect 47780 10810 47808 11494
rect 48320 11280 48372 11286
rect 48320 11222 48372 11228
rect 47952 11008 48004 11014
rect 47952 10950 48004 10956
rect 48228 11008 48280 11014
rect 48228 10950 48280 10956
rect 47964 10810 47992 10950
rect 47768 10804 47820 10810
rect 47768 10746 47820 10752
rect 47952 10804 48004 10810
rect 47952 10746 48004 10752
rect 48240 10674 48268 10950
rect 48228 10668 48280 10674
rect 48228 10610 48280 10616
rect 48136 10464 48188 10470
rect 48136 10406 48188 10412
rect 47492 9648 47544 9654
rect 47492 9590 47544 9596
rect 47768 9444 47820 9450
rect 47768 9386 47820 9392
rect 47124 9376 47176 9382
rect 47124 9318 47176 9324
rect 46940 9172 46992 9178
rect 46940 9114 46992 9120
rect 47136 9042 47164 9318
rect 46756 9036 46808 9042
rect 46756 8978 46808 8984
rect 47124 9036 47176 9042
rect 47124 8978 47176 8984
rect 46768 7546 46796 8978
rect 46756 7540 46808 7546
rect 46756 7482 46808 7488
rect 46664 6860 46716 6866
rect 46664 6802 46716 6808
rect 46768 6798 46796 7482
rect 47136 7206 47164 8978
rect 47780 8838 47808 9386
rect 48044 8968 48096 8974
rect 48044 8910 48096 8916
rect 47768 8832 47820 8838
rect 47768 8774 47820 8780
rect 47780 8430 47808 8774
rect 48056 8634 48084 8910
rect 48044 8628 48096 8634
rect 48044 8570 48096 8576
rect 47952 8492 48004 8498
rect 47952 8434 48004 8440
rect 47768 8424 47820 8430
rect 47768 8366 47820 8372
rect 47964 8090 47992 8434
rect 47952 8084 48004 8090
rect 47952 8026 48004 8032
rect 47584 7812 47636 7818
rect 47584 7754 47636 7760
rect 47596 7546 47624 7754
rect 47584 7540 47636 7546
rect 47584 7482 47636 7488
rect 47124 7200 47176 7206
rect 47124 7142 47176 7148
rect 47860 6860 47912 6866
rect 47860 6802 47912 6808
rect 46756 6792 46808 6798
rect 47308 6792 47360 6798
rect 46808 6740 46888 6746
rect 46756 6734 46888 6740
rect 47308 6734 47360 6740
rect 45836 6724 45888 6730
rect 45836 6666 45888 6672
rect 46480 6724 46532 6730
rect 46480 6666 46532 6672
rect 46664 6724 46716 6730
rect 46768 6718 46888 6734
rect 46664 6666 46716 6672
rect 45744 6656 45796 6662
rect 45744 6598 45796 6604
rect 45756 6458 45784 6598
rect 45744 6452 45796 6458
rect 45744 6394 45796 6400
rect 45652 5364 45704 5370
rect 45652 5306 45704 5312
rect 45376 5024 45428 5030
rect 45376 4966 45428 4972
rect 45284 4480 45336 4486
rect 45284 4422 45336 4428
rect 45296 4214 45324 4422
rect 45284 4208 45336 4214
rect 45284 4150 45336 4156
rect 45192 4140 45244 4146
rect 45112 4100 45192 4128
rect 45192 4082 45244 4088
rect 45098 4040 45154 4049
rect 45098 3975 45154 3984
rect 45112 3602 45140 3975
rect 45284 3936 45336 3942
rect 45284 3878 45336 3884
rect 45008 3596 45060 3602
rect 45008 3538 45060 3544
rect 45100 3596 45152 3602
rect 45100 3538 45152 3544
rect 45008 3392 45060 3398
rect 45008 3334 45060 3340
rect 45020 3194 45048 3334
rect 45008 3188 45060 3194
rect 45008 3130 45060 3136
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 45112 800 45140 3062
rect 45296 3058 45324 3878
rect 45388 3602 45416 4966
rect 45744 4072 45796 4078
rect 45744 4014 45796 4020
rect 45756 3738 45784 4014
rect 45848 4010 45876 6666
rect 46204 6112 46256 6118
rect 46204 6054 46256 6060
rect 46572 6112 46624 6118
rect 46572 6054 46624 6060
rect 46020 5636 46072 5642
rect 46020 5578 46072 5584
rect 46032 4826 46060 5578
rect 46216 5166 46244 6054
rect 46584 5370 46612 6054
rect 46572 5364 46624 5370
rect 46572 5306 46624 5312
rect 46204 5160 46256 5166
rect 46204 5102 46256 5108
rect 46204 5024 46256 5030
rect 46204 4966 46256 4972
rect 46480 5024 46532 5030
rect 46480 4966 46532 4972
rect 46020 4820 46072 4826
rect 46020 4762 46072 4768
rect 45928 4616 45980 4622
rect 45928 4558 45980 4564
rect 45940 4282 45968 4558
rect 45928 4276 45980 4282
rect 45928 4218 45980 4224
rect 46216 4146 46244 4966
rect 46492 4826 46520 4966
rect 46480 4820 46532 4826
rect 46480 4762 46532 4768
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 45836 4004 45888 4010
rect 45836 3946 45888 3952
rect 45744 3732 45796 3738
rect 45744 3674 45796 3680
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 46216 3534 46244 4082
rect 46676 4078 46704 6666
rect 46756 4480 46808 4486
rect 46756 4422 46808 4428
rect 46768 4282 46796 4422
rect 46756 4276 46808 4282
rect 46756 4218 46808 4224
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 46860 3602 46888 6718
rect 47124 6248 47176 6254
rect 47124 6190 47176 6196
rect 47136 5778 47164 6190
rect 47124 5772 47176 5778
rect 47124 5714 47176 5720
rect 47320 5710 47348 6734
rect 47492 6656 47544 6662
rect 47492 6598 47544 6604
rect 47308 5704 47360 5710
rect 47308 5646 47360 5652
rect 47504 5302 47532 6598
rect 47676 6112 47728 6118
rect 47676 6054 47728 6060
rect 47492 5296 47544 5302
rect 47492 5238 47544 5244
rect 47504 4706 47532 5238
rect 47688 5166 47716 6054
rect 47872 5846 47900 6802
rect 48044 6656 48096 6662
rect 48044 6598 48096 6604
rect 47860 5840 47912 5846
rect 47860 5782 47912 5788
rect 47768 5772 47820 5778
rect 47768 5714 47820 5720
rect 47780 5234 47808 5714
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 47676 5160 47728 5166
rect 47676 5102 47728 5108
rect 47504 4678 47624 4706
rect 47308 4616 47360 4622
rect 47308 4558 47360 4564
rect 47492 4616 47544 4622
rect 47492 4558 47544 4564
rect 47216 4140 47268 4146
rect 47216 4082 47268 4088
rect 46938 3632 46994 3641
rect 46848 3596 46900 3602
rect 46938 3567 46994 3576
rect 46848 3538 46900 3544
rect 46204 3528 46256 3534
rect 46204 3470 46256 3476
rect 45652 3392 45704 3398
rect 45652 3334 45704 3340
rect 46204 3392 46256 3398
rect 46204 3334 46256 3340
rect 45284 3052 45336 3058
rect 45284 2994 45336 3000
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45572 2514 45600 2790
rect 45664 2650 45692 3334
rect 45836 2984 45888 2990
rect 45836 2926 45888 2932
rect 45652 2644 45704 2650
rect 45652 2586 45704 2592
rect 45560 2508 45612 2514
rect 45560 2450 45612 2456
rect 45848 1578 45876 2926
rect 45664 1550 45876 1578
rect 45664 800 45692 1550
rect 46216 800 46244 3334
rect 46952 3058 46980 3567
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 46940 3052 46992 3058
rect 46940 2994 46992 3000
rect 47044 2854 47072 3470
rect 47228 3194 47256 4082
rect 47320 4010 47348 4558
rect 47308 4004 47360 4010
rect 47308 3946 47360 3952
rect 47320 3602 47348 3946
rect 47308 3596 47360 3602
rect 47308 3538 47360 3544
rect 47504 3398 47532 4558
rect 47596 4078 47624 4678
rect 47872 4298 47900 5782
rect 47952 5568 48004 5574
rect 47952 5510 48004 5516
rect 47780 4270 47900 4298
rect 47964 4282 47992 5510
rect 47952 4276 48004 4282
rect 47584 4072 47636 4078
rect 47584 4014 47636 4020
rect 47780 3670 47808 4270
rect 47952 4218 48004 4224
rect 47860 4072 47912 4078
rect 47860 4014 47912 4020
rect 47872 3738 47900 4014
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47768 3664 47820 3670
rect 47768 3606 47820 3612
rect 47492 3392 47544 3398
rect 47492 3334 47544 3340
rect 47216 3188 47268 3194
rect 47216 3130 47268 3136
rect 48056 2990 48084 6598
rect 48148 6186 48176 10406
rect 48240 8906 48268 10610
rect 48332 10062 48360 11222
rect 48424 10538 48452 11630
rect 48504 11144 48556 11150
rect 48504 11086 48556 11092
rect 48516 10810 48544 11086
rect 48792 11014 48820 12038
rect 48780 11008 48832 11014
rect 48780 10950 48832 10956
rect 48504 10804 48556 10810
rect 48504 10746 48556 10752
rect 48412 10532 48464 10538
rect 48412 10474 48464 10480
rect 48412 10192 48464 10198
rect 48412 10134 48464 10140
rect 48320 10056 48372 10062
rect 48320 9998 48372 10004
rect 48424 9586 48452 10134
rect 48792 9722 48820 10950
rect 48884 10146 48912 12406
rect 49436 12102 49464 12786
rect 49424 12096 49476 12102
rect 49424 12038 49476 12044
rect 49608 11688 49660 11694
rect 49608 11630 49660 11636
rect 49516 11076 49568 11082
rect 49516 11018 49568 11024
rect 49148 11008 49200 11014
rect 49148 10950 49200 10956
rect 49160 10606 49188 10950
rect 49528 10674 49556 11018
rect 49620 10690 49648 11630
rect 49516 10668 49568 10674
rect 49620 10662 49740 10690
rect 49712 10656 49740 10662
rect 49792 10668 49844 10674
rect 49712 10628 49792 10656
rect 49516 10610 49568 10616
rect 49792 10610 49844 10616
rect 49148 10600 49200 10606
rect 49148 10542 49200 10548
rect 49608 10600 49660 10606
rect 49608 10542 49660 10548
rect 49620 10266 49648 10542
rect 49608 10260 49660 10266
rect 49608 10202 49660 10208
rect 48884 10118 49004 10146
rect 48780 9716 48832 9722
rect 48780 9658 48832 9664
rect 48412 9580 48464 9586
rect 48412 9522 48464 9528
rect 48688 9376 48740 9382
rect 48688 9318 48740 9324
rect 48700 9042 48728 9318
rect 48688 9036 48740 9042
rect 48688 8978 48740 8984
rect 48228 8900 48280 8906
rect 48228 8842 48280 8848
rect 48240 8634 48268 8842
rect 48688 8832 48740 8838
rect 48688 8774 48740 8780
rect 48228 8628 48280 8634
rect 48228 8570 48280 8576
rect 48320 8288 48372 8294
rect 48320 8230 48372 8236
rect 48332 7410 48360 8230
rect 48596 7812 48648 7818
rect 48596 7754 48648 7760
rect 48608 7546 48636 7754
rect 48596 7540 48648 7546
rect 48596 7482 48648 7488
rect 48700 7410 48728 8774
rect 48320 7404 48372 7410
rect 48320 7346 48372 7352
rect 48688 7404 48740 7410
rect 48688 7346 48740 7352
rect 48780 7336 48832 7342
rect 48780 7278 48832 7284
rect 48792 6905 48820 7278
rect 48778 6896 48834 6905
rect 48504 6860 48556 6866
rect 48778 6831 48834 6840
rect 48504 6802 48556 6808
rect 48320 6656 48372 6662
rect 48320 6598 48372 6604
rect 48332 6322 48360 6598
rect 48320 6316 48372 6322
rect 48320 6258 48372 6264
rect 48136 6180 48188 6186
rect 48136 6122 48188 6128
rect 48516 6118 48544 6802
rect 48792 6458 48820 6831
rect 48780 6452 48832 6458
rect 48780 6394 48832 6400
rect 48504 6112 48556 6118
rect 48504 6054 48556 6060
rect 48516 4826 48544 6054
rect 48872 5704 48924 5710
rect 48872 5646 48924 5652
rect 48884 5030 48912 5646
rect 48872 5024 48924 5030
rect 48872 4966 48924 4972
rect 48504 4820 48556 4826
rect 48504 4762 48556 4768
rect 48688 4752 48740 4758
rect 48688 4694 48740 4700
rect 48412 4140 48464 4146
rect 48412 4082 48464 4088
rect 48596 4140 48648 4146
rect 48596 4082 48648 4088
rect 48320 3936 48372 3942
rect 48320 3878 48372 3884
rect 48136 3528 48188 3534
rect 48136 3470 48188 3476
rect 48044 2984 48096 2990
rect 48044 2926 48096 2932
rect 47032 2848 47084 2854
rect 47032 2790 47084 2796
rect 47044 2514 47072 2790
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 47308 2372 47360 2378
rect 47308 2314 47360 2320
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46768 800 46796 2246
rect 47320 800 47348 2314
rect 47872 870 47992 898
rect 47872 800 47900 870
rect 44652 734 44956 762
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 47964 762 47992 870
rect 48148 762 48176 3470
rect 48332 3194 48360 3878
rect 48424 3398 48452 4082
rect 48608 3738 48636 4082
rect 48700 3942 48728 4694
rect 48688 3936 48740 3942
rect 48688 3878 48740 3884
rect 48596 3732 48648 3738
rect 48596 3674 48648 3680
rect 48976 3618 49004 10118
rect 49896 10062 49924 17478
rect 50528 16720 50580 16726
rect 50528 16662 50580 16668
rect 49976 16584 50028 16590
rect 49976 16526 50028 16532
rect 49988 15706 50016 16526
rect 50160 16448 50212 16454
rect 50160 16390 50212 16396
rect 50172 16182 50200 16390
rect 50160 16176 50212 16182
rect 50160 16118 50212 16124
rect 49976 15700 50028 15706
rect 49976 15642 50028 15648
rect 50436 15360 50488 15366
rect 50436 15302 50488 15308
rect 49976 14952 50028 14958
rect 49976 14894 50028 14900
rect 49988 12782 50016 14894
rect 50448 14260 50476 15302
rect 50540 14550 50568 16662
rect 50620 15904 50672 15910
rect 50620 15846 50672 15852
rect 50712 15904 50764 15910
rect 50712 15846 50764 15852
rect 50632 15026 50660 15846
rect 50724 15502 50752 15846
rect 50712 15496 50764 15502
rect 50712 15438 50764 15444
rect 50896 15088 50948 15094
rect 50896 15030 50948 15036
rect 50620 15020 50672 15026
rect 50620 14962 50672 14968
rect 50804 14816 50856 14822
rect 50804 14758 50856 14764
rect 50528 14544 50580 14550
rect 50528 14486 50580 14492
rect 50528 14272 50580 14278
rect 50448 14232 50528 14260
rect 50528 14214 50580 14220
rect 50344 13388 50396 13394
rect 50344 13330 50396 13336
rect 49976 12776 50028 12782
rect 49976 12718 50028 12724
rect 49988 11762 50016 12718
rect 49976 11756 50028 11762
rect 49976 11698 50028 11704
rect 49988 10606 50016 11698
rect 50356 11218 50384 13330
rect 50540 13190 50568 14214
rect 50620 14068 50672 14074
rect 50620 14010 50672 14016
rect 50528 13184 50580 13190
rect 50528 13126 50580 13132
rect 50540 12986 50568 13126
rect 50528 12980 50580 12986
rect 50528 12922 50580 12928
rect 50632 12850 50660 14010
rect 50816 13190 50844 14758
rect 50908 14346 50936 15030
rect 50896 14340 50948 14346
rect 50896 14282 50948 14288
rect 50908 14006 50936 14282
rect 50896 14000 50948 14006
rect 50896 13942 50948 13948
rect 51264 13864 51316 13870
rect 51264 13806 51316 13812
rect 51172 13728 51224 13734
rect 51172 13670 51224 13676
rect 51184 13326 51212 13670
rect 51276 13530 51304 13806
rect 51264 13524 51316 13530
rect 51264 13466 51316 13472
rect 51172 13320 51224 13326
rect 51172 13262 51224 13268
rect 50804 13184 50856 13190
rect 50804 13126 50856 13132
rect 51080 12980 51132 12986
rect 51080 12922 51132 12928
rect 50620 12844 50672 12850
rect 50620 12786 50672 12792
rect 50436 12776 50488 12782
rect 50436 12718 50488 12724
rect 50448 12374 50476 12718
rect 50436 12368 50488 12374
rect 50436 12310 50488 12316
rect 50804 11688 50856 11694
rect 50804 11630 50856 11636
rect 50712 11552 50764 11558
rect 50712 11494 50764 11500
rect 50724 11354 50752 11494
rect 50712 11348 50764 11354
rect 50712 11290 50764 11296
rect 50344 11212 50396 11218
rect 50344 11154 50396 11160
rect 50436 11076 50488 11082
rect 50436 11018 50488 11024
rect 49976 10600 50028 10606
rect 49976 10542 50028 10548
rect 49988 10266 50016 10542
rect 50160 10464 50212 10470
rect 50160 10406 50212 10412
rect 49976 10260 50028 10266
rect 49976 10202 50028 10208
rect 49884 10056 49936 10062
rect 49884 9998 49936 10004
rect 49424 9988 49476 9994
rect 49424 9930 49476 9936
rect 49056 9716 49108 9722
rect 49056 9658 49108 9664
rect 49068 8498 49096 9658
rect 49332 8968 49384 8974
rect 49332 8910 49384 8916
rect 49148 8832 49200 8838
rect 49148 8774 49200 8780
rect 49056 8492 49108 8498
rect 49056 8434 49108 8440
rect 49160 7546 49188 8774
rect 49344 8498 49372 8910
rect 49332 8492 49384 8498
rect 49332 8434 49384 8440
rect 49240 8424 49292 8430
rect 49240 8366 49292 8372
rect 49252 7818 49280 8366
rect 49240 7812 49292 7818
rect 49240 7754 49292 7760
rect 49148 7540 49200 7546
rect 49148 7482 49200 7488
rect 49056 6656 49108 6662
rect 49056 6598 49108 6604
rect 49068 3738 49096 6598
rect 49436 4758 49464 9930
rect 49976 9920 50028 9926
rect 49976 9862 50028 9868
rect 49988 9722 50016 9862
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 49792 9376 49844 9382
rect 49792 9318 49844 9324
rect 49608 9104 49660 9110
rect 49608 9046 49660 9052
rect 49620 8430 49648 9046
rect 49804 9042 49832 9318
rect 49792 9036 49844 9042
rect 49792 8978 49844 8984
rect 49608 8424 49660 8430
rect 49608 8366 49660 8372
rect 49804 6662 49832 8978
rect 50172 8566 50200 10406
rect 50448 9674 50476 11018
rect 50816 10810 50844 11630
rect 50804 10804 50856 10810
rect 50804 10746 50856 10752
rect 50528 10464 50580 10470
rect 50528 10406 50580 10412
rect 50540 9926 50568 10406
rect 50528 9920 50580 9926
rect 50528 9862 50580 9868
rect 50356 9646 50476 9674
rect 50356 8906 50384 9646
rect 51092 9178 51120 12922
rect 51368 12782 51396 19110
rect 51504 19068 51812 19077
rect 51504 19066 51510 19068
rect 51566 19066 51590 19068
rect 51646 19066 51670 19068
rect 51726 19066 51750 19068
rect 51806 19066 51812 19068
rect 51566 19014 51568 19066
rect 51748 19014 51750 19066
rect 51504 19012 51510 19014
rect 51566 19012 51590 19014
rect 51646 19012 51670 19014
rect 51726 19012 51750 19014
rect 51806 19012 51812 19014
rect 51504 19003 51812 19012
rect 52196 18698 52224 19110
rect 52184 18692 52236 18698
rect 52184 18634 52236 18640
rect 51908 18624 51960 18630
rect 51908 18566 51960 18572
rect 51504 17980 51812 17989
rect 51504 17978 51510 17980
rect 51566 17978 51590 17980
rect 51646 17978 51670 17980
rect 51726 17978 51750 17980
rect 51806 17978 51812 17980
rect 51566 17926 51568 17978
rect 51748 17926 51750 17978
rect 51504 17924 51510 17926
rect 51566 17924 51590 17926
rect 51646 17924 51670 17926
rect 51726 17924 51750 17926
rect 51806 17924 51812 17926
rect 51504 17915 51812 17924
rect 51920 17610 51948 18566
rect 51908 17604 51960 17610
rect 51908 17546 51960 17552
rect 52000 17536 52052 17542
rect 52000 17478 52052 17484
rect 51504 16892 51812 16901
rect 51504 16890 51510 16892
rect 51566 16890 51590 16892
rect 51646 16890 51670 16892
rect 51726 16890 51750 16892
rect 51806 16890 51812 16892
rect 51566 16838 51568 16890
rect 51748 16838 51750 16890
rect 51504 16836 51510 16838
rect 51566 16836 51590 16838
rect 51646 16836 51670 16838
rect 51726 16836 51750 16838
rect 51806 16836 51812 16838
rect 51504 16827 51812 16836
rect 52012 16250 52040 17478
rect 52000 16244 52052 16250
rect 52000 16186 52052 16192
rect 51504 15804 51812 15813
rect 51504 15802 51510 15804
rect 51566 15802 51590 15804
rect 51646 15802 51670 15804
rect 51726 15802 51750 15804
rect 51806 15802 51812 15804
rect 51566 15750 51568 15802
rect 51748 15750 51750 15802
rect 51504 15748 51510 15750
rect 51566 15748 51590 15750
rect 51646 15748 51670 15750
rect 51726 15748 51750 15750
rect 51806 15748 51812 15750
rect 51504 15739 51812 15748
rect 52000 15020 52052 15026
rect 52000 14962 52052 14968
rect 51504 14716 51812 14725
rect 51504 14714 51510 14716
rect 51566 14714 51590 14716
rect 51646 14714 51670 14716
rect 51726 14714 51750 14716
rect 51806 14714 51812 14716
rect 51566 14662 51568 14714
rect 51748 14662 51750 14714
rect 51504 14660 51510 14662
rect 51566 14660 51590 14662
rect 51646 14660 51670 14662
rect 51726 14660 51750 14662
rect 51806 14660 51812 14662
rect 51504 14651 51812 14660
rect 52012 14618 52040 14962
rect 52092 14816 52144 14822
rect 52092 14758 52144 14764
rect 52000 14612 52052 14618
rect 52000 14554 52052 14560
rect 52104 14482 52132 14758
rect 52092 14476 52144 14482
rect 52092 14418 52144 14424
rect 52196 14362 52224 18634
rect 52564 18426 52592 19110
rect 52736 18624 52788 18630
rect 52736 18566 52788 18572
rect 52828 18624 52880 18630
rect 52828 18566 52880 18572
rect 52552 18420 52604 18426
rect 52552 18362 52604 18368
rect 52564 18290 52592 18362
rect 52552 18284 52604 18290
rect 52552 18226 52604 18232
rect 52748 17882 52776 18566
rect 52840 18426 52868 18566
rect 52932 18426 52960 19110
rect 53024 18698 53052 20334
rect 53392 19990 53420 21422
rect 54484 21344 54536 21350
rect 54484 21286 54536 21292
rect 55956 21344 56008 21350
rect 55956 21286 56008 21292
rect 56048 21344 56100 21350
rect 56048 21286 56100 21292
rect 53840 21004 53892 21010
rect 53840 20946 53892 20952
rect 53472 20936 53524 20942
rect 53472 20878 53524 20884
rect 53484 20330 53512 20878
rect 53748 20800 53800 20806
rect 53748 20742 53800 20748
rect 53760 20534 53788 20742
rect 53748 20528 53800 20534
rect 53748 20470 53800 20476
rect 53852 20398 53880 20946
rect 54496 20398 54524 21286
rect 55968 21010 55996 21286
rect 54668 21004 54720 21010
rect 54668 20946 54720 20952
rect 55956 21004 56008 21010
rect 55956 20946 56008 20952
rect 54680 20466 54708 20946
rect 55036 20800 55088 20806
rect 55036 20742 55088 20748
rect 55588 20800 55640 20806
rect 55588 20742 55640 20748
rect 54668 20460 54720 20466
rect 54668 20402 54720 20408
rect 53840 20392 53892 20398
rect 53840 20334 53892 20340
rect 54484 20392 54536 20398
rect 54484 20334 54536 20340
rect 54760 20392 54812 20398
rect 54760 20334 54812 20340
rect 53472 20324 53524 20330
rect 53472 20266 53524 20272
rect 53380 19984 53432 19990
rect 53380 19926 53432 19932
rect 53392 19718 53420 19926
rect 53380 19712 53432 19718
rect 53380 19654 53432 19660
rect 54300 19712 54352 19718
rect 54300 19654 54352 19660
rect 54312 18970 54340 19654
rect 54300 18964 54352 18970
rect 54300 18906 54352 18912
rect 53656 18760 53708 18766
rect 53656 18702 53708 18708
rect 53012 18692 53064 18698
rect 53012 18634 53064 18640
rect 52828 18420 52880 18426
rect 52828 18362 52880 18368
rect 52920 18420 52972 18426
rect 52920 18362 52972 18368
rect 53024 18358 53052 18634
rect 53668 18426 53696 18702
rect 53656 18420 53708 18426
rect 53656 18362 53708 18368
rect 53012 18352 53064 18358
rect 53012 18294 53064 18300
rect 52828 18216 52880 18222
rect 52828 18158 52880 18164
rect 52736 17876 52788 17882
rect 52736 17818 52788 17824
rect 52552 15904 52604 15910
rect 52552 15846 52604 15852
rect 52104 14334 52224 14362
rect 51504 13628 51812 13637
rect 51504 13626 51510 13628
rect 51566 13626 51590 13628
rect 51646 13626 51670 13628
rect 51726 13626 51750 13628
rect 51806 13626 51812 13628
rect 51566 13574 51568 13626
rect 51748 13574 51750 13626
rect 51504 13572 51510 13574
rect 51566 13572 51590 13574
rect 51646 13572 51670 13574
rect 51726 13572 51750 13574
rect 51806 13572 51812 13574
rect 51504 13563 51812 13572
rect 51540 13388 51592 13394
rect 51540 13330 51592 13336
rect 51552 12986 51580 13330
rect 51540 12980 51592 12986
rect 51540 12922 51592 12928
rect 51356 12776 51408 12782
rect 51356 12718 51408 12724
rect 51368 12434 51396 12718
rect 51504 12540 51812 12549
rect 51504 12538 51510 12540
rect 51566 12538 51590 12540
rect 51646 12538 51670 12540
rect 51726 12538 51750 12540
rect 51806 12538 51812 12540
rect 51566 12486 51568 12538
rect 51748 12486 51750 12538
rect 51504 12484 51510 12486
rect 51566 12484 51590 12486
rect 51646 12484 51670 12486
rect 51726 12484 51750 12486
rect 51806 12484 51812 12486
rect 51504 12475 51812 12484
rect 51276 12406 51396 12434
rect 51276 11558 51304 12406
rect 51540 12300 51592 12306
rect 51540 12242 51592 12248
rect 51552 11898 51580 12242
rect 51540 11892 51592 11898
rect 51540 11834 51592 11840
rect 51264 11552 51316 11558
rect 51264 11494 51316 11500
rect 51172 11280 51224 11286
rect 51172 11222 51224 11228
rect 51184 9586 51212 11222
rect 51276 11218 51304 11494
rect 51504 11452 51812 11461
rect 51504 11450 51510 11452
rect 51566 11450 51590 11452
rect 51646 11450 51670 11452
rect 51726 11450 51750 11452
rect 51806 11450 51812 11452
rect 51566 11398 51568 11450
rect 51748 11398 51750 11450
rect 51504 11396 51510 11398
rect 51566 11396 51590 11398
rect 51646 11396 51670 11398
rect 51726 11396 51750 11398
rect 51806 11396 51812 11398
rect 51504 11387 51812 11396
rect 51264 11212 51316 11218
rect 51264 11154 51316 11160
rect 51172 9580 51224 9586
rect 51172 9522 51224 9528
rect 51172 9444 51224 9450
rect 51172 9386 51224 9392
rect 51080 9172 51132 9178
rect 51080 9114 51132 9120
rect 51184 9058 51212 9386
rect 51276 9110 51304 11154
rect 51356 11144 51408 11150
rect 51356 11086 51408 11092
rect 51368 10266 51396 11086
rect 51504 10364 51812 10373
rect 51504 10362 51510 10364
rect 51566 10362 51590 10364
rect 51646 10362 51670 10364
rect 51726 10362 51750 10364
rect 51806 10362 51812 10364
rect 51566 10310 51568 10362
rect 51748 10310 51750 10362
rect 51504 10308 51510 10310
rect 51566 10308 51590 10310
rect 51646 10308 51670 10310
rect 51726 10308 51750 10310
rect 51806 10308 51812 10310
rect 51504 10299 51812 10308
rect 51356 10260 51408 10266
rect 51356 10202 51408 10208
rect 51816 9988 51868 9994
rect 51816 9930 51868 9936
rect 51828 9722 51856 9930
rect 51816 9716 51868 9722
rect 51816 9658 51868 9664
rect 51504 9276 51812 9285
rect 51504 9274 51510 9276
rect 51566 9274 51590 9276
rect 51646 9274 51670 9276
rect 51726 9274 51750 9276
rect 51806 9274 51812 9276
rect 51566 9222 51568 9274
rect 51748 9222 51750 9274
rect 51504 9220 51510 9222
rect 51566 9220 51590 9222
rect 51646 9220 51670 9222
rect 51726 9220 51750 9222
rect 51806 9220 51812 9222
rect 51504 9211 51812 9220
rect 51092 9030 51212 9058
rect 51264 9104 51316 9110
rect 51264 9046 51316 9052
rect 51092 8974 51120 9030
rect 51080 8968 51132 8974
rect 51080 8910 51132 8916
rect 50344 8900 50396 8906
rect 50344 8842 50396 8848
rect 50160 8560 50212 8566
rect 50160 8502 50212 8508
rect 49884 8424 49936 8430
rect 49884 8366 49936 8372
rect 50252 8424 50304 8430
rect 50252 8366 50304 8372
rect 49896 7750 49924 8366
rect 50160 8356 50212 8362
rect 50160 8298 50212 8304
rect 50172 8022 50200 8298
rect 50264 8090 50292 8366
rect 50252 8084 50304 8090
rect 50252 8026 50304 8032
rect 50160 8016 50212 8022
rect 50160 7958 50212 7964
rect 49884 7744 49936 7750
rect 49884 7686 49936 7692
rect 49896 7410 49924 7686
rect 50264 7410 50292 8026
rect 49884 7404 49936 7410
rect 49884 7346 49936 7352
rect 50252 7404 50304 7410
rect 50252 7346 50304 7352
rect 49896 6730 49924 7346
rect 49884 6724 49936 6730
rect 49884 6666 49936 6672
rect 49792 6656 49844 6662
rect 49792 6598 49844 6604
rect 50252 6656 50304 6662
rect 50252 6598 50304 6604
rect 49608 6316 49660 6322
rect 49608 6258 49660 6264
rect 49620 5574 49648 6258
rect 49792 6112 49844 6118
rect 49712 6072 49792 6100
rect 49712 5710 49740 6072
rect 49792 6054 49844 6060
rect 50264 5778 50292 6598
rect 50252 5772 50304 5778
rect 50252 5714 50304 5720
rect 49700 5704 49752 5710
rect 49700 5646 49752 5652
rect 50160 5704 50212 5710
rect 50160 5646 50212 5652
rect 49608 5568 49660 5574
rect 49608 5510 49660 5516
rect 49424 4752 49476 4758
rect 49424 4694 49476 4700
rect 49620 4486 49648 5510
rect 50172 5234 50200 5646
rect 50160 5228 50212 5234
rect 50160 5170 50212 5176
rect 50172 4826 50200 5170
rect 50356 5166 50384 8842
rect 50896 8832 50948 8838
rect 50896 8774 50948 8780
rect 50908 8634 50936 8774
rect 50896 8628 50948 8634
rect 50896 8570 50948 8576
rect 50804 6656 50856 6662
rect 50804 6598 50856 6604
rect 51092 6610 51120 8910
rect 51172 8900 51224 8906
rect 51172 8842 51224 8848
rect 51184 8634 51212 8842
rect 51172 8628 51224 8634
rect 51172 8570 51224 8576
rect 51276 8480 51304 9046
rect 51356 8900 51408 8906
rect 51356 8842 51408 8848
rect 51184 8452 51304 8480
rect 51184 6730 51212 8452
rect 51264 8356 51316 8362
rect 51264 8298 51316 8304
rect 51172 6724 51224 6730
rect 51172 6666 51224 6672
rect 50436 5704 50488 5710
rect 50436 5646 50488 5652
rect 50448 5302 50476 5646
rect 50436 5296 50488 5302
rect 50436 5238 50488 5244
rect 50344 5160 50396 5166
rect 50344 5102 50396 5108
rect 50160 4820 50212 4826
rect 50160 4762 50212 4768
rect 50816 4758 50844 6598
rect 51092 6582 51212 6610
rect 51080 6248 51132 6254
rect 51080 6190 51132 6196
rect 51092 5914 51120 6190
rect 51080 5908 51132 5914
rect 51080 5850 51132 5856
rect 51080 5568 51132 5574
rect 51080 5510 51132 5516
rect 51092 5370 51120 5510
rect 51080 5364 51132 5370
rect 51080 5306 51132 5312
rect 50896 5228 50948 5234
rect 50948 5188 51028 5216
rect 50896 5170 50948 5176
rect 50804 4752 50856 4758
rect 50804 4694 50856 4700
rect 49700 4616 49752 4622
rect 49700 4558 49752 4564
rect 49608 4480 49660 4486
rect 49608 4422 49660 4428
rect 49620 4146 49648 4422
rect 49712 4282 49740 4558
rect 50528 4480 50580 4486
rect 50528 4422 50580 4428
rect 50804 4480 50856 4486
rect 50804 4422 50856 4428
rect 50896 4480 50948 4486
rect 50896 4422 50948 4428
rect 49700 4276 49752 4282
rect 49700 4218 49752 4224
rect 49884 4276 49936 4282
rect 49884 4218 49936 4224
rect 49792 4208 49844 4214
rect 49792 4150 49844 4156
rect 49608 4140 49660 4146
rect 49608 4082 49660 4088
rect 49700 3936 49752 3942
rect 49700 3878 49752 3884
rect 49056 3732 49108 3738
rect 49056 3674 49108 3680
rect 48872 3596 48924 3602
rect 48976 3590 49648 3618
rect 48872 3538 48924 3544
rect 48412 3392 48464 3398
rect 48412 3334 48464 3340
rect 48320 3188 48372 3194
rect 48320 3130 48372 3136
rect 48884 3058 48912 3538
rect 49424 3460 49476 3466
rect 49424 3402 49476 3408
rect 49436 3194 49464 3402
rect 49424 3188 49476 3194
rect 49424 3130 49476 3136
rect 49620 3058 49648 3590
rect 49712 3398 49740 3878
rect 49700 3392 49752 3398
rect 49700 3334 49752 3340
rect 48872 3052 48924 3058
rect 48872 2994 48924 3000
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48412 2848 48464 2854
rect 48412 2790 48464 2796
rect 48332 2446 48360 2790
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 48424 800 48452 2790
rect 49804 2650 49832 4150
rect 49896 3602 49924 4218
rect 50540 4146 50568 4422
rect 50816 4282 50844 4422
rect 50908 4282 50936 4422
rect 50804 4276 50856 4282
rect 50804 4218 50856 4224
rect 50896 4276 50948 4282
rect 50896 4218 50948 4224
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4140 50580 4146
rect 50528 4082 50580 4088
rect 50356 3602 50384 4082
rect 49884 3596 49936 3602
rect 49884 3538 49936 3544
rect 50344 3596 50396 3602
rect 50344 3538 50396 3544
rect 50252 3460 50304 3466
rect 50252 3402 50304 3408
rect 50264 3210 50292 3402
rect 50080 3182 50292 3210
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 49240 2508 49292 2514
rect 49240 2450 49292 2456
rect 48976 870 49096 898
rect 48976 800 49004 870
rect 47964 734 48176 762
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49068 762 49096 870
rect 49252 762 49280 2450
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49712 1442 49740 2382
rect 49528 1414 49740 1442
rect 49528 800 49556 1414
rect 50080 800 50108 3182
rect 50356 3126 50384 3538
rect 50712 3528 50764 3534
rect 50712 3470 50764 3476
rect 50724 3194 50752 3470
rect 50712 3188 50764 3194
rect 50712 3130 50764 3136
rect 50344 3120 50396 3126
rect 50344 3062 50396 3068
rect 50632 3046 50752 3074
rect 50252 2848 50304 2854
rect 50252 2790 50304 2796
rect 50264 2446 50292 2790
rect 50252 2440 50304 2446
rect 50252 2382 50304 2388
rect 50632 800 50660 3046
rect 50724 2990 50752 3046
rect 50712 2984 50764 2990
rect 50712 2926 50764 2932
rect 51000 2310 51028 5188
rect 51184 5030 51212 6582
rect 51172 5024 51224 5030
rect 51092 4972 51172 4978
rect 51092 4966 51224 4972
rect 51092 4950 51212 4966
rect 51092 4078 51120 4950
rect 51172 4684 51224 4690
rect 51172 4626 51224 4632
rect 51080 4072 51132 4078
rect 51080 4014 51132 4020
rect 51184 2650 51212 4626
rect 51276 4146 51304 8298
rect 51368 4826 51396 8842
rect 52104 8537 52132 14334
rect 52368 13456 52420 13462
rect 52368 13398 52420 13404
rect 52276 13320 52328 13326
rect 52274 13288 52276 13297
rect 52328 13288 52330 13297
rect 52274 13223 52330 13232
rect 52276 12980 52328 12986
rect 52276 12922 52328 12928
rect 52184 12640 52236 12646
rect 52184 12582 52236 12588
rect 52196 12306 52224 12582
rect 52184 12300 52236 12306
rect 52184 12242 52236 12248
rect 52288 11098 52316 12922
rect 52196 11070 52316 11098
rect 52090 8528 52146 8537
rect 52090 8463 52146 8472
rect 51908 8288 51960 8294
rect 51908 8230 51960 8236
rect 51504 8188 51812 8197
rect 51504 8186 51510 8188
rect 51566 8186 51590 8188
rect 51646 8186 51670 8188
rect 51726 8186 51750 8188
rect 51806 8186 51812 8188
rect 51566 8134 51568 8186
rect 51748 8134 51750 8186
rect 51504 8132 51510 8134
rect 51566 8132 51590 8134
rect 51646 8132 51670 8134
rect 51726 8132 51750 8134
rect 51806 8132 51812 8134
rect 51504 8123 51812 8132
rect 51920 7886 51948 8230
rect 51908 7880 51960 7886
rect 51908 7822 51960 7828
rect 52000 7744 52052 7750
rect 52000 7686 52052 7692
rect 52012 7546 52040 7686
rect 52000 7540 52052 7546
rect 52000 7482 52052 7488
rect 52012 7206 52040 7482
rect 52196 7410 52224 11070
rect 52276 11008 52328 11014
rect 52276 10950 52328 10956
rect 52288 10198 52316 10950
rect 52276 10192 52328 10198
rect 52276 10134 52328 10140
rect 52276 9444 52328 9450
rect 52276 9386 52328 9392
rect 52288 9042 52316 9386
rect 52276 9036 52328 9042
rect 52276 8978 52328 8984
rect 52184 7404 52236 7410
rect 52184 7346 52236 7352
rect 52000 7200 52052 7206
rect 52000 7142 52052 7148
rect 51504 7100 51812 7109
rect 51504 7098 51510 7100
rect 51566 7098 51590 7100
rect 51646 7098 51670 7100
rect 51726 7098 51750 7100
rect 51806 7098 51812 7100
rect 51566 7046 51568 7098
rect 51748 7046 51750 7098
rect 51504 7044 51510 7046
rect 51566 7044 51590 7046
rect 51646 7044 51670 7046
rect 51726 7044 51750 7046
rect 51806 7044 51812 7046
rect 51504 7035 51812 7044
rect 51908 6792 51960 6798
rect 51908 6734 51960 6740
rect 51920 6458 51948 6734
rect 52012 6662 52040 7142
rect 52000 6656 52052 6662
rect 52000 6598 52052 6604
rect 52276 6656 52328 6662
rect 52276 6598 52328 6604
rect 51908 6452 51960 6458
rect 51908 6394 51960 6400
rect 51504 6012 51812 6021
rect 51504 6010 51510 6012
rect 51566 6010 51590 6012
rect 51646 6010 51670 6012
rect 51726 6010 51750 6012
rect 51806 6010 51812 6012
rect 51566 5958 51568 6010
rect 51748 5958 51750 6010
rect 51504 5956 51510 5958
rect 51566 5956 51590 5958
rect 51646 5956 51670 5958
rect 51726 5956 51750 5958
rect 51806 5956 51812 5958
rect 51504 5947 51812 5956
rect 52288 5642 52316 6598
rect 52276 5636 52328 5642
rect 52276 5578 52328 5584
rect 51504 4924 51812 4933
rect 51504 4922 51510 4924
rect 51566 4922 51590 4924
rect 51646 4922 51670 4924
rect 51726 4922 51750 4924
rect 51806 4922 51812 4924
rect 51566 4870 51568 4922
rect 51748 4870 51750 4922
rect 51504 4868 51510 4870
rect 51566 4868 51590 4870
rect 51646 4868 51670 4870
rect 51726 4868 51750 4870
rect 51806 4868 51812 4870
rect 51504 4859 51812 4868
rect 51356 4820 51408 4826
rect 51356 4762 51408 4768
rect 51448 4616 51500 4622
rect 51448 4558 51500 4564
rect 52000 4616 52052 4622
rect 52000 4558 52052 4564
rect 52092 4616 52144 4622
rect 52092 4558 52144 4564
rect 51356 4548 51408 4554
rect 51356 4490 51408 4496
rect 51264 4140 51316 4146
rect 51264 4082 51316 4088
rect 51368 3738 51396 4490
rect 51460 4282 51488 4558
rect 51448 4276 51500 4282
rect 51448 4218 51500 4224
rect 51908 3936 51960 3942
rect 51908 3878 51960 3884
rect 51504 3836 51812 3845
rect 51504 3834 51510 3836
rect 51566 3834 51590 3836
rect 51646 3834 51670 3836
rect 51726 3834 51750 3836
rect 51806 3834 51812 3836
rect 51566 3782 51568 3834
rect 51748 3782 51750 3834
rect 51504 3780 51510 3782
rect 51566 3780 51590 3782
rect 51646 3780 51670 3782
rect 51726 3780 51750 3782
rect 51806 3780 51812 3782
rect 51504 3771 51812 3780
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 51920 3534 51948 3878
rect 52012 3738 52040 4558
rect 52000 3732 52052 3738
rect 52000 3674 52052 3680
rect 51908 3528 51960 3534
rect 51908 3470 51960 3476
rect 52000 3528 52052 3534
rect 52000 3470 52052 3476
rect 51724 3392 51776 3398
rect 51776 3340 51948 3346
rect 51724 3334 51948 3340
rect 51736 3318 51948 3334
rect 51504 2748 51812 2757
rect 51504 2746 51510 2748
rect 51566 2746 51590 2748
rect 51646 2746 51670 2748
rect 51726 2746 51750 2748
rect 51806 2746 51812 2748
rect 51566 2694 51568 2746
rect 51748 2694 51750 2746
rect 51504 2692 51510 2694
rect 51566 2692 51590 2694
rect 51646 2692 51670 2694
rect 51726 2692 51750 2694
rect 51806 2692 51812 2694
rect 51504 2683 51812 2692
rect 51920 2650 51948 3318
rect 51172 2644 51224 2650
rect 51172 2586 51224 2592
rect 51908 2644 51960 2650
rect 51908 2586 51960 2592
rect 52012 2514 52040 3470
rect 52000 2508 52052 2514
rect 52000 2450 52052 2456
rect 51356 2372 51408 2378
rect 51356 2314 51408 2320
rect 50988 2304 51040 2310
rect 50988 2246 51040 2252
rect 51368 1306 51396 2314
rect 51184 1278 51396 1306
rect 51184 800 51212 1278
rect 51736 870 51856 898
rect 51736 800 51764 870
rect 49068 734 49280 762
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 51828 762 51856 870
rect 52104 762 52132 4558
rect 52380 3058 52408 13398
rect 52460 13184 52512 13190
rect 52460 13126 52512 13132
rect 52472 12782 52500 13126
rect 52460 12776 52512 12782
rect 52460 12718 52512 12724
rect 52472 12442 52500 12718
rect 52460 12436 52512 12442
rect 52460 12378 52512 12384
rect 52460 10668 52512 10674
rect 52460 10610 52512 10616
rect 52472 10130 52500 10610
rect 52460 10124 52512 10130
rect 52460 10066 52512 10072
rect 52564 7478 52592 15846
rect 52644 15156 52696 15162
rect 52644 15098 52696 15104
rect 52656 14074 52684 15098
rect 52644 14068 52696 14074
rect 52644 14010 52696 14016
rect 52644 11008 52696 11014
rect 52644 10950 52696 10956
rect 52656 10742 52684 10950
rect 52644 10736 52696 10742
rect 52644 10678 52696 10684
rect 52840 10577 52868 18158
rect 54312 18068 54340 18906
rect 54496 18612 54524 20334
rect 54772 19990 54800 20334
rect 54944 20324 54996 20330
rect 54944 20266 54996 20272
rect 54760 19984 54812 19990
rect 54760 19926 54812 19932
rect 54956 19718 54984 20266
rect 54944 19712 54996 19718
rect 54944 19654 54996 19660
rect 54576 18624 54628 18630
rect 54496 18584 54576 18612
rect 54576 18566 54628 18572
rect 54588 18290 54616 18566
rect 54576 18284 54628 18290
rect 54576 18226 54628 18232
rect 54392 18080 54444 18086
rect 54312 18040 54392 18068
rect 54312 17882 54340 18040
rect 54392 18022 54444 18028
rect 54300 17876 54352 17882
rect 54300 17818 54352 17824
rect 54300 17536 54352 17542
rect 54300 17478 54352 17484
rect 53196 16992 53248 16998
rect 53196 16934 53248 16940
rect 53104 16448 53156 16454
rect 53104 16390 53156 16396
rect 53116 15434 53144 16390
rect 53208 16250 53236 16934
rect 53840 16584 53892 16590
rect 53840 16526 53892 16532
rect 53852 16250 53880 16526
rect 53196 16244 53248 16250
rect 53196 16186 53248 16192
rect 53840 16244 53892 16250
rect 53840 16186 53892 16192
rect 53208 15434 53236 16186
rect 53748 16040 53800 16046
rect 53748 15982 53800 15988
rect 53760 15434 53788 15982
rect 54116 15904 54168 15910
rect 54116 15846 54168 15852
rect 54208 15904 54260 15910
rect 54208 15846 54260 15852
rect 53104 15428 53156 15434
rect 53104 15370 53156 15376
rect 53196 15428 53248 15434
rect 53196 15370 53248 15376
rect 53748 15428 53800 15434
rect 53748 15370 53800 15376
rect 53208 15162 53236 15370
rect 53196 15156 53248 15162
rect 53196 15098 53248 15104
rect 53656 14408 53708 14414
rect 53656 14350 53708 14356
rect 53012 14272 53064 14278
rect 53012 14214 53064 14220
rect 53024 13326 53052 14214
rect 53668 14074 53696 14350
rect 53656 14068 53708 14074
rect 53656 14010 53708 14016
rect 53760 13954 53788 15370
rect 54128 15094 54156 15846
rect 54220 15706 54248 15846
rect 54208 15700 54260 15706
rect 54208 15642 54260 15648
rect 54312 15586 54340 17478
rect 54588 16658 54616 18226
rect 54852 18216 54904 18222
rect 54852 18158 54904 18164
rect 54864 17746 54892 18158
rect 54852 17740 54904 17746
rect 54852 17682 54904 17688
rect 54576 16652 54628 16658
rect 54576 16594 54628 16600
rect 54220 15558 54340 15586
rect 54116 15088 54168 15094
rect 54116 15030 54168 15036
rect 53668 13926 53788 13954
rect 53668 13870 53696 13926
rect 53656 13864 53708 13870
rect 53656 13806 53708 13812
rect 53012 13320 53064 13326
rect 53012 13262 53064 13268
rect 54116 13320 54168 13326
rect 54116 13262 54168 13268
rect 54128 12442 54156 13262
rect 54116 12436 54168 12442
rect 54116 12378 54168 12384
rect 53012 11144 53064 11150
rect 53012 11086 53064 11092
rect 53024 10674 53052 11086
rect 53012 10668 53064 10674
rect 53012 10610 53064 10616
rect 53196 10668 53248 10674
rect 53196 10610 53248 10616
rect 52826 10568 52882 10577
rect 52826 10503 52882 10512
rect 52644 9920 52696 9926
rect 52644 9862 52696 9868
rect 52552 7472 52604 7478
rect 52552 7414 52604 7420
rect 52656 7206 52684 9862
rect 53208 9722 53236 10610
rect 53840 10260 53892 10266
rect 53840 10202 53892 10208
rect 53196 9716 53248 9722
rect 53196 9658 53248 9664
rect 53852 9586 53880 10202
rect 54024 9988 54076 9994
rect 54024 9930 54076 9936
rect 54036 9586 54064 9930
rect 54116 9920 54168 9926
rect 54116 9862 54168 9868
rect 53840 9580 53892 9586
rect 53840 9522 53892 9528
rect 54024 9580 54076 9586
rect 54024 9522 54076 9528
rect 54128 9466 54156 9862
rect 53760 9438 54156 9466
rect 53012 9376 53064 9382
rect 53012 9318 53064 9324
rect 53472 9376 53524 9382
rect 53472 9318 53524 9324
rect 53024 8974 53052 9318
rect 53012 8968 53064 8974
rect 53012 8910 53064 8916
rect 52920 8832 52972 8838
rect 52920 8774 52972 8780
rect 52932 8634 52960 8774
rect 52920 8628 52972 8634
rect 52920 8570 52972 8576
rect 52828 8492 52880 8498
rect 52828 8434 52880 8440
rect 52840 8090 52868 8434
rect 52828 8084 52880 8090
rect 52828 8026 52880 8032
rect 52644 7200 52696 7206
rect 52644 7142 52696 7148
rect 52656 6866 52684 7142
rect 52460 6860 52512 6866
rect 52460 6802 52512 6808
rect 52644 6860 52696 6866
rect 52644 6802 52696 6808
rect 52472 4690 52500 6802
rect 52552 6316 52604 6322
rect 52552 6258 52604 6264
rect 52564 5370 52592 6258
rect 52552 5364 52604 5370
rect 52552 5306 52604 5312
rect 52656 5302 52684 6802
rect 52840 6322 52868 8026
rect 53024 7834 53052 8910
rect 52932 7806 53052 7834
rect 52932 7206 52960 7806
rect 53484 7546 53512 9318
rect 53760 8838 53788 9438
rect 53932 9104 53984 9110
rect 53932 9046 53984 9052
rect 53748 8832 53800 8838
rect 53746 8800 53748 8809
rect 53800 8800 53802 8809
rect 53746 8735 53802 8744
rect 53760 7834 53788 8735
rect 53944 7954 53972 9046
rect 54024 8968 54076 8974
rect 54024 8910 54076 8916
rect 54036 8378 54064 8910
rect 54036 8350 54156 8378
rect 54024 8288 54076 8294
rect 54024 8230 54076 8236
rect 53932 7948 53984 7954
rect 53932 7890 53984 7896
rect 53760 7806 53880 7834
rect 53472 7540 53524 7546
rect 53472 7482 53524 7488
rect 52920 7200 52972 7206
rect 52920 7142 52972 7148
rect 52828 6316 52880 6322
rect 52828 6258 52880 6264
rect 52840 5710 52868 6258
rect 52828 5704 52880 5710
rect 52734 5672 52790 5681
rect 52828 5646 52880 5652
rect 52734 5607 52736 5616
rect 52788 5607 52790 5616
rect 52736 5578 52788 5584
rect 52644 5296 52696 5302
rect 52644 5238 52696 5244
rect 52552 5024 52604 5030
rect 52552 4966 52604 4972
rect 52564 4826 52592 4966
rect 52552 4820 52604 4826
rect 52552 4762 52604 4768
rect 52460 4684 52512 4690
rect 52460 4626 52512 4632
rect 52564 4010 52592 4762
rect 52736 4480 52788 4486
rect 52736 4422 52788 4428
rect 52748 4146 52776 4422
rect 52736 4140 52788 4146
rect 52736 4082 52788 4088
rect 52644 4072 52696 4078
rect 52644 4014 52696 4020
rect 52552 4004 52604 4010
rect 52552 3946 52604 3952
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 52564 2990 52592 3946
rect 52552 2984 52604 2990
rect 52552 2926 52604 2932
rect 52184 2916 52236 2922
rect 52184 2858 52236 2864
rect 52196 2446 52224 2858
rect 52656 2774 52684 4014
rect 52840 3534 52868 5646
rect 52932 4078 52960 7142
rect 53196 6928 53248 6934
rect 53196 6870 53248 6876
rect 53104 6656 53156 6662
rect 53104 6598 53156 6604
rect 53116 6458 53144 6598
rect 53208 6458 53236 6870
rect 53104 6452 53156 6458
rect 53104 6394 53156 6400
rect 53196 6452 53248 6458
rect 53196 6394 53248 6400
rect 53116 5302 53144 6394
rect 53380 5908 53432 5914
rect 53380 5850 53432 5856
rect 53104 5296 53156 5302
rect 53104 5238 53156 5244
rect 53012 5160 53064 5166
rect 53012 5102 53064 5108
rect 52920 4072 52972 4078
rect 52920 4014 52972 4020
rect 52828 3528 52880 3534
rect 52828 3470 52880 3476
rect 52840 3058 52868 3470
rect 52828 3052 52880 3058
rect 52828 2994 52880 3000
rect 52656 2746 52776 2774
rect 52460 2508 52512 2514
rect 52288 2468 52460 2496
rect 52184 2440 52236 2446
rect 52184 2382 52236 2388
rect 52288 800 52316 2468
rect 52460 2450 52512 2456
rect 52748 2446 52776 2746
rect 53024 2632 53052 5102
rect 53116 4622 53144 5238
rect 53392 5234 53420 5850
rect 53380 5228 53432 5234
rect 53380 5170 53432 5176
rect 53852 5030 53880 7806
rect 54036 7546 54064 8230
rect 54128 7546 54156 8350
rect 54024 7540 54076 7546
rect 54024 7482 54076 7488
rect 54116 7540 54168 7546
rect 54116 7482 54168 7488
rect 54220 7313 54248 15558
rect 54484 15360 54536 15366
rect 54484 15302 54536 15308
rect 54300 14612 54352 14618
rect 54300 14554 54352 14560
rect 54312 13954 54340 14554
rect 54312 13926 54432 13954
rect 54300 12436 54352 12442
rect 54300 12378 54352 12384
rect 54312 9024 54340 12378
rect 54404 10130 54432 13926
rect 54496 12306 54524 15302
rect 54484 12300 54536 12306
rect 54484 12242 54536 12248
rect 54588 11898 54616 16594
rect 54668 16040 54720 16046
rect 54668 15982 54720 15988
rect 54680 15706 54708 15982
rect 54668 15700 54720 15706
rect 54668 15642 54720 15648
rect 54852 15564 54904 15570
rect 54852 15506 54904 15512
rect 54760 15360 54812 15366
rect 54760 15302 54812 15308
rect 54772 15162 54800 15302
rect 54760 15156 54812 15162
rect 54760 15098 54812 15104
rect 54864 14618 54892 15506
rect 54852 14612 54904 14618
rect 54852 14554 54904 14560
rect 54944 13864 54996 13870
rect 54944 13806 54996 13812
rect 54760 13728 54812 13734
rect 54760 13670 54812 13676
rect 54772 13394 54800 13670
rect 54956 13394 54984 13806
rect 54760 13388 54812 13394
rect 54760 13330 54812 13336
rect 54944 13388 54996 13394
rect 54944 13330 54996 13336
rect 54944 13184 54996 13190
rect 54944 13126 54996 13132
rect 54956 12986 54984 13126
rect 54944 12980 54996 12986
rect 54944 12922 54996 12928
rect 55048 12434 55076 20742
rect 55404 20392 55456 20398
rect 55404 20334 55456 20340
rect 55496 20392 55548 20398
rect 55496 20334 55548 20340
rect 55416 19854 55444 20334
rect 55508 20058 55536 20334
rect 55496 20052 55548 20058
rect 55496 19994 55548 20000
rect 55404 19848 55456 19854
rect 55404 19790 55456 19796
rect 55416 19514 55444 19790
rect 55404 19508 55456 19514
rect 55404 19450 55456 19456
rect 55600 18630 55628 20742
rect 55772 20256 55824 20262
rect 55772 20198 55824 20204
rect 55784 18766 55812 20198
rect 55864 19780 55916 19786
rect 55864 19722 55916 19728
rect 55876 19514 55904 19722
rect 55864 19508 55916 19514
rect 55864 19450 55916 19456
rect 55772 18760 55824 18766
rect 55772 18702 55824 18708
rect 55588 18624 55640 18630
rect 55588 18566 55640 18572
rect 55680 18624 55732 18630
rect 55680 18566 55732 18572
rect 55600 18306 55628 18566
rect 55692 18426 55720 18566
rect 55680 18420 55732 18426
rect 55680 18362 55732 18368
rect 55600 18278 55720 18306
rect 55692 17542 55720 18278
rect 55680 17536 55732 17542
rect 55680 17478 55732 17484
rect 55692 17066 55720 17478
rect 55680 17060 55732 17066
rect 55680 17002 55732 17008
rect 55772 16516 55824 16522
rect 55772 16458 55824 16464
rect 55784 16250 55812 16458
rect 55772 16244 55824 16250
rect 55772 16186 55824 16192
rect 55784 15570 55812 16186
rect 55772 15564 55824 15570
rect 55772 15506 55824 15512
rect 55220 14816 55272 14822
rect 55220 14758 55272 14764
rect 55784 14770 55812 15506
rect 55968 15450 55996 20946
rect 56060 20534 56088 21286
rect 56612 21146 56640 21422
rect 56600 21140 56652 21146
rect 56600 21082 56652 21088
rect 57520 20936 57572 20942
rect 57520 20878 57572 20884
rect 56784 20868 56836 20874
rect 56784 20810 56836 20816
rect 56140 20800 56192 20806
rect 56140 20742 56192 20748
rect 56048 20528 56100 20534
rect 56048 20470 56100 20476
rect 56152 19310 56180 20742
rect 56796 20058 56824 20810
rect 57532 20602 57560 20878
rect 58726 20700 59034 20709
rect 58726 20698 58732 20700
rect 58788 20698 58812 20700
rect 58868 20698 58892 20700
rect 58948 20698 58972 20700
rect 59028 20698 59034 20700
rect 58788 20646 58790 20698
rect 58970 20646 58972 20698
rect 58726 20644 58732 20646
rect 58788 20644 58812 20646
rect 58868 20644 58892 20646
rect 58948 20644 58972 20646
rect 59028 20644 59034 20646
rect 58726 20635 59034 20644
rect 57520 20596 57572 20602
rect 57520 20538 57572 20544
rect 56784 20052 56836 20058
rect 56784 19994 56836 20000
rect 58726 19612 59034 19621
rect 58726 19610 58732 19612
rect 58788 19610 58812 19612
rect 58868 19610 58892 19612
rect 58948 19610 58972 19612
rect 59028 19610 59034 19612
rect 58788 19558 58790 19610
rect 58970 19558 58972 19610
rect 58726 19556 58732 19558
rect 58788 19556 58812 19558
rect 58868 19556 58892 19558
rect 58948 19556 58972 19558
rect 59028 19556 59034 19558
rect 58726 19547 59034 19556
rect 56140 19304 56192 19310
rect 56140 19246 56192 19252
rect 58164 18896 58216 18902
rect 58164 18838 58216 18844
rect 56324 18828 56376 18834
rect 56324 18770 56376 18776
rect 56232 18624 56284 18630
rect 56232 18566 56284 18572
rect 56244 18358 56272 18566
rect 56232 18352 56284 18358
rect 56232 18294 56284 18300
rect 56140 18080 56192 18086
rect 56140 18022 56192 18028
rect 56152 17678 56180 18022
rect 56140 17672 56192 17678
rect 56140 17614 56192 17620
rect 56152 16998 56180 17614
rect 56140 16992 56192 16998
rect 56140 16934 56192 16940
rect 56048 15972 56100 15978
rect 56048 15914 56100 15920
rect 56060 15570 56088 15914
rect 56152 15910 56180 16934
rect 56140 15904 56192 15910
rect 56140 15846 56192 15852
rect 56048 15564 56100 15570
rect 56048 15506 56100 15512
rect 55968 15422 56088 15450
rect 55128 13184 55180 13190
rect 55128 13126 55180 13132
rect 55140 12918 55168 13126
rect 55232 12986 55260 14758
rect 55784 14742 55996 14770
rect 55312 13864 55364 13870
rect 55312 13806 55364 13812
rect 55324 13462 55352 13806
rect 55312 13456 55364 13462
rect 55312 13398 55364 13404
rect 55220 12980 55272 12986
rect 55220 12922 55272 12928
rect 55128 12912 55180 12918
rect 55128 12854 55180 12860
rect 55232 12646 55260 12922
rect 55324 12714 55352 13398
rect 55968 13326 55996 14742
rect 55956 13320 56008 13326
rect 55956 13262 56008 13268
rect 55968 12850 55996 13262
rect 55956 12844 56008 12850
rect 55956 12786 56008 12792
rect 55312 12708 55364 12714
rect 55312 12650 55364 12656
rect 55220 12640 55272 12646
rect 55220 12582 55272 12588
rect 54772 12406 55076 12434
rect 54576 11892 54628 11898
rect 54576 11834 54628 11840
rect 54576 10600 54628 10606
rect 54576 10542 54628 10548
rect 54484 10464 54536 10470
rect 54484 10406 54536 10412
rect 54392 10124 54444 10130
rect 54392 10066 54444 10072
rect 54392 9036 54444 9042
rect 54312 8996 54392 9024
rect 54392 8978 54444 8984
rect 54206 7304 54262 7313
rect 54206 7239 54262 7248
rect 54404 7002 54432 8978
rect 54496 7886 54524 10406
rect 54588 9586 54616 10542
rect 54576 9580 54628 9586
rect 54576 9522 54628 9528
rect 54668 8968 54720 8974
rect 54668 8910 54720 8916
rect 54680 8430 54708 8910
rect 54668 8424 54720 8430
rect 54668 8366 54720 8372
rect 54484 7880 54536 7886
rect 54484 7822 54536 7828
rect 54772 7206 54800 12406
rect 55128 11892 55180 11898
rect 55128 11834 55180 11840
rect 55036 11144 55088 11150
rect 55036 11086 55088 11092
rect 55048 10266 55076 11086
rect 55140 10674 55168 11834
rect 55232 11762 55260 12582
rect 55220 11756 55272 11762
rect 55220 11698 55272 11704
rect 55128 10668 55180 10674
rect 55128 10610 55180 10616
rect 55036 10260 55088 10266
rect 55036 10202 55088 10208
rect 55140 9058 55168 10610
rect 55232 10470 55260 11698
rect 55404 11280 55456 11286
rect 55404 11222 55456 11228
rect 55416 10674 55444 11222
rect 55404 10668 55456 10674
rect 55404 10610 55456 10616
rect 55220 10464 55272 10470
rect 55220 10406 55272 10412
rect 54956 9030 55168 9058
rect 54956 8514 54984 9030
rect 55232 8786 55260 10406
rect 55416 10130 55444 10610
rect 55404 10124 55456 10130
rect 55404 10066 55456 10072
rect 55864 9512 55916 9518
rect 55864 9454 55916 9460
rect 55876 9178 55904 9454
rect 55864 9172 55916 9178
rect 55864 9114 55916 9120
rect 56060 9081 56088 15422
rect 56152 14822 56180 15846
rect 56232 15496 56284 15502
rect 56232 15438 56284 15444
rect 56336 15450 56364 18770
rect 56600 18760 56652 18766
rect 56600 18702 56652 18708
rect 56612 17882 56640 18702
rect 56968 18624 57020 18630
rect 56968 18566 57020 18572
rect 57244 18624 57296 18630
rect 57244 18566 57296 18572
rect 56692 18420 56744 18426
rect 56692 18362 56744 18368
rect 56704 17882 56732 18362
rect 56600 17876 56652 17882
rect 56600 17818 56652 17824
rect 56692 17876 56744 17882
rect 56692 17818 56744 17824
rect 56980 17678 57008 18566
rect 57256 18426 57284 18566
rect 57244 18420 57296 18426
rect 57244 18362 57296 18368
rect 57704 18216 57756 18222
rect 57704 18158 57756 18164
rect 57336 18080 57388 18086
rect 57336 18022 57388 18028
rect 56968 17672 57020 17678
rect 56968 17614 57020 17620
rect 57348 17338 57376 18022
rect 57716 17882 57744 18158
rect 57704 17876 57756 17882
rect 57704 17818 57756 17824
rect 57336 17332 57388 17338
rect 57336 17274 57388 17280
rect 56876 17128 56928 17134
rect 56876 17070 56928 17076
rect 57704 17128 57756 17134
rect 57704 17070 57756 17076
rect 56784 16448 56836 16454
rect 56784 16390 56836 16396
rect 56796 15638 56824 16390
rect 56784 15632 56836 15638
rect 56784 15574 56836 15580
rect 56508 15564 56560 15570
rect 56508 15506 56560 15512
rect 56600 15564 56652 15570
rect 56600 15506 56652 15512
rect 56244 15026 56272 15438
rect 56336 15422 56456 15450
rect 56324 15360 56376 15366
rect 56324 15302 56376 15308
rect 56232 15020 56284 15026
rect 56232 14962 56284 14968
rect 56140 14816 56192 14822
rect 56140 14758 56192 14764
rect 56152 13734 56180 14758
rect 56336 13734 56364 15302
rect 56140 13728 56192 13734
rect 56140 13670 56192 13676
rect 56324 13728 56376 13734
rect 56324 13670 56376 13676
rect 56152 12850 56180 13670
rect 56428 12866 56456 15422
rect 56520 13394 56548 15506
rect 56612 13954 56640 15506
rect 56796 15366 56824 15574
rect 56784 15360 56836 15366
rect 56784 15302 56836 15308
rect 56796 14278 56824 15302
rect 56784 14272 56836 14278
rect 56784 14214 56836 14220
rect 56612 13926 56732 13954
rect 56508 13388 56560 13394
rect 56508 13330 56560 13336
rect 56600 13388 56652 13394
rect 56600 13330 56652 13336
rect 56520 12986 56548 13330
rect 56508 12980 56560 12986
rect 56508 12922 56560 12928
rect 56612 12866 56640 13330
rect 56704 13297 56732 13926
rect 56690 13288 56746 13297
rect 56690 13223 56746 13232
rect 56140 12844 56192 12850
rect 56140 12786 56192 12792
rect 56428 12838 56640 12866
rect 56232 12096 56284 12102
rect 56232 12038 56284 12044
rect 56244 9654 56272 12038
rect 56428 10810 56456 12838
rect 56600 11552 56652 11558
rect 56600 11494 56652 11500
rect 56612 11150 56640 11494
rect 56600 11144 56652 11150
rect 56600 11086 56652 11092
rect 56600 11008 56652 11014
rect 56600 10950 56652 10956
rect 56416 10804 56468 10810
rect 56416 10746 56468 10752
rect 56612 10674 56640 10950
rect 56704 10690 56732 13223
rect 56796 12986 56824 14214
rect 56784 12980 56836 12986
rect 56784 12922 56836 12928
rect 56796 12102 56824 12922
rect 56784 12096 56836 12102
rect 56784 12038 56836 12044
rect 56600 10668 56652 10674
rect 56704 10662 56824 10690
rect 56600 10610 56652 10616
rect 56692 10600 56744 10606
rect 56692 10542 56744 10548
rect 56324 10464 56376 10470
rect 56324 10406 56376 10412
rect 56600 10464 56652 10470
rect 56600 10406 56652 10412
rect 56336 9926 56364 10406
rect 56324 9920 56376 9926
rect 56324 9862 56376 9868
rect 56232 9648 56284 9654
rect 56232 9590 56284 9596
rect 56324 9376 56376 9382
rect 56324 9318 56376 9324
rect 56046 9072 56102 9081
rect 56046 9007 56102 9016
rect 55232 8758 55352 8786
rect 55220 8628 55272 8634
rect 55220 8570 55272 8576
rect 54864 8498 54984 8514
rect 54852 8492 54984 8498
rect 54904 8486 54984 8492
rect 54852 8434 54904 8440
rect 54956 8022 54984 8486
rect 55128 8424 55180 8430
rect 55128 8366 55180 8372
rect 55140 8090 55168 8366
rect 55128 8084 55180 8090
rect 55128 8026 55180 8032
rect 54944 8016 54996 8022
rect 54944 7958 54996 7964
rect 54760 7200 54812 7206
rect 54760 7142 54812 7148
rect 54392 6996 54444 7002
rect 54392 6938 54444 6944
rect 54116 6656 54168 6662
rect 54116 6598 54168 6604
rect 54128 6458 54156 6598
rect 54116 6452 54168 6458
rect 54116 6394 54168 6400
rect 54956 6322 54984 7958
rect 55140 7410 55168 8026
rect 55232 7954 55260 8570
rect 55324 8430 55352 8758
rect 56336 8498 56364 9318
rect 56324 8492 56376 8498
rect 56324 8434 56376 8440
rect 55312 8424 55364 8430
rect 55312 8366 55364 8372
rect 56140 8424 56192 8430
rect 56140 8366 56192 8372
rect 55220 7948 55272 7954
rect 55220 7890 55272 7896
rect 55864 7948 55916 7954
rect 55864 7890 55916 7896
rect 55312 7744 55364 7750
rect 55312 7686 55364 7692
rect 55128 7404 55180 7410
rect 55128 7346 55180 7352
rect 54944 6316 54996 6322
rect 54944 6258 54996 6264
rect 54024 5636 54076 5642
rect 54024 5578 54076 5584
rect 54036 5370 54064 5578
rect 54956 5370 54984 6258
rect 55220 6248 55272 6254
rect 55220 6190 55272 6196
rect 55232 5914 55260 6190
rect 55220 5908 55272 5914
rect 55220 5850 55272 5856
rect 54024 5364 54076 5370
rect 54024 5306 54076 5312
rect 54944 5364 54996 5370
rect 54944 5306 54996 5312
rect 53748 5024 53800 5030
rect 53748 4966 53800 4972
rect 53840 5024 53892 5030
rect 53840 4966 53892 4972
rect 53104 4616 53156 4622
rect 53104 4558 53156 4564
rect 53116 4078 53144 4558
rect 53196 4480 53248 4486
rect 53196 4422 53248 4428
rect 53564 4480 53616 4486
rect 53564 4422 53616 4428
rect 53104 4072 53156 4078
rect 53104 4014 53156 4020
rect 53208 3738 53236 4422
rect 53196 3732 53248 3738
rect 53196 3674 53248 3680
rect 53576 3126 53604 4422
rect 53564 3120 53616 3126
rect 53564 3062 53616 3068
rect 53380 2848 53432 2854
rect 53380 2790 53432 2796
rect 52840 2604 53052 2632
rect 52736 2440 52788 2446
rect 52736 2382 52788 2388
rect 52840 800 52868 2604
rect 53392 800 53420 2790
rect 53760 2514 53788 4966
rect 54024 4684 54076 4690
rect 54024 4626 54076 4632
rect 53932 4208 53984 4214
rect 53932 4150 53984 4156
rect 53944 3738 53972 4150
rect 54036 4078 54064 4626
rect 54116 4616 54168 4622
rect 54116 4558 54168 4564
rect 54128 4078 54156 4558
rect 54956 4162 54984 5306
rect 55220 5092 55272 5098
rect 55220 5034 55272 5040
rect 54772 4146 54984 4162
rect 54760 4140 54984 4146
rect 54812 4134 54984 4140
rect 54760 4082 54812 4088
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54116 4072 54168 4078
rect 54116 4014 54168 4020
rect 54852 4072 54904 4078
rect 54852 4014 54904 4020
rect 55036 4072 55088 4078
rect 55036 4014 55088 4020
rect 54024 3936 54076 3942
rect 54024 3878 54076 3884
rect 53932 3732 53984 3738
rect 53932 3674 53984 3680
rect 54036 3194 54064 3878
rect 54864 3534 54892 4014
rect 55048 3738 55076 4014
rect 55232 3738 55260 5034
rect 55324 4282 55352 7686
rect 55588 7472 55640 7478
rect 55588 7414 55640 7420
rect 55496 7200 55548 7206
rect 55496 7142 55548 7148
rect 55508 6905 55536 7142
rect 55600 7002 55628 7414
rect 55876 7342 55904 7890
rect 56152 7750 56180 8366
rect 56140 7744 56192 7750
rect 56140 7686 56192 7692
rect 56508 7744 56560 7750
rect 56508 7686 56560 7692
rect 56520 7342 56548 7686
rect 55864 7336 55916 7342
rect 55864 7278 55916 7284
rect 56508 7336 56560 7342
rect 56508 7278 56560 7284
rect 55876 7041 55904 7278
rect 55862 7032 55918 7041
rect 55588 6996 55640 7002
rect 55862 6967 55918 6976
rect 55588 6938 55640 6944
rect 55494 6896 55550 6905
rect 55494 6831 55496 6840
rect 55548 6831 55550 6840
rect 55496 6802 55548 6808
rect 55600 6254 55628 6938
rect 56612 6934 56640 10406
rect 56704 10266 56732 10542
rect 56796 10470 56824 10662
rect 56784 10464 56836 10470
rect 56784 10406 56836 10412
rect 56692 10260 56744 10266
rect 56692 10202 56744 10208
rect 56692 9648 56744 9654
rect 56692 9590 56744 9596
rect 56704 9178 56732 9590
rect 56784 9512 56836 9518
rect 56784 9454 56836 9460
rect 56692 9172 56744 9178
rect 56692 9114 56744 9120
rect 56600 6928 56652 6934
rect 56600 6870 56652 6876
rect 55956 6656 56008 6662
rect 55956 6598 56008 6604
rect 55588 6248 55640 6254
rect 55588 6190 55640 6196
rect 55404 5024 55456 5030
rect 55404 4966 55456 4972
rect 55312 4276 55364 4282
rect 55312 4218 55364 4224
rect 55416 3754 55444 4966
rect 55496 4616 55548 4622
rect 55496 4558 55548 4564
rect 55508 4282 55536 4558
rect 55496 4276 55548 4282
rect 55496 4218 55548 4224
rect 55600 4078 55628 6190
rect 55864 6112 55916 6118
rect 55864 6054 55916 6060
rect 55680 5636 55732 5642
rect 55680 5578 55732 5584
rect 55692 5370 55720 5578
rect 55680 5364 55732 5370
rect 55680 5306 55732 5312
rect 55680 4616 55732 4622
rect 55680 4558 55732 4564
rect 55772 4616 55824 4622
rect 55772 4558 55824 4564
rect 55588 4072 55640 4078
rect 55588 4014 55640 4020
rect 55036 3732 55088 3738
rect 55036 3674 55088 3680
rect 55220 3732 55272 3738
rect 55220 3674 55272 3680
rect 55324 3726 55444 3754
rect 54852 3528 54904 3534
rect 54852 3470 54904 3476
rect 54116 3392 54168 3398
rect 54116 3334 54168 3340
rect 54128 3194 54156 3334
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 54116 3188 54168 3194
rect 54116 3130 54168 3136
rect 54484 3052 54536 3058
rect 54484 2994 54536 3000
rect 53932 2984 53984 2990
rect 53932 2926 53984 2932
rect 53748 2508 53800 2514
rect 53748 2450 53800 2456
rect 53944 800 53972 2926
rect 54496 800 54524 2994
rect 55036 2984 55088 2990
rect 55036 2926 55088 2932
rect 55048 800 55076 2926
rect 55324 2650 55352 3726
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55312 2644 55364 2650
rect 55312 2586 55364 2592
rect 55416 2514 55444 2790
rect 55404 2508 55456 2514
rect 55404 2450 55456 2456
rect 55692 2446 55720 4558
rect 55784 4078 55812 4558
rect 55876 4214 55904 6054
rect 55968 5234 55996 6598
rect 56704 6338 56732 9114
rect 56796 9110 56824 9454
rect 56784 9104 56836 9110
rect 56784 9046 56836 9052
rect 56796 7546 56824 9046
rect 56888 8945 56916 17070
rect 57060 16652 57112 16658
rect 57060 16594 57112 16600
rect 56968 10668 57020 10674
rect 56968 10610 57020 10616
rect 56980 9518 57008 10610
rect 57072 9518 57100 16594
rect 57428 16448 57480 16454
rect 57428 16390 57480 16396
rect 57440 16250 57468 16390
rect 57716 16250 57744 17070
rect 57888 16992 57940 16998
rect 57888 16934 57940 16940
rect 57900 16590 57928 16934
rect 57888 16584 57940 16590
rect 57888 16526 57940 16532
rect 57428 16244 57480 16250
rect 57428 16186 57480 16192
rect 57704 16244 57756 16250
rect 57704 16186 57756 16192
rect 57152 16108 57204 16114
rect 57152 16050 57204 16056
rect 57164 15570 57192 16050
rect 57716 15706 57744 16186
rect 57888 15904 57940 15910
rect 57888 15846 57940 15852
rect 57900 15706 57928 15846
rect 57244 15700 57296 15706
rect 57244 15642 57296 15648
rect 57704 15700 57756 15706
rect 57704 15642 57756 15648
rect 57888 15700 57940 15706
rect 57888 15642 57940 15648
rect 57256 15570 57284 15642
rect 57152 15564 57204 15570
rect 57152 15506 57204 15512
rect 57244 15564 57296 15570
rect 57244 15506 57296 15512
rect 57164 15162 57192 15506
rect 57980 15360 58032 15366
rect 57980 15302 58032 15308
rect 57152 15156 57204 15162
rect 57152 15098 57204 15104
rect 57992 15026 58020 15302
rect 57980 15020 58032 15026
rect 57980 14962 58032 14968
rect 57888 14340 57940 14346
rect 57888 14282 57940 14288
rect 57336 14272 57388 14278
rect 57336 14214 57388 14220
rect 57348 14074 57376 14214
rect 57900 14074 57928 14282
rect 57336 14068 57388 14074
rect 57336 14010 57388 14016
rect 57888 14068 57940 14074
rect 57888 14010 57940 14016
rect 57704 13796 57756 13802
rect 57704 13738 57756 13744
rect 57612 13728 57664 13734
rect 57612 13670 57664 13676
rect 57624 13326 57652 13670
rect 57716 13394 57744 13738
rect 57704 13388 57756 13394
rect 57704 13330 57756 13336
rect 57152 13320 57204 13326
rect 57152 13262 57204 13268
rect 57612 13320 57664 13326
rect 57612 13262 57664 13268
rect 57164 12986 57192 13262
rect 57520 13184 57572 13190
rect 57520 13126 57572 13132
rect 57152 12980 57204 12986
rect 57152 12922 57204 12928
rect 57244 12844 57296 12850
rect 57244 12786 57296 12792
rect 57256 12442 57284 12786
rect 57244 12436 57296 12442
rect 57532 12434 57560 13126
rect 57612 12640 57664 12646
rect 57612 12582 57664 12588
rect 57244 12378 57296 12384
rect 57440 12406 57560 12434
rect 57152 11688 57204 11694
rect 57152 11630 57204 11636
rect 56968 9512 57020 9518
rect 56968 9454 57020 9460
rect 57060 9512 57112 9518
rect 57060 9454 57112 9460
rect 56874 8936 56930 8945
rect 56874 8871 56930 8880
rect 56876 8832 56928 8838
rect 56874 8800 56876 8809
rect 56980 8820 57008 9454
rect 57164 9382 57192 11630
rect 57152 9376 57204 9382
rect 57152 9318 57204 9324
rect 57244 9036 57296 9042
rect 57244 8978 57296 8984
rect 56928 8800 57008 8820
rect 56930 8792 57008 8800
rect 56874 8735 56930 8744
rect 56784 7540 56836 7546
rect 56784 7482 56836 7488
rect 56796 6866 56824 7482
rect 56784 6860 56836 6866
rect 56784 6802 56836 6808
rect 56784 6656 56836 6662
rect 56784 6598 56836 6604
rect 56968 6656 57020 6662
rect 56968 6598 57020 6604
rect 56612 6310 56732 6338
rect 56508 5636 56560 5642
rect 56508 5578 56560 5584
rect 55956 5228 56008 5234
rect 55956 5170 56008 5176
rect 56140 5160 56192 5166
rect 56140 5102 56192 5108
rect 55956 4752 56008 4758
rect 55956 4694 56008 4700
rect 55864 4208 55916 4214
rect 55864 4150 55916 4156
rect 55968 4146 55996 4694
rect 56048 4480 56100 4486
rect 56048 4422 56100 4428
rect 55956 4140 56008 4146
rect 55956 4082 56008 4088
rect 55772 4072 55824 4078
rect 55772 4014 55824 4020
rect 55956 4004 56008 4010
rect 55956 3946 56008 3952
rect 55968 3194 55996 3946
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 56060 2774 56088 4422
rect 55784 2746 56088 2774
rect 55784 2650 55812 2746
rect 55772 2644 55824 2650
rect 55772 2586 55824 2592
rect 55772 2508 55824 2514
rect 55772 2450 55824 2456
rect 55680 2440 55732 2446
rect 55680 2382 55732 2388
rect 55784 1170 55812 2450
rect 55600 1142 55812 1170
rect 55600 800 55628 1142
rect 56152 800 56180 5102
rect 56520 4758 56548 5578
rect 56612 5166 56640 6310
rect 56692 6248 56744 6254
rect 56692 6190 56744 6196
rect 56704 5914 56732 6190
rect 56796 5914 56824 6598
rect 56692 5908 56744 5914
rect 56692 5850 56744 5856
rect 56784 5908 56836 5914
rect 56784 5850 56836 5856
rect 56704 5710 56732 5850
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56980 5234 57008 6598
rect 56968 5228 57020 5234
rect 56968 5170 57020 5176
rect 57152 5228 57204 5234
rect 57152 5170 57204 5176
rect 56600 5160 56652 5166
rect 56600 5102 56652 5108
rect 56508 4752 56560 4758
rect 56508 4694 56560 4700
rect 56600 4548 56652 4554
rect 56600 4490 56652 4496
rect 56416 4480 56468 4486
rect 56416 4422 56468 4428
rect 56428 4282 56456 4422
rect 56416 4276 56468 4282
rect 56416 4218 56468 4224
rect 56612 2394 56640 4490
rect 56980 4214 57008 5170
rect 57164 4826 57192 5170
rect 57152 4820 57204 4826
rect 57152 4762 57204 4768
rect 57060 4480 57112 4486
rect 57060 4422 57112 4428
rect 56968 4208 57020 4214
rect 56968 4150 57020 4156
rect 56692 4072 56744 4078
rect 56690 4040 56692 4049
rect 56744 4040 56746 4049
rect 56690 3975 56746 3984
rect 57072 3534 57100 4422
rect 57256 4078 57284 8978
rect 57336 5296 57388 5302
rect 57336 5238 57388 5244
rect 57440 5250 57468 12406
rect 57624 12238 57652 12582
rect 57612 12232 57664 12238
rect 57612 12174 57664 12180
rect 57612 12096 57664 12102
rect 57612 12038 57664 12044
rect 57520 9580 57572 9586
rect 57520 9522 57572 9528
rect 57532 9042 57560 9522
rect 57520 9036 57572 9042
rect 57520 8978 57572 8984
rect 57624 7546 57652 12038
rect 57796 11076 57848 11082
rect 57796 11018 57848 11024
rect 57704 10056 57756 10062
rect 57704 9998 57756 10004
rect 57716 8294 57744 9998
rect 57808 9654 57836 11018
rect 57888 10464 57940 10470
rect 57888 10406 57940 10412
rect 57900 10266 57928 10406
rect 57888 10260 57940 10266
rect 57888 10202 57940 10208
rect 57796 9648 57848 9654
rect 57796 9590 57848 9596
rect 57796 8900 57848 8906
rect 57796 8842 57848 8848
rect 57808 8634 57836 8842
rect 57888 8832 57940 8838
rect 57888 8774 57940 8780
rect 58072 8832 58124 8838
rect 58072 8774 58124 8780
rect 57796 8628 57848 8634
rect 57796 8570 57848 8576
rect 57704 8288 57756 8294
rect 57704 8230 57756 8236
rect 57716 7954 57744 8230
rect 57704 7948 57756 7954
rect 57704 7890 57756 7896
rect 57612 7540 57664 7546
rect 57612 7482 57664 7488
rect 57612 7404 57664 7410
rect 57612 7346 57664 7352
rect 57520 6656 57572 6662
rect 57520 6598 57572 6604
rect 57532 6458 57560 6598
rect 57520 6452 57572 6458
rect 57520 6394 57572 6400
rect 57520 5568 57572 5574
rect 57520 5510 57572 5516
rect 57532 5370 57560 5510
rect 57624 5370 57652 7346
rect 57716 6322 57744 7890
rect 57900 7546 57928 8774
rect 58084 7954 58112 8774
rect 58072 7948 58124 7954
rect 58072 7890 58124 7896
rect 57888 7540 57940 7546
rect 57888 7482 57940 7488
rect 58072 7472 58124 7478
rect 58072 7414 58124 7420
rect 57888 6860 57940 6866
rect 57888 6802 57940 6808
rect 57900 6458 57928 6802
rect 57980 6724 58032 6730
rect 57980 6666 58032 6672
rect 57888 6452 57940 6458
rect 57888 6394 57940 6400
rect 57704 6316 57756 6322
rect 57704 6258 57756 6264
rect 57716 5778 57744 6258
rect 57704 5772 57756 5778
rect 57704 5714 57756 5720
rect 57520 5364 57572 5370
rect 57520 5306 57572 5312
rect 57612 5364 57664 5370
rect 57612 5306 57664 5312
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57060 3528 57112 3534
rect 57060 3470 57112 3476
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 57164 2650 57192 3470
rect 57152 2644 57204 2650
rect 57152 2586 57204 2592
rect 56612 2366 56732 2394
rect 56704 800 56732 2366
rect 57256 800 57284 3538
rect 57348 2938 57376 5238
rect 57440 5222 57652 5250
rect 57428 4548 57480 4554
rect 57428 4490 57480 4496
rect 57440 3074 57468 4490
rect 57520 3936 57572 3942
rect 57520 3878 57572 3884
rect 57532 3194 57560 3878
rect 57520 3188 57572 3194
rect 57520 3130 57572 3136
rect 57440 3046 57560 3074
rect 57348 2910 57468 2938
rect 57440 2854 57468 2910
rect 57428 2848 57480 2854
rect 57428 2790 57480 2796
rect 57532 2446 57560 3046
rect 57624 2514 57652 5222
rect 57716 4826 57744 5714
rect 57796 5024 57848 5030
rect 57796 4966 57848 4972
rect 57704 4820 57756 4826
rect 57704 4762 57756 4768
rect 57716 3194 57744 4762
rect 57808 4622 57836 4966
rect 57796 4616 57848 4622
rect 57796 4558 57848 4564
rect 57992 4128 58020 6666
rect 57808 4100 58020 4128
rect 57704 3188 57756 3194
rect 57704 3130 57756 3136
rect 57704 3052 57756 3058
rect 57704 2994 57756 3000
rect 57716 2650 57744 2994
rect 57704 2644 57756 2650
rect 57704 2586 57756 2592
rect 57612 2508 57664 2514
rect 57612 2450 57664 2456
rect 57520 2440 57572 2446
rect 57520 2382 57572 2388
rect 57808 800 57836 4100
rect 57888 3460 57940 3466
rect 57888 3402 57940 3408
rect 57900 3194 57928 3402
rect 57888 3188 57940 3194
rect 57888 3130 57940 3136
rect 57980 2916 58032 2922
rect 57980 2858 58032 2864
rect 57992 2514 58020 2858
rect 57980 2508 58032 2514
rect 57980 2450 58032 2456
rect 51828 734 52132 762
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58084 762 58112 7414
rect 58176 4622 58204 18838
rect 58726 18524 59034 18533
rect 58726 18522 58732 18524
rect 58788 18522 58812 18524
rect 58868 18522 58892 18524
rect 58948 18522 58972 18524
rect 59028 18522 59034 18524
rect 58788 18470 58790 18522
rect 58970 18470 58972 18522
rect 58726 18468 58732 18470
rect 58788 18468 58812 18470
rect 58868 18468 58892 18470
rect 58948 18468 58972 18470
rect 59028 18468 59034 18470
rect 58726 18459 59034 18468
rect 58348 17672 58400 17678
rect 58348 17614 58400 17620
rect 58360 17338 58388 17614
rect 58726 17436 59034 17445
rect 58726 17434 58732 17436
rect 58788 17434 58812 17436
rect 58868 17434 58892 17436
rect 58948 17434 58972 17436
rect 59028 17434 59034 17436
rect 58788 17382 58790 17434
rect 58970 17382 58972 17434
rect 58726 17380 58732 17382
rect 58788 17380 58812 17382
rect 58868 17380 58892 17382
rect 58948 17380 58972 17382
rect 59028 17380 59034 17382
rect 58726 17371 59034 17380
rect 58348 17332 58400 17338
rect 58348 17274 58400 17280
rect 58256 17060 58308 17066
rect 58256 17002 58308 17008
rect 58268 9654 58296 17002
rect 58726 16348 59034 16357
rect 58726 16346 58732 16348
rect 58788 16346 58812 16348
rect 58868 16346 58892 16348
rect 58948 16346 58972 16348
rect 59028 16346 59034 16348
rect 58788 16294 58790 16346
rect 58970 16294 58972 16346
rect 58726 16292 58732 16294
rect 58788 16292 58812 16294
rect 58868 16292 58892 16294
rect 58948 16292 58972 16294
rect 59028 16292 59034 16294
rect 58726 16283 59034 16292
rect 58726 15260 59034 15269
rect 58726 15258 58732 15260
rect 58788 15258 58812 15260
rect 58868 15258 58892 15260
rect 58948 15258 58972 15260
rect 59028 15258 59034 15260
rect 58788 15206 58790 15258
rect 58970 15206 58972 15258
rect 58726 15204 58732 15206
rect 58788 15204 58812 15206
rect 58868 15204 58892 15206
rect 58948 15204 58972 15206
rect 59028 15204 59034 15206
rect 58726 15195 59034 15204
rect 58726 14172 59034 14181
rect 58726 14170 58732 14172
rect 58788 14170 58812 14172
rect 58868 14170 58892 14172
rect 58948 14170 58972 14172
rect 59028 14170 59034 14172
rect 58788 14118 58790 14170
rect 58970 14118 58972 14170
rect 58726 14116 58732 14118
rect 58788 14116 58812 14118
rect 58868 14116 58892 14118
rect 58948 14116 58972 14118
rect 59028 14116 59034 14118
rect 58726 14107 59034 14116
rect 58726 13084 59034 13093
rect 58726 13082 58732 13084
rect 58788 13082 58812 13084
rect 58868 13082 58892 13084
rect 58948 13082 58972 13084
rect 59028 13082 59034 13084
rect 58788 13030 58790 13082
rect 58970 13030 58972 13082
rect 58726 13028 58732 13030
rect 58788 13028 58812 13030
rect 58868 13028 58892 13030
rect 58948 13028 58972 13030
rect 59028 13028 59034 13030
rect 58726 13019 59034 13028
rect 58726 11996 59034 12005
rect 58726 11994 58732 11996
rect 58788 11994 58812 11996
rect 58868 11994 58892 11996
rect 58948 11994 58972 11996
rect 59028 11994 59034 11996
rect 58788 11942 58790 11994
rect 58970 11942 58972 11994
rect 58726 11940 58732 11942
rect 58788 11940 58812 11942
rect 58868 11940 58892 11942
rect 58948 11940 58972 11942
rect 59028 11940 59034 11942
rect 58726 11931 59034 11940
rect 58726 10908 59034 10917
rect 58726 10906 58732 10908
rect 58788 10906 58812 10908
rect 58868 10906 58892 10908
rect 58948 10906 58972 10908
rect 59028 10906 59034 10908
rect 58788 10854 58790 10906
rect 58970 10854 58972 10906
rect 58726 10852 58732 10854
rect 58788 10852 58812 10854
rect 58868 10852 58892 10854
rect 58948 10852 58972 10854
rect 59028 10852 59034 10854
rect 58726 10843 59034 10852
rect 58726 9820 59034 9829
rect 58726 9818 58732 9820
rect 58788 9818 58812 9820
rect 58868 9818 58892 9820
rect 58948 9818 58972 9820
rect 59028 9818 59034 9820
rect 58788 9766 58790 9818
rect 58970 9766 58972 9818
rect 58726 9764 58732 9766
rect 58788 9764 58812 9766
rect 58868 9764 58892 9766
rect 58948 9764 58972 9766
rect 59028 9764 59034 9766
rect 58726 9755 59034 9764
rect 58256 9648 58308 9654
rect 58256 9590 58308 9596
rect 58440 9580 58492 9586
rect 58440 9522 58492 9528
rect 58256 7268 58308 7274
rect 58256 7210 58308 7216
rect 58268 5710 58296 7210
rect 58348 6656 58400 6662
rect 58348 6598 58400 6604
rect 58256 5704 58308 5710
rect 58256 5646 58308 5652
rect 58164 4616 58216 4622
rect 58164 4558 58216 4564
rect 58360 2378 58388 6598
rect 58452 5914 58480 9522
rect 58726 8732 59034 8741
rect 58726 8730 58732 8732
rect 58788 8730 58812 8732
rect 58868 8730 58892 8732
rect 58948 8730 58972 8732
rect 59028 8730 59034 8732
rect 58788 8678 58790 8730
rect 58970 8678 58972 8730
rect 58726 8676 58732 8678
rect 58788 8676 58812 8678
rect 58868 8676 58892 8678
rect 58948 8676 58972 8678
rect 59028 8676 59034 8678
rect 58726 8667 59034 8676
rect 58726 7644 59034 7653
rect 58726 7642 58732 7644
rect 58788 7642 58812 7644
rect 58868 7642 58892 7644
rect 58948 7642 58972 7644
rect 59028 7642 59034 7644
rect 58788 7590 58790 7642
rect 58970 7590 58972 7642
rect 58726 7588 58732 7590
rect 58788 7588 58812 7590
rect 58868 7588 58892 7590
rect 58948 7588 58972 7590
rect 59028 7588 59034 7590
rect 58726 7579 59034 7588
rect 58726 6556 59034 6565
rect 58726 6554 58732 6556
rect 58788 6554 58812 6556
rect 58868 6554 58892 6556
rect 58948 6554 58972 6556
rect 59028 6554 59034 6556
rect 58788 6502 58790 6554
rect 58970 6502 58972 6554
rect 58726 6500 58732 6502
rect 58788 6500 58812 6502
rect 58868 6500 58892 6502
rect 58948 6500 58972 6502
rect 59028 6500 59034 6502
rect 58726 6491 59034 6500
rect 58440 5908 58492 5914
rect 58440 5850 58492 5856
rect 58726 5468 59034 5477
rect 58726 5466 58732 5468
rect 58788 5466 58812 5468
rect 58868 5466 58892 5468
rect 58948 5466 58972 5468
rect 59028 5466 59034 5468
rect 58788 5414 58790 5466
rect 58970 5414 58972 5466
rect 58726 5412 58732 5414
rect 58788 5412 58812 5414
rect 58868 5412 58892 5414
rect 58948 5412 58972 5414
rect 59028 5412 59034 5414
rect 58726 5403 59034 5412
rect 58726 4380 59034 4389
rect 58726 4378 58732 4380
rect 58788 4378 58812 4380
rect 58868 4378 58892 4380
rect 58948 4378 58972 4380
rect 59028 4378 59034 4380
rect 58788 4326 58790 4378
rect 58970 4326 58972 4378
rect 58726 4324 58732 4326
rect 58788 4324 58812 4326
rect 58868 4324 58892 4326
rect 58948 4324 58972 4326
rect 59028 4324 59034 4326
rect 58726 4315 59034 4324
rect 58532 3664 58584 3670
rect 58532 3606 58584 3612
rect 58348 2372 58400 2378
rect 58348 2314 58400 2320
rect 58268 870 58388 898
rect 58268 762 58296 870
rect 58360 800 58388 870
rect 58084 734 58296 762
rect 58346 0 58402 800
rect 58544 762 58572 3606
rect 58726 3292 59034 3301
rect 58726 3290 58732 3292
rect 58788 3290 58812 3292
rect 58868 3290 58892 3292
rect 58948 3290 58972 3292
rect 59028 3290 59034 3292
rect 58788 3238 58790 3290
rect 58970 3238 58972 3290
rect 58726 3236 58732 3238
rect 58788 3236 58812 3238
rect 58868 3236 58892 3238
rect 58948 3236 58972 3238
rect 59028 3236 59034 3238
rect 58726 3227 59034 3236
rect 58726 2204 59034 2213
rect 58726 2202 58732 2204
rect 58788 2202 58812 2204
rect 58868 2202 58892 2204
rect 58948 2202 58972 2204
rect 59028 2202 59034 2204
rect 58788 2150 58790 2202
rect 58970 2150 58972 2202
rect 58726 2148 58732 2150
rect 58788 2148 58812 2150
rect 58868 2148 58892 2150
rect 58948 2148 58972 2150
rect 59028 2148 59034 2150
rect 58726 2139 59034 2148
rect 58820 870 58940 898
rect 58820 762 58848 870
rect 58912 800 58940 870
rect 58544 734 58848 762
rect 58898 0 58954 800
<< via2 >>
rect 15400 21786 15456 21788
rect 15480 21786 15536 21788
rect 15560 21786 15616 21788
rect 15640 21786 15696 21788
rect 15400 21734 15446 21786
rect 15446 21734 15456 21786
rect 15480 21734 15510 21786
rect 15510 21734 15522 21786
rect 15522 21734 15536 21786
rect 15560 21734 15574 21786
rect 15574 21734 15586 21786
rect 15586 21734 15616 21786
rect 15640 21734 15650 21786
rect 15650 21734 15696 21786
rect 15400 21732 15456 21734
rect 15480 21732 15536 21734
rect 15560 21732 15616 21734
rect 15640 21732 15696 21734
rect 29844 21786 29900 21788
rect 29924 21786 29980 21788
rect 30004 21786 30060 21788
rect 30084 21786 30140 21788
rect 29844 21734 29890 21786
rect 29890 21734 29900 21786
rect 29924 21734 29954 21786
rect 29954 21734 29966 21786
rect 29966 21734 29980 21786
rect 30004 21734 30018 21786
rect 30018 21734 30030 21786
rect 30030 21734 30060 21786
rect 30084 21734 30094 21786
rect 30094 21734 30140 21786
rect 29844 21732 29900 21734
rect 29924 21732 29980 21734
rect 30004 21732 30060 21734
rect 30084 21732 30140 21734
rect 44288 21786 44344 21788
rect 44368 21786 44424 21788
rect 44448 21786 44504 21788
rect 44528 21786 44584 21788
rect 44288 21734 44334 21786
rect 44334 21734 44344 21786
rect 44368 21734 44398 21786
rect 44398 21734 44410 21786
rect 44410 21734 44424 21786
rect 44448 21734 44462 21786
rect 44462 21734 44474 21786
rect 44474 21734 44504 21786
rect 44528 21734 44538 21786
rect 44538 21734 44584 21786
rect 44288 21732 44344 21734
rect 44368 21732 44424 21734
rect 44448 21732 44504 21734
rect 44528 21732 44584 21734
rect 58732 21786 58788 21788
rect 58812 21786 58868 21788
rect 58892 21786 58948 21788
rect 58972 21786 59028 21788
rect 58732 21734 58778 21786
rect 58778 21734 58788 21786
rect 58812 21734 58842 21786
rect 58842 21734 58854 21786
rect 58854 21734 58868 21786
rect 58892 21734 58906 21786
rect 58906 21734 58918 21786
rect 58918 21734 58948 21786
rect 58972 21734 58982 21786
rect 58982 21734 59028 21786
rect 58732 21732 58788 21734
rect 58812 21732 58868 21734
rect 58892 21732 58948 21734
rect 58972 21732 59028 21734
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 938 3440 994 3496
rect 1674 3304 1730 3360
rect 1858 3188 1914 3224
rect 1858 3168 1860 3188
rect 1860 3168 1912 3188
rect 1912 3168 1914 3188
rect 2134 3596 2190 3632
rect 2134 3576 2136 3596
rect 2136 3576 2188 3596
rect 2188 3576 2190 3596
rect 3790 4020 3792 4040
rect 3792 4020 3844 4040
rect 3844 4020 3846 4040
rect 3790 3984 3846 4020
rect 4250 4428 4252 4448
rect 4252 4428 4304 4448
rect 4304 4428 4306 4448
rect 4250 4392 4306 4428
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 5170 5244 5172 5264
rect 5172 5244 5224 5264
rect 5224 5244 5226 5264
rect 5170 5208 5226 5244
rect 4710 3712 4766 3768
rect 4894 3596 4950 3632
rect 4894 3576 4896 3596
rect 4896 3576 4948 3596
rect 4948 3576 4950 3596
rect 6182 5480 6238 5536
rect 6182 5072 6238 5128
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 6734 3732 6790 3768
rect 6734 3712 6736 3732
rect 6736 3712 6788 3732
rect 6788 3712 6790 3732
rect 6642 3304 6698 3360
rect 7286 3576 7342 3632
rect 6918 3188 6974 3224
rect 6918 3168 6920 3188
rect 6920 3168 6972 3188
rect 6972 3168 6974 3188
rect 8114 7284 8116 7304
rect 8116 7284 8168 7304
rect 8168 7284 8170 7304
rect 8114 7248 8170 7284
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 9218 8900 9274 8936
rect 9218 8880 9220 8900
rect 9220 8880 9272 8900
rect 9272 8880 9274 8900
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8758 5208 8814 5264
rect 8850 5072 8906 5128
rect 9494 9424 9550 9480
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 9218 4392 9274 4448
rect 10138 9016 10194 9072
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 10598 4156 10600 4176
rect 10600 4156 10652 4176
rect 10652 4156 10654 4176
rect 10598 4120 10654 4156
rect 12990 10532 13046 10568
rect 12990 10512 12992 10532
rect 12992 10512 13044 10532
rect 13044 10512 13046 10532
rect 13358 8492 13414 8528
rect 13358 8472 13360 8492
rect 13360 8472 13412 8492
rect 13412 8472 13414 8492
rect 15400 20698 15456 20700
rect 15480 20698 15536 20700
rect 15560 20698 15616 20700
rect 15640 20698 15696 20700
rect 15400 20646 15446 20698
rect 15446 20646 15456 20698
rect 15480 20646 15510 20698
rect 15510 20646 15522 20698
rect 15522 20646 15536 20698
rect 15560 20646 15574 20698
rect 15574 20646 15586 20698
rect 15586 20646 15616 20698
rect 15640 20646 15650 20698
rect 15650 20646 15696 20698
rect 15400 20644 15456 20646
rect 15480 20644 15536 20646
rect 15560 20644 15616 20646
rect 15640 20644 15696 20646
rect 15400 19610 15456 19612
rect 15480 19610 15536 19612
rect 15560 19610 15616 19612
rect 15640 19610 15696 19612
rect 15400 19558 15446 19610
rect 15446 19558 15456 19610
rect 15480 19558 15510 19610
rect 15510 19558 15522 19610
rect 15522 19558 15536 19610
rect 15560 19558 15574 19610
rect 15574 19558 15586 19610
rect 15586 19558 15616 19610
rect 15640 19558 15650 19610
rect 15650 19558 15696 19610
rect 15400 19556 15456 19558
rect 15480 19556 15536 19558
rect 15560 19556 15616 19558
rect 15640 19556 15696 19558
rect 15400 18522 15456 18524
rect 15480 18522 15536 18524
rect 15560 18522 15616 18524
rect 15640 18522 15696 18524
rect 15400 18470 15446 18522
rect 15446 18470 15456 18522
rect 15480 18470 15510 18522
rect 15510 18470 15522 18522
rect 15522 18470 15536 18522
rect 15560 18470 15574 18522
rect 15574 18470 15586 18522
rect 15586 18470 15616 18522
rect 15640 18470 15650 18522
rect 15650 18470 15696 18522
rect 15400 18468 15456 18470
rect 15480 18468 15536 18470
rect 15560 18468 15616 18470
rect 15640 18468 15696 18470
rect 22622 21242 22678 21244
rect 22702 21242 22758 21244
rect 22782 21242 22838 21244
rect 22862 21242 22918 21244
rect 22622 21190 22668 21242
rect 22668 21190 22678 21242
rect 22702 21190 22732 21242
rect 22732 21190 22744 21242
rect 22744 21190 22758 21242
rect 22782 21190 22796 21242
rect 22796 21190 22808 21242
rect 22808 21190 22838 21242
rect 22862 21190 22872 21242
rect 22872 21190 22918 21242
rect 22622 21188 22678 21190
rect 22702 21188 22758 21190
rect 22782 21188 22838 21190
rect 22862 21188 22918 21190
rect 15400 17434 15456 17436
rect 15480 17434 15536 17436
rect 15560 17434 15616 17436
rect 15640 17434 15696 17436
rect 15400 17382 15446 17434
rect 15446 17382 15456 17434
rect 15480 17382 15510 17434
rect 15510 17382 15522 17434
rect 15522 17382 15536 17434
rect 15560 17382 15574 17434
rect 15574 17382 15586 17434
rect 15586 17382 15616 17434
rect 15640 17382 15650 17434
rect 15650 17382 15696 17434
rect 15400 17380 15456 17382
rect 15480 17380 15536 17382
rect 15560 17380 15616 17382
rect 15640 17380 15696 17382
rect 15400 16346 15456 16348
rect 15480 16346 15536 16348
rect 15560 16346 15616 16348
rect 15640 16346 15696 16348
rect 15400 16294 15446 16346
rect 15446 16294 15456 16346
rect 15480 16294 15510 16346
rect 15510 16294 15522 16346
rect 15522 16294 15536 16346
rect 15560 16294 15574 16346
rect 15574 16294 15586 16346
rect 15586 16294 15616 16346
rect 15640 16294 15650 16346
rect 15650 16294 15696 16346
rect 15400 16292 15456 16294
rect 15480 16292 15536 16294
rect 15560 16292 15616 16294
rect 15640 16292 15696 16294
rect 15400 15258 15456 15260
rect 15480 15258 15536 15260
rect 15560 15258 15616 15260
rect 15640 15258 15696 15260
rect 15400 15206 15446 15258
rect 15446 15206 15456 15258
rect 15480 15206 15510 15258
rect 15510 15206 15522 15258
rect 15522 15206 15536 15258
rect 15560 15206 15574 15258
rect 15574 15206 15586 15258
rect 15586 15206 15616 15258
rect 15640 15206 15650 15258
rect 15650 15206 15696 15258
rect 15400 15204 15456 15206
rect 15480 15204 15536 15206
rect 15560 15204 15616 15206
rect 15640 15204 15696 15206
rect 15400 14170 15456 14172
rect 15480 14170 15536 14172
rect 15560 14170 15616 14172
rect 15640 14170 15696 14172
rect 15400 14118 15446 14170
rect 15446 14118 15456 14170
rect 15480 14118 15510 14170
rect 15510 14118 15522 14170
rect 15522 14118 15536 14170
rect 15560 14118 15574 14170
rect 15574 14118 15586 14170
rect 15586 14118 15616 14170
rect 15640 14118 15650 14170
rect 15650 14118 15696 14170
rect 15400 14116 15456 14118
rect 15480 14116 15536 14118
rect 15560 14116 15616 14118
rect 15640 14116 15696 14118
rect 15400 13082 15456 13084
rect 15480 13082 15536 13084
rect 15560 13082 15616 13084
rect 15640 13082 15696 13084
rect 15400 13030 15446 13082
rect 15446 13030 15456 13082
rect 15480 13030 15510 13082
rect 15510 13030 15522 13082
rect 15522 13030 15536 13082
rect 15560 13030 15574 13082
rect 15574 13030 15586 13082
rect 15586 13030 15616 13082
rect 15640 13030 15650 13082
rect 15650 13030 15696 13082
rect 15400 13028 15456 13030
rect 15480 13028 15536 13030
rect 15560 13028 15616 13030
rect 15640 13028 15696 13030
rect 15400 11994 15456 11996
rect 15480 11994 15536 11996
rect 15560 11994 15616 11996
rect 15640 11994 15696 11996
rect 15400 11942 15446 11994
rect 15446 11942 15456 11994
rect 15480 11942 15510 11994
rect 15510 11942 15522 11994
rect 15522 11942 15536 11994
rect 15560 11942 15574 11994
rect 15574 11942 15586 11994
rect 15586 11942 15616 11994
rect 15640 11942 15650 11994
rect 15650 11942 15696 11994
rect 15400 11940 15456 11942
rect 15480 11940 15536 11942
rect 15560 11940 15616 11942
rect 15640 11940 15696 11942
rect 15400 10906 15456 10908
rect 15480 10906 15536 10908
rect 15560 10906 15616 10908
rect 15640 10906 15696 10908
rect 15400 10854 15446 10906
rect 15446 10854 15456 10906
rect 15480 10854 15510 10906
rect 15510 10854 15522 10906
rect 15522 10854 15536 10906
rect 15560 10854 15574 10906
rect 15574 10854 15586 10906
rect 15586 10854 15616 10906
rect 15640 10854 15650 10906
rect 15650 10854 15696 10906
rect 15400 10852 15456 10854
rect 15480 10852 15536 10854
rect 15560 10852 15616 10854
rect 15640 10852 15696 10854
rect 15400 9818 15456 9820
rect 15480 9818 15536 9820
rect 15560 9818 15616 9820
rect 15640 9818 15696 9820
rect 15400 9766 15446 9818
rect 15446 9766 15456 9818
rect 15480 9766 15510 9818
rect 15510 9766 15522 9818
rect 15522 9766 15536 9818
rect 15560 9766 15574 9818
rect 15574 9766 15586 9818
rect 15586 9766 15616 9818
rect 15640 9766 15650 9818
rect 15650 9766 15696 9818
rect 15400 9764 15456 9766
rect 15480 9764 15536 9766
rect 15560 9764 15616 9766
rect 15640 9764 15696 9766
rect 15290 9460 15292 9480
rect 15292 9460 15344 9480
rect 15344 9460 15346 9480
rect 15290 9424 15346 9460
rect 15400 8730 15456 8732
rect 15480 8730 15536 8732
rect 15560 8730 15616 8732
rect 15640 8730 15696 8732
rect 15400 8678 15446 8730
rect 15446 8678 15456 8730
rect 15480 8678 15510 8730
rect 15510 8678 15522 8730
rect 15522 8678 15536 8730
rect 15560 8678 15574 8730
rect 15574 8678 15586 8730
rect 15586 8678 15616 8730
rect 15640 8678 15650 8730
rect 15650 8678 15696 8730
rect 15400 8676 15456 8678
rect 15480 8676 15536 8678
rect 15560 8676 15616 8678
rect 15640 8676 15696 8678
rect 15400 7642 15456 7644
rect 15480 7642 15536 7644
rect 15560 7642 15616 7644
rect 15640 7642 15696 7644
rect 15400 7590 15446 7642
rect 15446 7590 15456 7642
rect 15480 7590 15510 7642
rect 15510 7590 15522 7642
rect 15522 7590 15536 7642
rect 15560 7590 15574 7642
rect 15574 7590 15586 7642
rect 15586 7590 15616 7642
rect 15640 7590 15650 7642
rect 15650 7590 15696 7642
rect 15400 7588 15456 7590
rect 15480 7588 15536 7590
rect 15560 7588 15616 7590
rect 15640 7588 15696 7590
rect 15400 6554 15456 6556
rect 15480 6554 15536 6556
rect 15560 6554 15616 6556
rect 15640 6554 15696 6556
rect 15400 6502 15446 6554
rect 15446 6502 15456 6554
rect 15480 6502 15510 6554
rect 15510 6502 15522 6554
rect 15522 6502 15536 6554
rect 15560 6502 15574 6554
rect 15574 6502 15586 6554
rect 15586 6502 15616 6554
rect 15640 6502 15650 6554
rect 15650 6502 15696 6554
rect 15400 6500 15456 6502
rect 15480 6500 15536 6502
rect 15560 6500 15616 6502
rect 15640 6500 15696 6502
rect 15400 5466 15456 5468
rect 15480 5466 15536 5468
rect 15560 5466 15616 5468
rect 15640 5466 15696 5468
rect 15400 5414 15446 5466
rect 15446 5414 15456 5466
rect 15480 5414 15510 5466
rect 15510 5414 15522 5466
rect 15522 5414 15536 5466
rect 15560 5414 15574 5466
rect 15574 5414 15586 5466
rect 15586 5414 15616 5466
rect 15640 5414 15650 5466
rect 15650 5414 15696 5466
rect 15400 5412 15456 5414
rect 15480 5412 15536 5414
rect 15560 5412 15616 5414
rect 15640 5412 15696 5414
rect 15400 4378 15456 4380
rect 15480 4378 15536 4380
rect 15560 4378 15616 4380
rect 15640 4378 15696 4380
rect 15400 4326 15446 4378
rect 15446 4326 15456 4378
rect 15480 4326 15510 4378
rect 15510 4326 15522 4378
rect 15522 4326 15536 4378
rect 15560 4326 15574 4378
rect 15574 4326 15586 4378
rect 15586 4326 15616 4378
rect 15640 4326 15650 4378
rect 15650 4326 15696 4378
rect 15400 4324 15456 4326
rect 15480 4324 15536 4326
rect 15560 4324 15616 4326
rect 15640 4324 15696 4326
rect 15400 3290 15456 3292
rect 15480 3290 15536 3292
rect 15560 3290 15616 3292
rect 15640 3290 15696 3292
rect 15400 3238 15446 3290
rect 15446 3238 15456 3290
rect 15480 3238 15510 3290
rect 15510 3238 15522 3290
rect 15522 3238 15536 3290
rect 15560 3238 15574 3290
rect 15574 3238 15586 3290
rect 15586 3238 15616 3290
rect 15640 3238 15650 3290
rect 15650 3238 15696 3290
rect 15400 3236 15456 3238
rect 15480 3236 15536 3238
rect 15560 3236 15616 3238
rect 15640 3236 15696 3238
rect 16026 3340 16028 3360
rect 16028 3340 16080 3360
rect 16080 3340 16082 3360
rect 16026 3304 16082 3340
rect 15400 2202 15456 2204
rect 15480 2202 15536 2204
rect 15560 2202 15616 2204
rect 15640 2202 15696 2204
rect 15400 2150 15446 2202
rect 15446 2150 15456 2202
rect 15480 2150 15510 2202
rect 15510 2150 15522 2202
rect 15522 2150 15536 2202
rect 15560 2150 15574 2202
rect 15574 2150 15586 2202
rect 15586 2150 15616 2202
rect 15640 2150 15650 2202
rect 15650 2150 15696 2202
rect 15400 2148 15456 2150
rect 15480 2148 15536 2150
rect 15560 2148 15616 2150
rect 15640 2148 15696 2150
rect 19982 10668 20038 10704
rect 19982 10648 19984 10668
rect 19984 10648 20036 10668
rect 20036 10648 20038 10668
rect 22622 20154 22678 20156
rect 22702 20154 22758 20156
rect 22782 20154 22838 20156
rect 22862 20154 22918 20156
rect 22622 20102 22668 20154
rect 22668 20102 22678 20154
rect 22702 20102 22732 20154
rect 22732 20102 22744 20154
rect 22744 20102 22758 20154
rect 22782 20102 22796 20154
rect 22796 20102 22808 20154
rect 22808 20102 22838 20154
rect 22862 20102 22872 20154
rect 22872 20102 22918 20154
rect 22622 20100 22678 20102
rect 22702 20100 22758 20102
rect 22782 20100 22838 20102
rect 22862 20100 22918 20102
rect 22622 19066 22678 19068
rect 22702 19066 22758 19068
rect 22782 19066 22838 19068
rect 22862 19066 22918 19068
rect 22622 19014 22668 19066
rect 22668 19014 22678 19066
rect 22702 19014 22732 19066
rect 22732 19014 22744 19066
rect 22744 19014 22758 19066
rect 22782 19014 22796 19066
rect 22796 19014 22808 19066
rect 22808 19014 22838 19066
rect 22862 19014 22872 19066
rect 22872 19014 22918 19066
rect 22622 19012 22678 19014
rect 22702 19012 22758 19014
rect 22782 19012 22838 19014
rect 22862 19012 22918 19014
rect 22622 17978 22678 17980
rect 22702 17978 22758 17980
rect 22782 17978 22838 17980
rect 22862 17978 22918 17980
rect 22622 17926 22668 17978
rect 22668 17926 22678 17978
rect 22702 17926 22732 17978
rect 22732 17926 22744 17978
rect 22744 17926 22758 17978
rect 22782 17926 22796 17978
rect 22796 17926 22808 17978
rect 22808 17926 22838 17978
rect 22862 17926 22872 17978
rect 22872 17926 22918 17978
rect 22622 17924 22678 17926
rect 22702 17924 22758 17926
rect 22782 17924 22838 17926
rect 22862 17924 22918 17926
rect 22622 16890 22678 16892
rect 22702 16890 22758 16892
rect 22782 16890 22838 16892
rect 22862 16890 22918 16892
rect 22622 16838 22668 16890
rect 22668 16838 22678 16890
rect 22702 16838 22732 16890
rect 22732 16838 22744 16890
rect 22744 16838 22758 16890
rect 22782 16838 22796 16890
rect 22796 16838 22808 16890
rect 22808 16838 22838 16890
rect 22862 16838 22872 16890
rect 22872 16838 22918 16890
rect 22622 16836 22678 16838
rect 22702 16836 22758 16838
rect 22782 16836 22838 16838
rect 22862 16836 22918 16838
rect 22622 15802 22678 15804
rect 22702 15802 22758 15804
rect 22782 15802 22838 15804
rect 22862 15802 22918 15804
rect 22622 15750 22668 15802
rect 22668 15750 22678 15802
rect 22702 15750 22732 15802
rect 22732 15750 22744 15802
rect 22744 15750 22758 15802
rect 22782 15750 22796 15802
rect 22796 15750 22808 15802
rect 22808 15750 22838 15802
rect 22862 15750 22872 15802
rect 22872 15750 22918 15802
rect 22622 15748 22678 15750
rect 22702 15748 22758 15750
rect 22782 15748 22838 15750
rect 22862 15748 22918 15750
rect 22622 14714 22678 14716
rect 22702 14714 22758 14716
rect 22782 14714 22838 14716
rect 22862 14714 22918 14716
rect 22622 14662 22668 14714
rect 22668 14662 22678 14714
rect 22702 14662 22732 14714
rect 22732 14662 22744 14714
rect 22744 14662 22758 14714
rect 22782 14662 22796 14714
rect 22796 14662 22808 14714
rect 22808 14662 22838 14714
rect 22862 14662 22872 14714
rect 22872 14662 22918 14714
rect 22622 14660 22678 14662
rect 22702 14660 22758 14662
rect 22782 14660 22838 14662
rect 22862 14660 22918 14662
rect 22622 13626 22678 13628
rect 22702 13626 22758 13628
rect 22782 13626 22838 13628
rect 22862 13626 22918 13628
rect 22622 13574 22668 13626
rect 22668 13574 22678 13626
rect 22702 13574 22732 13626
rect 22732 13574 22744 13626
rect 22744 13574 22758 13626
rect 22782 13574 22796 13626
rect 22796 13574 22808 13626
rect 22808 13574 22838 13626
rect 22862 13574 22872 13626
rect 22872 13574 22918 13626
rect 22622 13572 22678 13574
rect 22702 13572 22758 13574
rect 22782 13572 22838 13574
rect 22862 13572 22918 13574
rect 22622 12538 22678 12540
rect 22702 12538 22758 12540
rect 22782 12538 22838 12540
rect 22862 12538 22918 12540
rect 22622 12486 22668 12538
rect 22668 12486 22678 12538
rect 22702 12486 22732 12538
rect 22732 12486 22744 12538
rect 22744 12486 22758 12538
rect 22782 12486 22796 12538
rect 22796 12486 22808 12538
rect 22808 12486 22838 12538
rect 22862 12486 22872 12538
rect 22872 12486 22918 12538
rect 22622 12484 22678 12486
rect 22702 12484 22758 12486
rect 22782 12484 22838 12486
rect 22862 12484 22918 12486
rect 22622 11450 22678 11452
rect 22702 11450 22758 11452
rect 22782 11450 22838 11452
rect 22862 11450 22918 11452
rect 22622 11398 22668 11450
rect 22668 11398 22678 11450
rect 22702 11398 22732 11450
rect 22732 11398 22744 11450
rect 22744 11398 22758 11450
rect 22782 11398 22796 11450
rect 22796 11398 22808 11450
rect 22808 11398 22838 11450
rect 22862 11398 22872 11450
rect 22872 11398 22918 11450
rect 22622 11396 22678 11398
rect 22702 11396 22758 11398
rect 22782 11396 22838 11398
rect 22862 11396 22918 11398
rect 22622 10362 22678 10364
rect 22702 10362 22758 10364
rect 22782 10362 22838 10364
rect 22862 10362 22918 10364
rect 22622 10310 22668 10362
rect 22668 10310 22678 10362
rect 22702 10310 22732 10362
rect 22732 10310 22744 10362
rect 22744 10310 22758 10362
rect 22782 10310 22796 10362
rect 22796 10310 22808 10362
rect 22808 10310 22838 10362
rect 22862 10310 22872 10362
rect 22872 10310 22918 10362
rect 22622 10308 22678 10310
rect 22702 10308 22758 10310
rect 22782 10308 22838 10310
rect 22862 10308 22918 10310
rect 22006 9832 22062 9888
rect 24674 20440 24730 20496
rect 22190 9832 22246 9888
rect 22622 9274 22678 9276
rect 22702 9274 22758 9276
rect 22782 9274 22838 9276
rect 22862 9274 22918 9276
rect 22622 9222 22668 9274
rect 22668 9222 22678 9274
rect 22702 9222 22732 9274
rect 22732 9222 22744 9274
rect 22744 9222 22758 9274
rect 22782 9222 22796 9274
rect 22796 9222 22808 9274
rect 22808 9222 22838 9274
rect 22862 9222 22872 9274
rect 22872 9222 22918 9274
rect 22622 9220 22678 9222
rect 22702 9220 22758 9222
rect 22782 9220 22838 9222
rect 22862 9220 22918 9222
rect 22622 8186 22678 8188
rect 22702 8186 22758 8188
rect 22782 8186 22838 8188
rect 22862 8186 22918 8188
rect 22622 8134 22668 8186
rect 22668 8134 22678 8186
rect 22702 8134 22732 8186
rect 22732 8134 22744 8186
rect 22744 8134 22758 8186
rect 22782 8134 22796 8186
rect 22796 8134 22808 8186
rect 22808 8134 22838 8186
rect 22862 8134 22872 8186
rect 22872 8134 22918 8186
rect 22622 8132 22678 8134
rect 22702 8132 22758 8134
rect 22782 8132 22838 8134
rect 22862 8132 22918 8134
rect 22622 7098 22678 7100
rect 22702 7098 22758 7100
rect 22782 7098 22838 7100
rect 22862 7098 22918 7100
rect 22622 7046 22668 7098
rect 22668 7046 22678 7098
rect 22702 7046 22732 7098
rect 22732 7046 22744 7098
rect 22744 7046 22758 7098
rect 22782 7046 22796 7098
rect 22796 7046 22808 7098
rect 22808 7046 22838 7098
rect 22862 7046 22872 7098
rect 22872 7046 22918 7098
rect 22622 7044 22678 7046
rect 22702 7044 22758 7046
rect 22782 7044 22838 7046
rect 22862 7044 22918 7046
rect 22622 6010 22678 6012
rect 22702 6010 22758 6012
rect 22782 6010 22838 6012
rect 22862 6010 22918 6012
rect 22622 5958 22668 6010
rect 22668 5958 22678 6010
rect 22702 5958 22732 6010
rect 22732 5958 22744 6010
rect 22744 5958 22758 6010
rect 22782 5958 22796 6010
rect 22796 5958 22808 6010
rect 22808 5958 22838 6010
rect 22862 5958 22872 6010
rect 22872 5958 22918 6010
rect 22622 5956 22678 5958
rect 22702 5956 22758 5958
rect 22782 5956 22838 5958
rect 22862 5956 22918 5958
rect 22622 4922 22678 4924
rect 22702 4922 22758 4924
rect 22782 4922 22838 4924
rect 22862 4922 22918 4924
rect 22622 4870 22668 4922
rect 22668 4870 22678 4922
rect 22702 4870 22732 4922
rect 22732 4870 22744 4922
rect 22744 4870 22758 4922
rect 22782 4870 22796 4922
rect 22796 4870 22808 4922
rect 22808 4870 22838 4922
rect 22862 4870 22872 4922
rect 22872 4870 22918 4922
rect 22622 4868 22678 4870
rect 22702 4868 22758 4870
rect 22782 4868 22838 4870
rect 22862 4868 22918 4870
rect 22622 3834 22678 3836
rect 22702 3834 22758 3836
rect 22782 3834 22838 3836
rect 22862 3834 22918 3836
rect 22622 3782 22668 3834
rect 22668 3782 22678 3834
rect 22702 3782 22732 3834
rect 22732 3782 22744 3834
rect 22744 3782 22758 3834
rect 22782 3782 22796 3834
rect 22796 3782 22808 3834
rect 22808 3782 22838 3834
rect 22862 3782 22872 3834
rect 22872 3782 22918 3834
rect 22622 3780 22678 3782
rect 22702 3780 22758 3782
rect 22782 3780 22838 3782
rect 22862 3780 22918 3782
rect 22622 2746 22678 2748
rect 22702 2746 22758 2748
rect 22782 2746 22838 2748
rect 22862 2746 22918 2748
rect 22622 2694 22668 2746
rect 22668 2694 22678 2746
rect 22702 2694 22732 2746
rect 22732 2694 22744 2746
rect 22744 2694 22758 2746
rect 22782 2694 22796 2746
rect 22796 2694 22808 2746
rect 22808 2694 22838 2746
rect 22862 2694 22872 2746
rect 22872 2694 22918 2746
rect 22622 2692 22678 2694
rect 22702 2692 22758 2694
rect 22782 2692 22838 2694
rect 22862 2692 22918 2694
rect 29844 20698 29900 20700
rect 29924 20698 29980 20700
rect 30004 20698 30060 20700
rect 30084 20698 30140 20700
rect 29844 20646 29890 20698
rect 29890 20646 29900 20698
rect 29924 20646 29954 20698
rect 29954 20646 29966 20698
rect 29966 20646 29980 20698
rect 30004 20646 30018 20698
rect 30018 20646 30030 20698
rect 30030 20646 30060 20698
rect 30084 20646 30094 20698
rect 30094 20646 30140 20698
rect 29844 20644 29900 20646
rect 29924 20644 29980 20646
rect 30004 20644 30060 20646
rect 30084 20644 30140 20646
rect 29844 19610 29900 19612
rect 29924 19610 29980 19612
rect 30004 19610 30060 19612
rect 30084 19610 30140 19612
rect 29844 19558 29890 19610
rect 29890 19558 29900 19610
rect 29924 19558 29954 19610
rect 29954 19558 29966 19610
rect 29966 19558 29980 19610
rect 30004 19558 30018 19610
rect 30018 19558 30030 19610
rect 30030 19558 30060 19610
rect 30084 19558 30094 19610
rect 30094 19558 30140 19610
rect 29844 19556 29900 19558
rect 29924 19556 29980 19558
rect 30004 19556 30060 19558
rect 30084 19556 30140 19558
rect 29844 18522 29900 18524
rect 29924 18522 29980 18524
rect 30004 18522 30060 18524
rect 30084 18522 30140 18524
rect 29844 18470 29890 18522
rect 29890 18470 29900 18522
rect 29924 18470 29954 18522
rect 29954 18470 29966 18522
rect 29966 18470 29980 18522
rect 30004 18470 30018 18522
rect 30018 18470 30030 18522
rect 30030 18470 30060 18522
rect 30084 18470 30094 18522
rect 30094 18470 30140 18522
rect 29844 18468 29900 18470
rect 29924 18468 29980 18470
rect 30004 18468 30060 18470
rect 30084 18468 30140 18470
rect 27710 9868 27712 9888
rect 27712 9868 27764 9888
rect 27764 9868 27766 9888
rect 27710 9832 27766 9868
rect 29844 17434 29900 17436
rect 29924 17434 29980 17436
rect 30004 17434 30060 17436
rect 30084 17434 30140 17436
rect 29844 17382 29890 17434
rect 29890 17382 29900 17434
rect 29924 17382 29954 17434
rect 29954 17382 29966 17434
rect 29966 17382 29980 17434
rect 30004 17382 30018 17434
rect 30018 17382 30030 17434
rect 30030 17382 30060 17434
rect 30084 17382 30094 17434
rect 30094 17382 30140 17434
rect 29844 17380 29900 17382
rect 29924 17380 29980 17382
rect 30004 17380 30060 17382
rect 30084 17380 30140 17382
rect 29844 16346 29900 16348
rect 29924 16346 29980 16348
rect 30004 16346 30060 16348
rect 30084 16346 30140 16348
rect 29844 16294 29890 16346
rect 29890 16294 29900 16346
rect 29924 16294 29954 16346
rect 29954 16294 29966 16346
rect 29966 16294 29980 16346
rect 30004 16294 30018 16346
rect 30018 16294 30030 16346
rect 30030 16294 30060 16346
rect 30084 16294 30094 16346
rect 30094 16294 30140 16346
rect 29844 16292 29900 16294
rect 29924 16292 29980 16294
rect 30004 16292 30060 16294
rect 30084 16292 30140 16294
rect 29844 15258 29900 15260
rect 29924 15258 29980 15260
rect 30004 15258 30060 15260
rect 30084 15258 30140 15260
rect 29844 15206 29890 15258
rect 29890 15206 29900 15258
rect 29924 15206 29954 15258
rect 29954 15206 29966 15258
rect 29966 15206 29980 15258
rect 30004 15206 30018 15258
rect 30018 15206 30030 15258
rect 30030 15206 30060 15258
rect 30084 15206 30094 15258
rect 30094 15206 30140 15258
rect 29844 15204 29900 15206
rect 29924 15204 29980 15206
rect 30004 15204 30060 15206
rect 30084 15204 30140 15206
rect 29844 14170 29900 14172
rect 29924 14170 29980 14172
rect 30004 14170 30060 14172
rect 30084 14170 30140 14172
rect 29844 14118 29890 14170
rect 29890 14118 29900 14170
rect 29924 14118 29954 14170
rect 29954 14118 29966 14170
rect 29966 14118 29980 14170
rect 30004 14118 30018 14170
rect 30018 14118 30030 14170
rect 30030 14118 30060 14170
rect 30084 14118 30094 14170
rect 30094 14118 30140 14170
rect 29844 14116 29900 14118
rect 29924 14116 29980 14118
rect 30004 14116 30060 14118
rect 30084 14116 30140 14118
rect 29844 13082 29900 13084
rect 29924 13082 29980 13084
rect 30004 13082 30060 13084
rect 30084 13082 30140 13084
rect 29844 13030 29890 13082
rect 29890 13030 29900 13082
rect 29924 13030 29954 13082
rect 29954 13030 29966 13082
rect 29966 13030 29980 13082
rect 30004 13030 30018 13082
rect 30018 13030 30030 13082
rect 30030 13030 30060 13082
rect 30084 13030 30094 13082
rect 30094 13030 30140 13082
rect 29844 13028 29900 13030
rect 29924 13028 29980 13030
rect 30004 13028 30060 13030
rect 30084 13028 30140 13030
rect 27342 3304 27398 3360
rect 27802 2896 27858 2952
rect 29844 11994 29900 11996
rect 29924 11994 29980 11996
rect 30004 11994 30060 11996
rect 30084 11994 30140 11996
rect 29844 11942 29890 11994
rect 29890 11942 29900 11994
rect 29924 11942 29954 11994
rect 29954 11942 29966 11994
rect 29966 11942 29980 11994
rect 30004 11942 30018 11994
rect 30018 11942 30030 11994
rect 30030 11942 30060 11994
rect 30084 11942 30094 11994
rect 30094 11942 30140 11994
rect 29844 11940 29900 11942
rect 29924 11940 29980 11942
rect 30004 11940 30060 11942
rect 30084 11940 30140 11942
rect 29844 10906 29900 10908
rect 29924 10906 29980 10908
rect 30004 10906 30060 10908
rect 30084 10906 30140 10908
rect 29844 10854 29890 10906
rect 29890 10854 29900 10906
rect 29924 10854 29954 10906
rect 29954 10854 29966 10906
rect 29966 10854 29980 10906
rect 30004 10854 30018 10906
rect 30018 10854 30030 10906
rect 30030 10854 30060 10906
rect 30084 10854 30094 10906
rect 30094 10854 30140 10906
rect 29844 10852 29900 10854
rect 29924 10852 29980 10854
rect 30004 10852 30060 10854
rect 30084 10852 30140 10854
rect 29844 9818 29900 9820
rect 29924 9818 29980 9820
rect 30004 9818 30060 9820
rect 30084 9818 30140 9820
rect 29844 9766 29890 9818
rect 29890 9766 29900 9818
rect 29924 9766 29954 9818
rect 29954 9766 29966 9818
rect 29966 9766 29980 9818
rect 30004 9766 30018 9818
rect 30018 9766 30030 9818
rect 30030 9766 30060 9818
rect 30084 9766 30094 9818
rect 30094 9766 30140 9818
rect 29844 9764 29900 9766
rect 29924 9764 29980 9766
rect 30004 9764 30060 9766
rect 30084 9764 30140 9766
rect 31114 12960 31170 13016
rect 37066 21242 37122 21244
rect 37146 21242 37202 21244
rect 37226 21242 37282 21244
rect 37306 21242 37362 21244
rect 37066 21190 37112 21242
rect 37112 21190 37122 21242
rect 37146 21190 37176 21242
rect 37176 21190 37188 21242
rect 37188 21190 37202 21242
rect 37226 21190 37240 21242
rect 37240 21190 37252 21242
rect 37252 21190 37282 21242
rect 37306 21190 37316 21242
rect 37316 21190 37362 21242
rect 37066 21188 37122 21190
rect 37146 21188 37202 21190
rect 37226 21188 37282 21190
rect 37306 21188 37362 21190
rect 30654 10648 30710 10704
rect 29844 8730 29900 8732
rect 29924 8730 29980 8732
rect 30004 8730 30060 8732
rect 30084 8730 30140 8732
rect 29844 8678 29890 8730
rect 29890 8678 29900 8730
rect 29924 8678 29954 8730
rect 29954 8678 29966 8730
rect 29966 8678 29980 8730
rect 30004 8678 30018 8730
rect 30018 8678 30030 8730
rect 30030 8678 30060 8730
rect 30084 8678 30094 8730
rect 30094 8678 30140 8730
rect 29844 8676 29900 8678
rect 29924 8676 29980 8678
rect 30004 8676 30060 8678
rect 30084 8676 30140 8678
rect 29844 7642 29900 7644
rect 29924 7642 29980 7644
rect 30004 7642 30060 7644
rect 30084 7642 30140 7644
rect 29844 7590 29890 7642
rect 29890 7590 29900 7642
rect 29924 7590 29954 7642
rect 29954 7590 29966 7642
rect 29966 7590 29980 7642
rect 30004 7590 30018 7642
rect 30018 7590 30030 7642
rect 30030 7590 30060 7642
rect 30084 7590 30094 7642
rect 30094 7590 30140 7642
rect 29844 7588 29900 7590
rect 29924 7588 29980 7590
rect 30004 7588 30060 7590
rect 30084 7588 30140 7590
rect 29550 3440 29606 3496
rect 30746 9424 30802 9480
rect 30194 6876 30196 6896
rect 30196 6876 30248 6896
rect 30248 6876 30250 6896
rect 30194 6840 30250 6876
rect 29844 6554 29900 6556
rect 29924 6554 29980 6556
rect 30004 6554 30060 6556
rect 30084 6554 30140 6556
rect 29844 6502 29890 6554
rect 29890 6502 29900 6554
rect 29924 6502 29954 6554
rect 29954 6502 29966 6554
rect 29966 6502 29980 6554
rect 30004 6502 30018 6554
rect 30018 6502 30030 6554
rect 30030 6502 30060 6554
rect 30084 6502 30094 6554
rect 30094 6502 30140 6554
rect 29844 6500 29900 6502
rect 29924 6500 29980 6502
rect 30004 6500 30060 6502
rect 30084 6500 30140 6502
rect 29844 5466 29900 5468
rect 29924 5466 29980 5468
rect 30004 5466 30060 5468
rect 30084 5466 30140 5468
rect 29844 5414 29890 5466
rect 29890 5414 29900 5466
rect 29924 5414 29954 5466
rect 29954 5414 29966 5466
rect 29966 5414 29980 5466
rect 30004 5414 30018 5466
rect 30018 5414 30030 5466
rect 30030 5414 30060 5466
rect 30084 5414 30094 5466
rect 30094 5414 30140 5466
rect 29844 5412 29900 5414
rect 29924 5412 29980 5414
rect 30004 5412 30060 5414
rect 30084 5412 30140 5414
rect 31298 6840 31354 6896
rect 29844 4378 29900 4380
rect 29924 4378 29980 4380
rect 30004 4378 30060 4380
rect 30084 4378 30140 4380
rect 29844 4326 29890 4378
rect 29890 4326 29900 4378
rect 29924 4326 29954 4378
rect 29954 4326 29966 4378
rect 29966 4326 29980 4378
rect 30004 4326 30018 4378
rect 30018 4326 30030 4378
rect 30030 4326 30060 4378
rect 30084 4326 30094 4378
rect 30094 4326 30140 4378
rect 29844 4324 29900 4326
rect 29924 4324 29980 4326
rect 30004 4324 30060 4326
rect 30084 4324 30140 4326
rect 30378 4120 30434 4176
rect 31482 5208 31538 5264
rect 29844 3290 29900 3292
rect 29924 3290 29980 3292
rect 30004 3290 30060 3292
rect 30084 3290 30140 3292
rect 29844 3238 29890 3290
rect 29890 3238 29900 3290
rect 29924 3238 29954 3290
rect 29954 3238 29966 3290
rect 29966 3238 29980 3290
rect 30004 3238 30018 3290
rect 30018 3238 30030 3290
rect 30030 3238 30060 3290
rect 30084 3238 30094 3290
rect 30094 3238 30140 3290
rect 29844 3236 29900 3238
rect 29924 3236 29980 3238
rect 30004 3236 30060 3238
rect 30084 3236 30140 3238
rect 30286 3984 30342 4040
rect 29844 2202 29900 2204
rect 29924 2202 29980 2204
rect 30004 2202 30060 2204
rect 30084 2202 30140 2204
rect 29844 2150 29890 2202
rect 29890 2150 29900 2202
rect 29924 2150 29954 2202
rect 29954 2150 29966 2202
rect 29966 2150 29980 2202
rect 30004 2150 30018 2202
rect 30018 2150 30030 2202
rect 30030 2150 30060 2202
rect 30084 2150 30094 2202
rect 30094 2150 30140 2202
rect 29844 2148 29900 2150
rect 29924 2148 29980 2150
rect 30004 2148 30060 2150
rect 30084 2148 30140 2150
rect 32310 4936 32366 4992
rect 32770 4936 32826 4992
rect 33230 4140 33286 4176
rect 33230 4120 33232 4140
rect 33232 4120 33284 4140
rect 33284 4120 33286 4140
rect 37066 20154 37122 20156
rect 37146 20154 37202 20156
rect 37226 20154 37282 20156
rect 37306 20154 37362 20156
rect 37066 20102 37112 20154
rect 37112 20102 37122 20154
rect 37146 20102 37176 20154
rect 37176 20102 37188 20154
rect 37188 20102 37202 20154
rect 37226 20102 37240 20154
rect 37240 20102 37252 20154
rect 37252 20102 37282 20154
rect 37306 20102 37316 20154
rect 37316 20102 37362 20154
rect 37066 20100 37122 20102
rect 37146 20100 37202 20102
rect 37226 20100 37282 20102
rect 37306 20100 37362 20102
rect 37066 19066 37122 19068
rect 37146 19066 37202 19068
rect 37226 19066 37282 19068
rect 37306 19066 37362 19068
rect 37066 19014 37112 19066
rect 37112 19014 37122 19066
rect 37146 19014 37176 19066
rect 37176 19014 37188 19066
rect 37188 19014 37202 19066
rect 37226 19014 37240 19066
rect 37240 19014 37252 19066
rect 37252 19014 37282 19066
rect 37306 19014 37316 19066
rect 37316 19014 37362 19066
rect 37066 19012 37122 19014
rect 37146 19012 37202 19014
rect 37226 19012 37282 19014
rect 37306 19012 37362 19014
rect 35438 16632 35494 16688
rect 35806 13404 35808 13424
rect 35808 13404 35860 13424
rect 35860 13404 35862 13424
rect 35530 12724 35532 12744
rect 35532 12724 35584 12744
rect 35584 12724 35586 12744
rect 35530 12688 35586 12724
rect 34978 6876 34980 6896
rect 34980 6876 35032 6896
rect 35032 6876 35034 6896
rect 34978 6840 35034 6876
rect 34886 5244 34888 5264
rect 34888 5244 34940 5264
rect 34940 5244 34942 5264
rect 34886 5208 34942 5244
rect 35162 4548 35218 4584
rect 35162 4528 35164 4548
rect 35164 4528 35216 4548
rect 35216 4528 35218 4548
rect 35806 13368 35862 13404
rect 37066 17978 37122 17980
rect 37146 17978 37202 17980
rect 37226 17978 37282 17980
rect 37306 17978 37362 17980
rect 37066 17926 37112 17978
rect 37112 17926 37122 17978
rect 37146 17926 37176 17978
rect 37176 17926 37188 17978
rect 37188 17926 37202 17978
rect 37226 17926 37240 17978
rect 37240 17926 37252 17978
rect 37252 17926 37282 17978
rect 37306 17926 37316 17978
rect 37316 17926 37362 17978
rect 37066 17924 37122 17926
rect 37146 17924 37202 17926
rect 37226 17924 37282 17926
rect 37306 17924 37362 17926
rect 37066 16890 37122 16892
rect 37146 16890 37202 16892
rect 37226 16890 37282 16892
rect 37306 16890 37362 16892
rect 37066 16838 37112 16890
rect 37112 16838 37122 16890
rect 37146 16838 37176 16890
rect 37176 16838 37188 16890
rect 37188 16838 37202 16890
rect 37226 16838 37240 16890
rect 37240 16838 37252 16890
rect 37252 16838 37282 16890
rect 37306 16838 37316 16890
rect 37316 16838 37362 16890
rect 37066 16836 37122 16838
rect 37146 16836 37202 16838
rect 37226 16836 37282 16838
rect 37306 16836 37362 16838
rect 37066 15802 37122 15804
rect 37146 15802 37202 15804
rect 37226 15802 37282 15804
rect 37306 15802 37362 15804
rect 37066 15750 37112 15802
rect 37112 15750 37122 15802
rect 37146 15750 37176 15802
rect 37176 15750 37188 15802
rect 37188 15750 37202 15802
rect 37226 15750 37240 15802
rect 37240 15750 37252 15802
rect 37252 15750 37282 15802
rect 37306 15750 37316 15802
rect 37316 15750 37362 15802
rect 37066 15748 37122 15750
rect 37146 15748 37202 15750
rect 37226 15748 37282 15750
rect 37306 15748 37362 15750
rect 35714 7384 35770 7440
rect 37066 14714 37122 14716
rect 37146 14714 37202 14716
rect 37226 14714 37282 14716
rect 37306 14714 37362 14716
rect 37066 14662 37112 14714
rect 37112 14662 37122 14714
rect 37146 14662 37176 14714
rect 37176 14662 37188 14714
rect 37188 14662 37202 14714
rect 37226 14662 37240 14714
rect 37240 14662 37252 14714
rect 37252 14662 37282 14714
rect 37306 14662 37316 14714
rect 37316 14662 37362 14714
rect 37066 14660 37122 14662
rect 37146 14660 37202 14662
rect 37226 14660 37282 14662
rect 37306 14660 37362 14662
rect 37066 13626 37122 13628
rect 37146 13626 37202 13628
rect 37226 13626 37282 13628
rect 37306 13626 37362 13628
rect 37066 13574 37112 13626
rect 37112 13574 37122 13626
rect 37146 13574 37176 13626
rect 37176 13574 37188 13626
rect 37188 13574 37202 13626
rect 37226 13574 37240 13626
rect 37240 13574 37252 13626
rect 37252 13574 37282 13626
rect 37306 13574 37316 13626
rect 37316 13574 37362 13626
rect 37066 13572 37122 13574
rect 37146 13572 37202 13574
rect 37226 13572 37282 13574
rect 37306 13572 37362 13574
rect 37066 12538 37122 12540
rect 37146 12538 37202 12540
rect 37226 12538 37282 12540
rect 37306 12538 37362 12540
rect 37066 12486 37112 12538
rect 37112 12486 37122 12538
rect 37146 12486 37176 12538
rect 37176 12486 37188 12538
rect 37188 12486 37202 12538
rect 37226 12486 37240 12538
rect 37240 12486 37252 12538
rect 37252 12486 37282 12538
rect 37306 12486 37316 12538
rect 37316 12486 37362 12538
rect 37066 12484 37122 12486
rect 37146 12484 37202 12486
rect 37226 12484 37282 12486
rect 37306 12484 37362 12486
rect 40038 19760 40094 19816
rect 37066 11450 37122 11452
rect 37146 11450 37202 11452
rect 37226 11450 37282 11452
rect 37306 11450 37362 11452
rect 37066 11398 37112 11450
rect 37112 11398 37122 11450
rect 37146 11398 37176 11450
rect 37176 11398 37188 11450
rect 37188 11398 37202 11450
rect 37226 11398 37240 11450
rect 37240 11398 37252 11450
rect 37252 11398 37282 11450
rect 37306 11398 37316 11450
rect 37316 11398 37362 11450
rect 37066 11396 37122 11398
rect 37146 11396 37202 11398
rect 37226 11396 37282 11398
rect 37306 11396 37362 11398
rect 37066 10362 37122 10364
rect 37146 10362 37202 10364
rect 37226 10362 37282 10364
rect 37306 10362 37362 10364
rect 37066 10310 37112 10362
rect 37112 10310 37122 10362
rect 37146 10310 37176 10362
rect 37176 10310 37188 10362
rect 37188 10310 37202 10362
rect 37226 10310 37240 10362
rect 37240 10310 37252 10362
rect 37252 10310 37282 10362
rect 37306 10310 37316 10362
rect 37316 10310 37362 10362
rect 37066 10308 37122 10310
rect 37146 10308 37202 10310
rect 37226 10308 37282 10310
rect 37306 10308 37362 10310
rect 35346 4020 35348 4040
rect 35348 4020 35400 4040
rect 35400 4020 35402 4040
rect 35346 3984 35402 4020
rect 38290 9424 38346 9480
rect 38842 13368 38898 13424
rect 37066 9274 37122 9276
rect 37146 9274 37202 9276
rect 37226 9274 37282 9276
rect 37306 9274 37362 9276
rect 37066 9222 37112 9274
rect 37112 9222 37122 9274
rect 37146 9222 37176 9274
rect 37176 9222 37188 9274
rect 37188 9222 37202 9274
rect 37226 9222 37240 9274
rect 37240 9222 37252 9274
rect 37252 9222 37282 9274
rect 37306 9222 37316 9274
rect 37316 9222 37362 9274
rect 37066 9220 37122 9222
rect 37146 9220 37202 9222
rect 37226 9220 37282 9222
rect 37306 9220 37362 9222
rect 37066 8186 37122 8188
rect 37146 8186 37202 8188
rect 37226 8186 37282 8188
rect 37306 8186 37362 8188
rect 37066 8134 37112 8186
rect 37112 8134 37122 8186
rect 37146 8134 37176 8186
rect 37176 8134 37188 8186
rect 37188 8134 37202 8186
rect 37226 8134 37240 8186
rect 37240 8134 37252 8186
rect 37252 8134 37282 8186
rect 37306 8134 37316 8186
rect 37316 8134 37362 8186
rect 37066 8132 37122 8134
rect 37146 8132 37202 8134
rect 37226 8132 37282 8134
rect 37306 8132 37362 8134
rect 37066 7098 37122 7100
rect 37146 7098 37202 7100
rect 37226 7098 37282 7100
rect 37306 7098 37362 7100
rect 37066 7046 37112 7098
rect 37112 7046 37122 7098
rect 37146 7046 37176 7098
rect 37176 7046 37188 7098
rect 37188 7046 37202 7098
rect 37226 7046 37240 7098
rect 37240 7046 37252 7098
rect 37252 7046 37282 7098
rect 37306 7046 37316 7098
rect 37316 7046 37362 7098
rect 37066 7044 37122 7046
rect 37146 7044 37202 7046
rect 37226 7044 37282 7046
rect 37306 7044 37362 7046
rect 37066 6010 37122 6012
rect 37146 6010 37202 6012
rect 37226 6010 37282 6012
rect 37306 6010 37362 6012
rect 37066 5958 37112 6010
rect 37112 5958 37122 6010
rect 37146 5958 37176 6010
rect 37176 5958 37188 6010
rect 37188 5958 37202 6010
rect 37226 5958 37240 6010
rect 37240 5958 37252 6010
rect 37252 5958 37282 6010
rect 37306 5958 37316 6010
rect 37316 5958 37362 6010
rect 37066 5956 37122 5958
rect 37146 5956 37202 5958
rect 37226 5956 37282 5958
rect 37306 5956 37362 5958
rect 37066 4922 37122 4924
rect 37146 4922 37202 4924
rect 37226 4922 37282 4924
rect 37306 4922 37362 4924
rect 37066 4870 37112 4922
rect 37112 4870 37122 4922
rect 37146 4870 37176 4922
rect 37176 4870 37188 4922
rect 37188 4870 37202 4922
rect 37226 4870 37240 4922
rect 37240 4870 37252 4922
rect 37252 4870 37282 4922
rect 37306 4870 37316 4922
rect 37316 4870 37362 4922
rect 37066 4868 37122 4870
rect 37146 4868 37202 4870
rect 37226 4868 37282 4870
rect 37306 4868 37362 4870
rect 38474 7404 38530 7440
rect 38474 7384 38476 7404
rect 38476 7384 38528 7404
rect 38528 7384 38530 7404
rect 36818 3848 36874 3904
rect 37066 3834 37122 3836
rect 37146 3834 37202 3836
rect 37226 3834 37282 3836
rect 37306 3834 37362 3836
rect 37066 3782 37112 3834
rect 37112 3782 37122 3834
rect 37146 3782 37176 3834
rect 37176 3782 37188 3834
rect 37188 3782 37202 3834
rect 37226 3782 37240 3834
rect 37240 3782 37252 3834
rect 37252 3782 37282 3834
rect 37306 3782 37316 3834
rect 37316 3782 37362 3834
rect 37066 3780 37122 3782
rect 37146 3780 37202 3782
rect 37226 3780 37282 3782
rect 37306 3780 37362 3782
rect 37066 2746 37122 2748
rect 37146 2746 37202 2748
rect 37226 2746 37282 2748
rect 37306 2746 37362 2748
rect 37066 2694 37112 2746
rect 37112 2694 37122 2746
rect 37146 2694 37176 2746
rect 37176 2694 37188 2746
rect 37188 2694 37202 2746
rect 37226 2694 37240 2746
rect 37240 2694 37252 2746
rect 37252 2694 37282 2746
rect 37306 2694 37316 2746
rect 37316 2694 37362 2746
rect 37066 2692 37122 2694
rect 37146 2692 37202 2694
rect 37226 2692 37282 2694
rect 37306 2692 37362 2694
rect 41050 12960 41106 13016
rect 40038 12688 40094 12744
rect 43718 19760 43774 19816
rect 44288 20698 44344 20700
rect 44368 20698 44424 20700
rect 44448 20698 44504 20700
rect 44528 20698 44584 20700
rect 44288 20646 44334 20698
rect 44334 20646 44344 20698
rect 44368 20646 44398 20698
rect 44398 20646 44410 20698
rect 44410 20646 44424 20698
rect 44448 20646 44462 20698
rect 44462 20646 44474 20698
rect 44474 20646 44504 20698
rect 44528 20646 44538 20698
rect 44538 20646 44584 20698
rect 44288 20644 44344 20646
rect 44368 20644 44424 20646
rect 44448 20644 44504 20646
rect 44528 20644 44584 20646
rect 44288 19610 44344 19612
rect 44368 19610 44424 19612
rect 44448 19610 44504 19612
rect 44528 19610 44584 19612
rect 44288 19558 44334 19610
rect 44334 19558 44344 19610
rect 44368 19558 44398 19610
rect 44398 19558 44410 19610
rect 44410 19558 44424 19610
rect 44448 19558 44462 19610
rect 44462 19558 44474 19610
rect 44474 19558 44504 19610
rect 44528 19558 44538 19610
rect 44538 19558 44584 19610
rect 44288 19556 44344 19558
rect 44368 19556 44424 19558
rect 44448 19556 44504 19558
rect 44528 19556 44584 19558
rect 40130 7112 40186 7168
rect 39854 6976 39910 7032
rect 39946 3984 40002 4040
rect 40682 7420 40684 7440
rect 40684 7420 40736 7440
rect 40736 7420 40738 7440
rect 40682 7384 40738 7420
rect 44288 18522 44344 18524
rect 44368 18522 44424 18524
rect 44448 18522 44504 18524
rect 44528 18522 44584 18524
rect 44288 18470 44334 18522
rect 44334 18470 44344 18522
rect 44368 18470 44398 18522
rect 44398 18470 44410 18522
rect 44410 18470 44424 18522
rect 44448 18470 44462 18522
rect 44462 18470 44474 18522
rect 44474 18470 44504 18522
rect 44528 18470 44538 18522
rect 44538 18470 44584 18522
rect 44288 18468 44344 18470
rect 44368 18468 44424 18470
rect 44448 18468 44504 18470
rect 44528 18468 44584 18470
rect 44288 17434 44344 17436
rect 44368 17434 44424 17436
rect 44448 17434 44504 17436
rect 44528 17434 44584 17436
rect 44288 17382 44334 17434
rect 44334 17382 44344 17434
rect 44368 17382 44398 17434
rect 44398 17382 44410 17434
rect 44410 17382 44424 17434
rect 44448 17382 44462 17434
rect 44462 17382 44474 17434
rect 44474 17382 44504 17434
rect 44528 17382 44538 17434
rect 44538 17382 44584 17434
rect 44288 17380 44344 17382
rect 44368 17380 44424 17382
rect 44448 17380 44504 17382
rect 44528 17380 44584 17382
rect 44288 16346 44344 16348
rect 44368 16346 44424 16348
rect 44448 16346 44504 16348
rect 44528 16346 44584 16348
rect 44288 16294 44334 16346
rect 44334 16294 44344 16346
rect 44368 16294 44398 16346
rect 44398 16294 44410 16346
rect 44410 16294 44424 16346
rect 44448 16294 44462 16346
rect 44462 16294 44474 16346
rect 44474 16294 44504 16346
rect 44528 16294 44538 16346
rect 44538 16294 44584 16346
rect 44288 16292 44344 16294
rect 44368 16292 44424 16294
rect 44448 16292 44504 16294
rect 44528 16292 44584 16294
rect 44288 15258 44344 15260
rect 44368 15258 44424 15260
rect 44448 15258 44504 15260
rect 44528 15258 44584 15260
rect 44288 15206 44334 15258
rect 44334 15206 44344 15258
rect 44368 15206 44398 15258
rect 44398 15206 44410 15258
rect 44410 15206 44424 15258
rect 44448 15206 44462 15258
rect 44462 15206 44474 15258
rect 44474 15206 44504 15258
rect 44528 15206 44538 15258
rect 44538 15206 44584 15258
rect 44288 15204 44344 15206
rect 44368 15204 44424 15206
rect 44448 15204 44504 15206
rect 44528 15204 44584 15206
rect 44288 14170 44344 14172
rect 44368 14170 44424 14172
rect 44448 14170 44504 14172
rect 44528 14170 44584 14172
rect 44288 14118 44334 14170
rect 44334 14118 44344 14170
rect 44368 14118 44398 14170
rect 44398 14118 44410 14170
rect 44410 14118 44424 14170
rect 44448 14118 44462 14170
rect 44462 14118 44474 14170
rect 44474 14118 44504 14170
rect 44528 14118 44538 14170
rect 44538 14118 44584 14170
rect 44288 14116 44344 14118
rect 44368 14116 44424 14118
rect 44448 14116 44504 14118
rect 44528 14116 44584 14118
rect 44288 13082 44344 13084
rect 44368 13082 44424 13084
rect 44448 13082 44504 13084
rect 44528 13082 44584 13084
rect 44288 13030 44334 13082
rect 44334 13030 44344 13082
rect 44368 13030 44398 13082
rect 44398 13030 44410 13082
rect 44410 13030 44424 13082
rect 44448 13030 44462 13082
rect 44462 13030 44474 13082
rect 44474 13030 44504 13082
rect 44528 13030 44538 13082
rect 44538 13030 44584 13082
rect 44288 13028 44344 13030
rect 44368 13028 44424 13030
rect 44448 13028 44504 13030
rect 44528 13028 44584 13030
rect 44288 11994 44344 11996
rect 44368 11994 44424 11996
rect 44448 11994 44504 11996
rect 44528 11994 44584 11996
rect 44288 11942 44334 11994
rect 44334 11942 44344 11994
rect 44368 11942 44398 11994
rect 44398 11942 44410 11994
rect 44410 11942 44424 11994
rect 44448 11942 44462 11994
rect 44462 11942 44474 11994
rect 44474 11942 44504 11994
rect 44528 11942 44538 11994
rect 44538 11942 44584 11994
rect 44288 11940 44344 11942
rect 44368 11940 44424 11942
rect 44448 11940 44504 11942
rect 44528 11940 44584 11942
rect 41050 4020 41052 4040
rect 41052 4020 41104 4040
rect 41104 4020 41106 4040
rect 41050 3984 41106 4020
rect 44288 10906 44344 10908
rect 44368 10906 44424 10908
rect 44448 10906 44504 10908
rect 44528 10906 44584 10908
rect 44288 10854 44334 10906
rect 44334 10854 44344 10906
rect 44368 10854 44398 10906
rect 44398 10854 44410 10906
rect 44410 10854 44424 10906
rect 44448 10854 44462 10906
rect 44462 10854 44474 10906
rect 44474 10854 44504 10906
rect 44528 10854 44538 10906
rect 44538 10854 44584 10906
rect 44288 10852 44344 10854
rect 44368 10852 44424 10854
rect 44448 10852 44504 10854
rect 44528 10852 44584 10854
rect 44288 9818 44344 9820
rect 44368 9818 44424 9820
rect 44448 9818 44504 9820
rect 44528 9818 44584 9820
rect 44288 9766 44334 9818
rect 44334 9766 44344 9818
rect 44368 9766 44398 9818
rect 44398 9766 44410 9818
rect 44410 9766 44424 9818
rect 44448 9766 44462 9818
rect 44462 9766 44474 9818
rect 44474 9766 44504 9818
rect 44528 9766 44538 9818
rect 44538 9766 44584 9818
rect 44288 9764 44344 9766
rect 44368 9764 44424 9766
rect 44448 9764 44504 9766
rect 44528 9764 44584 9766
rect 44288 8730 44344 8732
rect 44368 8730 44424 8732
rect 44448 8730 44504 8732
rect 44528 8730 44584 8732
rect 44288 8678 44334 8730
rect 44334 8678 44344 8730
rect 44368 8678 44398 8730
rect 44398 8678 44410 8730
rect 44410 8678 44424 8730
rect 44448 8678 44462 8730
rect 44462 8678 44474 8730
rect 44474 8678 44504 8730
rect 44528 8678 44538 8730
rect 44538 8678 44584 8730
rect 44288 8676 44344 8678
rect 44368 8676 44424 8678
rect 44448 8676 44504 8678
rect 44528 8676 44584 8678
rect 44288 7642 44344 7644
rect 44368 7642 44424 7644
rect 44448 7642 44504 7644
rect 44528 7642 44584 7644
rect 44288 7590 44334 7642
rect 44334 7590 44344 7642
rect 44368 7590 44398 7642
rect 44398 7590 44410 7642
rect 44410 7590 44424 7642
rect 44448 7590 44462 7642
rect 44462 7590 44474 7642
rect 44474 7590 44504 7642
rect 44528 7590 44538 7642
rect 44538 7590 44584 7642
rect 44288 7588 44344 7590
rect 44368 7588 44424 7590
rect 44448 7588 44504 7590
rect 44528 7588 44584 7590
rect 44086 7420 44088 7440
rect 44088 7420 44140 7440
rect 44140 7420 44142 7440
rect 44086 7384 44142 7420
rect 44288 6554 44344 6556
rect 44368 6554 44424 6556
rect 44448 6554 44504 6556
rect 44528 6554 44584 6556
rect 44288 6502 44334 6554
rect 44334 6502 44344 6554
rect 44368 6502 44398 6554
rect 44398 6502 44410 6554
rect 44410 6502 44424 6554
rect 44448 6502 44462 6554
rect 44462 6502 44474 6554
rect 44474 6502 44504 6554
rect 44528 6502 44538 6554
rect 44538 6502 44584 6554
rect 44288 6500 44344 6502
rect 44368 6500 44424 6502
rect 44448 6500 44504 6502
rect 44528 6500 44584 6502
rect 42890 4528 42946 4584
rect 42890 2896 42946 2952
rect 44178 5636 44234 5672
rect 44178 5616 44180 5636
rect 44180 5616 44232 5636
rect 44232 5616 44234 5636
rect 44288 5466 44344 5468
rect 44368 5466 44424 5468
rect 44448 5466 44504 5468
rect 44528 5466 44584 5468
rect 44288 5414 44334 5466
rect 44334 5414 44344 5466
rect 44368 5414 44398 5466
rect 44398 5414 44410 5466
rect 44410 5414 44424 5466
rect 44448 5414 44462 5466
rect 44462 5414 44474 5466
rect 44474 5414 44504 5466
rect 44528 5414 44538 5466
rect 44538 5414 44584 5466
rect 44288 5412 44344 5414
rect 44368 5412 44424 5414
rect 44448 5412 44504 5414
rect 44528 5412 44584 5414
rect 44288 4378 44344 4380
rect 44368 4378 44424 4380
rect 44448 4378 44504 4380
rect 44528 4378 44584 4380
rect 44288 4326 44334 4378
rect 44334 4326 44344 4378
rect 44368 4326 44398 4378
rect 44398 4326 44410 4378
rect 44410 4326 44424 4378
rect 44448 4326 44462 4378
rect 44462 4326 44474 4378
rect 44474 4326 44504 4378
rect 44528 4326 44538 4378
rect 44538 4326 44584 4378
rect 44288 4324 44344 4326
rect 44368 4324 44424 4326
rect 44448 4324 44504 4326
rect 44528 4324 44584 4326
rect 44288 3290 44344 3292
rect 44368 3290 44424 3292
rect 44448 3290 44504 3292
rect 44528 3290 44584 3292
rect 44288 3238 44334 3290
rect 44334 3238 44344 3290
rect 44368 3238 44398 3290
rect 44398 3238 44410 3290
rect 44410 3238 44424 3290
rect 44448 3238 44462 3290
rect 44462 3238 44474 3290
rect 44474 3238 44504 3290
rect 44528 3238 44538 3290
rect 44538 3238 44584 3290
rect 44288 3236 44344 3238
rect 44368 3236 44424 3238
rect 44448 3236 44504 3238
rect 44528 3236 44584 3238
rect 44822 7148 44824 7168
rect 44824 7148 44876 7168
rect 44876 7148 44878 7168
rect 44822 7112 44878 7148
rect 44914 6976 44970 7032
rect 44288 2202 44344 2204
rect 44368 2202 44424 2204
rect 44448 2202 44504 2204
rect 44528 2202 44584 2204
rect 44288 2150 44334 2202
rect 44334 2150 44344 2202
rect 44368 2150 44398 2202
rect 44398 2150 44410 2202
rect 44410 2150 44424 2202
rect 44448 2150 44462 2202
rect 44462 2150 44474 2202
rect 44474 2150 44504 2202
rect 44528 2150 44538 2202
rect 44538 2150 44584 2202
rect 44288 2148 44344 2150
rect 44368 2148 44424 2150
rect 44448 2148 44504 2150
rect 44528 2148 44584 2150
rect 51510 21242 51566 21244
rect 51590 21242 51646 21244
rect 51670 21242 51726 21244
rect 51750 21242 51806 21244
rect 51510 21190 51556 21242
rect 51556 21190 51566 21242
rect 51590 21190 51620 21242
rect 51620 21190 51632 21242
rect 51632 21190 51646 21242
rect 51670 21190 51684 21242
rect 51684 21190 51696 21242
rect 51696 21190 51726 21242
rect 51750 21190 51760 21242
rect 51760 21190 51806 21242
rect 51510 21188 51566 21190
rect 51590 21188 51646 21190
rect 51670 21188 51726 21190
rect 51750 21188 51806 21190
rect 51510 20154 51566 20156
rect 51590 20154 51646 20156
rect 51670 20154 51726 20156
rect 51750 20154 51806 20156
rect 51510 20102 51556 20154
rect 51556 20102 51566 20154
rect 51590 20102 51620 20154
rect 51620 20102 51632 20154
rect 51632 20102 51646 20154
rect 51670 20102 51684 20154
rect 51684 20102 51696 20154
rect 51696 20102 51726 20154
rect 51750 20102 51760 20154
rect 51760 20102 51806 20154
rect 51510 20100 51566 20102
rect 51590 20100 51646 20102
rect 51670 20100 51726 20102
rect 51750 20100 51806 20102
rect 52826 20440 52882 20496
rect 45098 3984 45154 4040
rect 46938 3576 46994 3632
rect 48778 6840 48834 6896
rect 51510 19066 51566 19068
rect 51590 19066 51646 19068
rect 51670 19066 51726 19068
rect 51750 19066 51806 19068
rect 51510 19014 51556 19066
rect 51556 19014 51566 19066
rect 51590 19014 51620 19066
rect 51620 19014 51632 19066
rect 51632 19014 51646 19066
rect 51670 19014 51684 19066
rect 51684 19014 51696 19066
rect 51696 19014 51726 19066
rect 51750 19014 51760 19066
rect 51760 19014 51806 19066
rect 51510 19012 51566 19014
rect 51590 19012 51646 19014
rect 51670 19012 51726 19014
rect 51750 19012 51806 19014
rect 51510 17978 51566 17980
rect 51590 17978 51646 17980
rect 51670 17978 51726 17980
rect 51750 17978 51806 17980
rect 51510 17926 51556 17978
rect 51556 17926 51566 17978
rect 51590 17926 51620 17978
rect 51620 17926 51632 17978
rect 51632 17926 51646 17978
rect 51670 17926 51684 17978
rect 51684 17926 51696 17978
rect 51696 17926 51726 17978
rect 51750 17926 51760 17978
rect 51760 17926 51806 17978
rect 51510 17924 51566 17926
rect 51590 17924 51646 17926
rect 51670 17924 51726 17926
rect 51750 17924 51806 17926
rect 51510 16890 51566 16892
rect 51590 16890 51646 16892
rect 51670 16890 51726 16892
rect 51750 16890 51806 16892
rect 51510 16838 51556 16890
rect 51556 16838 51566 16890
rect 51590 16838 51620 16890
rect 51620 16838 51632 16890
rect 51632 16838 51646 16890
rect 51670 16838 51684 16890
rect 51684 16838 51696 16890
rect 51696 16838 51726 16890
rect 51750 16838 51760 16890
rect 51760 16838 51806 16890
rect 51510 16836 51566 16838
rect 51590 16836 51646 16838
rect 51670 16836 51726 16838
rect 51750 16836 51806 16838
rect 51510 15802 51566 15804
rect 51590 15802 51646 15804
rect 51670 15802 51726 15804
rect 51750 15802 51806 15804
rect 51510 15750 51556 15802
rect 51556 15750 51566 15802
rect 51590 15750 51620 15802
rect 51620 15750 51632 15802
rect 51632 15750 51646 15802
rect 51670 15750 51684 15802
rect 51684 15750 51696 15802
rect 51696 15750 51726 15802
rect 51750 15750 51760 15802
rect 51760 15750 51806 15802
rect 51510 15748 51566 15750
rect 51590 15748 51646 15750
rect 51670 15748 51726 15750
rect 51750 15748 51806 15750
rect 51510 14714 51566 14716
rect 51590 14714 51646 14716
rect 51670 14714 51726 14716
rect 51750 14714 51806 14716
rect 51510 14662 51556 14714
rect 51556 14662 51566 14714
rect 51590 14662 51620 14714
rect 51620 14662 51632 14714
rect 51632 14662 51646 14714
rect 51670 14662 51684 14714
rect 51684 14662 51696 14714
rect 51696 14662 51726 14714
rect 51750 14662 51760 14714
rect 51760 14662 51806 14714
rect 51510 14660 51566 14662
rect 51590 14660 51646 14662
rect 51670 14660 51726 14662
rect 51750 14660 51806 14662
rect 51510 13626 51566 13628
rect 51590 13626 51646 13628
rect 51670 13626 51726 13628
rect 51750 13626 51806 13628
rect 51510 13574 51556 13626
rect 51556 13574 51566 13626
rect 51590 13574 51620 13626
rect 51620 13574 51632 13626
rect 51632 13574 51646 13626
rect 51670 13574 51684 13626
rect 51684 13574 51696 13626
rect 51696 13574 51726 13626
rect 51750 13574 51760 13626
rect 51760 13574 51806 13626
rect 51510 13572 51566 13574
rect 51590 13572 51646 13574
rect 51670 13572 51726 13574
rect 51750 13572 51806 13574
rect 51510 12538 51566 12540
rect 51590 12538 51646 12540
rect 51670 12538 51726 12540
rect 51750 12538 51806 12540
rect 51510 12486 51556 12538
rect 51556 12486 51566 12538
rect 51590 12486 51620 12538
rect 51620 12486 51632 12538
rect 51632 12486 51646 12538
rect 51670 12486 51684 12538
rect 51684 12486 51696 12538
rect 51696 12486 51726 12538
rect 51750 12486 51760 12538
rect 51760 12486 51806 12538
rect 51510 12484 51566 12486
rect 51590 12484 51646 12486
rect 51670 12484 51726 12486
rect 51750 12484 51806 12486
rect 51510 11450 51566 11452
rect 51590 11450 51646 11452
rect 51670 11450 51726 11452
rect 51750 11450 51806 11452
rect 51510 11398 51556 11450
rect 51556 11398 51566 11450
rect 51590 11398 51620 11450
rect 51620 11398 51632 11450
rect 51632 11398 51646 11450
rect 51670 11398 51684 11450
rect 51684 11398 51696 11450
rect 51696 11398 51726 11450
rect 51750 11398 51760 11450
rect 51760 11398 51806 11450
rect 51510 11396 51566 11398
rect 51590 11396 51646 11398
rect 51670 11396 51726 11398
rect 51750 11396 51806 11398
rect 51510 10362 51566 10364
rect 51590 10362 51646 10364
rect 51670 10362 51726 10364
rect 51750 10362 51806 10364
rect 51510 10310 51556 10362
rect 51556 10310 51566 10362
rect 51590 10310 51620 10362
rect 51620 10310 51632 10362
rect 51632 10310 51646 10362
rect 51670 10310 51684 10362
rect 51684 10310 51696 10362
rect 51696 10310 51726 10362
rect 51750 10310 51760 10362
rect 51760 10310 51806 10362
rect 51510 10308 51566 10310
rect 51590 10308 51646 10310
rect 51670 10308 51726 10310
rect 51750 10308 51806 10310
rect 51510 9274 51566 9276
rect 51590 9274 51646 9276
rect 51670 9274 51726 9276
rect 51750 9274 51806 9276
rect 51510 9222 51556 9274
rect 51556 9222 51566 9274
rect 51590 9222 51620 9274
rect 51620 9222 51632 9274
rect 51632 9222 51646 9274
rect 51670 9222 51684 9274
rect 51684 9222 51696 9274
rect 51696 9222 51726 9274
rect 51750 9222 51760 9274
rect 51760 9222 51806 9274
rect 51510 9220 51566 9222
rect 51590 9220 51646 9222
rect 51670 9220 51726 9222
rect 51750 9220 51806 9222
rect 52274 13268 52276 13288
rect 52276 13268 52328 13288
rect 52328 13268 52330 13288
rect 52274 13232 52330 13268
rect 52090 8472 52146 8528
rect 51510 8186 51566 8188
rect 51590 8186 51646 8188
rect 51670 8186 51726 8188
rect 51750 8186 51806 8188
rect 51510 8134 51556 8186
rect 51556 8134 51566 8186
rect 51590 8134 51620 8186
rect 51620 8134 51632 8186
rect 51632 8134 51646 8186
rect 51670 8134 51684 8186
rect 51684 8134 51696 8186
rect 51696 8134 51726 8186
rect 51750 8134 51760 8186
rect 51760 8134 51806 8186
rect 51510 8132 51566 8134
rect 51590 8132 51646 8134
rect 51670 8132 51726 8134
rect 51750 8132 51806 8134
rect 51510 7098 51566 7100
rect 51590 7098 51646 7100
rect 51670 7098 51726 7100
rect 51750 7098 51806 7100
rect 51510 7046 51556 7098
rect 51556 7046 51566 7098
rect 51590 7046 51620 7098
rect 51620 7046 51632 7098
rect 51632 7046 51646 7098
rect 51670 7046 51684 7098
rect 51684 7046 51696 7098
rect 51696 7046 51726 7098
rect 51750 7046 51760 7098
rect 51760 7046 51806 7098
rect 51510 7044 51566 7046
rect 51590 7044 51646 7046
rect 51670 7044 51726 7046
rect 51750 7044 51806 7046
rect 51510 6010 51566 6012
rect 51590 6010 51646 6012
rect 51670 6010 51726 6012
rect 51750 6010 51806 6012
rect 51510 5958 51556 6010
rect 51556 5958 51566 6010
rect 51590 5958 51620 6010
rect 51620 5958 51632 6010
rect 51632 5958 51646 6010
rect 51670 5958 51684 6010
rect 51684 5958 51696 6010
rect 51696 5958 51726 6010
rect 51750 5958 51760 6010
rect 51760 5958 51806 6010
rect 51510 5956 51566 5958
rect 51590 5956 51646 5958
rect 51670 5956 51726 5958
rect 51750 5956 51806 5958
rect 51510 4922 51566 4924
rect 51590 4922 51646 4924
rect 51670 4922 51726 4924
rect 51750 4922 51806 4924
rect 51510 4870 51556 4922
rect 51556 4870 51566 4922
rect 51590 4870 51620 4922
rect 51620 4870 51632 4922
rect 51632 4870 51646 4922
rect 51670 4870 51684 4922
rect 51684 4870 51696 4922
rect 51696 4870 51726 4922
rect 51750 4870 51760 4922
rect 51760 4870 51806 4922
rect 51510 4868 51566 4870
rect 51590 4868 51646 4870
rect 51670 4868 51726 4870
rect 51750 4868 51806 4870
rect 51510 3834 51566 3836
rect 51590 3834 51646 3836
rect 51670 3834 51726 3836
rect 51750 3834 51806 3836
rect 51510 3782 51556 3834
rect 51556 3782 51566 3834
rect 51590 3782 51620 3834
rect 51620 3782 51632 3834
rect 51632 3782 51646 3834
rect 51670 3782 51684 3834
rect 51684 3782 51696 3834
rect 51696 3782 51726 3834
rect 51750 3782 51760 3834
rect 51760 3782 51806 3834
rect 51510 3780 51566 3782
rect 51590 3780 51646 3782
rect 51670 3780 51726 3782
rect 51750 3780 51806 3782
rect 51510 2746 51566 2748
rect 51590 2746 51646 2748
rect 51670 2746 51726 2748
rect 51750 2746 51806 2748
rect 51510 2694 51556 2746
rect 51556 2694 51566 2746
rect 51590 2694 51620 2746
rect 51620 2694 51632 2746
rect 51632 2694 51646 2746
rect 51670 2694 51684 2746
rect 51684 2694 51696 2746
rect 51696 2694 51726 2746
rect 51750 2694 51760 2746
rect 51760 2694 51806 2746
rect 51510 2692 51566 2694
rect 51590 2692 51646 2694
rect 51670 2692 51726 2694
rect 51750 2692 51806 2694
rect 52826 10512 52882 10568
rect 53746 8780 53748 8800
rect 53748 8780 53800 8800
rect 53800 8780 53802 8800
rect 53746 8744 53802 8780
rect 52734 5636 52790 5672
rect 52734 5616 52736 5636
rect 52736 5616 52788 5636
rect 52788 5616 52790 5636
rect 58732 20698 58788 20700
rect 58812 20698 58868 20700
rect 58892 20698 58948 20700
rect 58972 20698 59028 20700
rect 58732 20646 58778 20698
rect 58778 20646 58788 20698
rect 58812 20646 58842 20698
rect 58842 20646 58854 20698
rect 58854 20646 58868 20698
rect 58892 20646 58906 20698
rect 58906 20646 58918 20698
rect 58918 20646 58948 20698
rect 58972 20646 58982 20698
rect 58982 20646 59028 20698
rect 58732 20644 58788 20646
rect 58812 20644 58868 20646
rect 58892 20644 58948 20646
rect 58972 20644 59028 20646
rect 58732 19610 58788 19612
rect 58812 19610 58868 19612
rect 58892 19610 58948 19612
rect 58972 19610 59028 19612
rect 58732 19558 58778 19610
rect 58778 19558 58788 19610
rect 58812 19558 58842 19610
rect 58842 19558 58854 19610
rect 58854 19558 58868 19610
rect 58892 19558 58906 19610
rect 58906 19558 58918 19610
rect 58918 19558 58948 19610
rect 58972 19558 58982 19610
rect 58982 19558 59028 19610
rect 58732 19556 58788 19558
rect 58812 19556 58868 19558
rect 58892 19556 58948 19558
rect 58972 19556 59028 19558
rect 54206 7248 54262 7304
rect 56690 13232 56746 13288
rect 56046 9016 56102 9072
rect 55862 6976 55918 7032
rect 55494 6860 55550 6896
rect 55494 6840 55496 6860
rect 55496 6840 55548 6860
rect 55548 6840 55550 6860
rect 56874 8880 56930 8936
rect 56874 8780 56876 8800
rect 56876 8780 56928 8800
rect 56928 8780 56930 8800
rect 56874 8744 56930 8780
rect 56690 4020 56692 4040
rect 56692 4020 56744 4040
rect 56744 4020 56746 4040
rect 56690 3984 56746 4020
rect 58732 18522 58788 18524
rect 58812 18522 58868 18524
rect 58892 18522 58948 18524
rect 58972 18522 59028 18524
rect 58732 18470 58778 18522
rect 58778 18470 58788 18522
rect 58812 18470 58842 18522
rect 58842 18470 58854 18522
rect 58854 18470 58868 18522
rect 58892 18470 58906 18522
rect 58906 18470 58918 18522
rect 58918 18470 58948 18522
rect 58972 18470 58982 18522
rect 58982 18470 59028 18522
rect 58732 18468 58788 18470
rect 58812 18468 58868 18470
rect 58892 18468 58948 18470
rect 58972 18468 59028 18470
rect 58732 17434 58788 17436
rect 58812 17434 58868 17436
rect 58892 17434 58948 17436
rect 58972 17434 59028 17436
rect 58732 17382 58778 17434
rect 58778 17382 58788 17434
rect 58812 17382 58842 17434
rect 58842 17382 58854 17434
rect 58854 17382 58868 17434
rect 58892 17382 58906 17434
rect 58906 17382 58918 17434
rect 58918 17382 58948 17434
rect 58972 17382 58982 17434
rect 58982 17382 59028 17434
rect 58732 17380 58788 17382
rect 58812 17380 58868 17382
rect 58892 17380 58948 17382
rect 58972 17380 59028 17382
rect 58732 16346 58788 16348
rect 58812 16346 58868 16348
rect 58892 16346 58948 16348
rect 58972 16346 59028 16348
rect 58732 16294 58778 16346
rect 58778 16294 58788 16346
rect 58812 16294 58842 16346
rect 58842 16294 58854 16346
rect 58854 16294 58868 16346
rect 58892 16294 58906 16346
rect 58906 16294 58918 16346
rect 58918 16294 58948 16346
rect 58972 16294 58982 16346
rect 58982 16294 59028 16346
rect 58732 16292 58788 16294
rect 58812 16292 58868 16294
rect 58892 16292 58948 16294
rect 58972 16292 59028 16294
rect 58732 15258 58788 15260
rect 58812 15258 58868 15260
rect 58892 15258 58948 15260
rect 58972 15258 59028 15260
rect 58732 15206 58778 15258
rect 58778 15206 58788 15258
rect 58812 15206 58842 15258
rect 58842 15206 58854 15258
rect 58854 15206 58868 15258
rect 58892 15206 58906 15258
rect 58906 15206 58918 15258
rect 58918 15206 58948 15258
rect 58972 15206 58982 15258
rect 58982 15206 59028 15258
rect 58732 15204 58788 15206
rect 58812 15204 58868 15206
rect 58892 15204 58948 15206
rect 58972 15204 59028 15206
rect 58732 14170 58788 14172
rect 58812 14170 58868 14172
rect 58892 14170 58948 14172
rect 58972 14170 59028 14172
rect 58732 14118 58778 14170
rect 58778 14118 58788 14170
rect 58812 14118 58842 14170
rect 58842 14118 58854 14170
rect 58854 14118 58868 14170
rect 58892 14118 58906 14170
rect 58906 14118 58918 14170
rect 58918 14118 58948 14170
rect 58972 14118 58982 14170
rect 58982 14118 59028 14170
rect 58732 14116 58788 14118
rect 58812 14116 58868 14118
rect 58892 14116 58948 14118
rect 58972 14116 59028 14118
rect 58732 13082 58788 13084
rect 58812 13082 58868 13084
rect 58892 13082 58948 13084
rect 58972 13082 59028 13084
rect 58732 13030 58778 13082
rect 58778 13030 58788 13082
rect 58812 13030 58842 13082
rect 58842 13030 58854 13082
rect 58854 13030 58868 13082
rect 58892 13030 58906 13082
rect 58906 13030 58918 13082
rect 58918 13030 58948 13082
rect 58972 13030 58982 13082
rect 58982 13030 59028 13082
rect 58732 13028 58788 13030
rect 58812 13028 58868 13030
rect 58892 13028 58948 13030
rect 58972 13028 59028 13030
rect 58732 11994 58788 11996
rect 58812 11994 58868 11996
rect 58892 11994 58948 11996
rect 58972 11994 59028 11996
rect 58732 11942 58778 11994
rect 58778 11942 58788 11994
rect 58812 11942 58842 11994
rect 58842 11942 58854 11994
rect 58854 11942 58868 11994
rect 58892 11942 58906 11994
rect 58906 11942 58918 11994
rect 58918 11942 58948 11994
rect 58972 11942 58982 11994
rect 58982 11942 59028 11994
rect 58732 11940 58788 11942
rect 58812 11940 58868 11942
rect 58892 11940 58948 11942
rect 58972 11940 59028 11942
rect 58732 10906 58788 10908
rect 58812 10906 58868 10908
rect 58892 10906 58948 10908
rect 58972 10906 59028 10908
rect 58732 10854 58778 10906
rect 58778 10854 58788 10906
rect 58812 10854 58842 10906
rect 58842 10854 58854 10906
rect 58854 10854 58868 10906
rect 58892 10854 58906 10906
rect 58906 10854 58918 10906
rect 58918 10854 58948 10906
rect 58972 10854 58982 10906
rect 58982 10854 59028 10906
rect 58732 10852 58788 10854
rect 58812 10852 58868 10854
rect 58892 10852 58948 10854
rect 58972 10852 59028 10854
rect 58732 9818 58788 9820
rect 58812 9818 58868 9820
rect 58892 9818 58948 9820
rect 58972 9818 59028 9820
rect 58732 9766 58778 9818
rect 58778 9766 58788 9818
rect 58812 9766 58842 9818
rect 58842 9766 58854 9818
rect 58854 9766 58868 9818
rect 58892 9766 58906 9818
rect 58906 9766 58918 9818
rect 58918 9766 58948 9818
rect 58972 9766 58982 9818
rect 58982 9766 59028 9818
rect 58732 9764 58788 9766
rect 58812 9764 58868 9766
rect 58892 9764 58948 9766
rect 58972 9764 59028 9766
rect 58732 8730 58788 8732
rect 58812 8730 58868 8732
rect 58892 8730 58948 8732
rect 58972 8730 59028 8732
rect 58732 8678 58778 8730
rect 58778 8678 58788 8730
rect 58812 8678 58842 8730
rect 58842 8678 58854 8730
rect 58854 8678 58868 8730
rect 58892 8678 58906 8730
rect 58906 8678 58918 8730
rect 58918 8678 58948 8730
rect 58972 8678 58982 8730
rect 58982 8678 59028 8730
rect 58732 8676 58788 8678
rect 58812 8676 58868 8678
rect 58892 8676 58948 8678
rect 58972 8676 59028 8678
rect 58732 7642 58788 7644
rect 58812 7642 58868 7644
rect 58892 7642 58948 7644
rect 58972 7642 59028 7644
rect 58732 7590 58778 7642
rect 58778 7590 58788 7642
rect 58812 7590 58842 7642
rect 58842 7590 58854 7642
rect 58854 7590 58868 7642
rect 58892 7590 58906 7642
rect 58906 7590 58918 7642
rect 58918 7590 58948 7642
rect 58972 7590 58982 7642
rect 58982 7590 59028 7642
rect 58732 7588 58788 7590
rect 58812 7588 58868 7590
rect 58892 7588 58948 7590
rect 58972 7588 59028 7590
rect 58732 6554 58788 6556
rect 58812 6554 58868 6556
rect 58892 6554 58948 6556
rect 58972 6554 59028 6556
rect 58732 6502 58778 6554
rect 58778 6502 58788 6554
rect 58812 6502 58842 6554
rect 58842 6502 58854 6554
rect 58854 6502 58868 6554
rect 58892 6502 58906 6554
rect 58906 6502 58918 6554
rect 58918 6502 58948 6554
rect 58972 6502 58982 6554
rect 58982 6502 59028 6554
rect 58732 6500 58788 6502
rect 58812 6500 58868 6502
rect 58892 6500 58948 6502
rect 58972 6500 59028 6502
rect 58732 5466 58788 5468
rect 58812 5466 58868 5468
rect 58892 5466 58948 5468
rect 58972 5466 59028 5468
rect 58732 5414 58778 5466
rect 58778 5414 58788 5466
rect 58812 5414 58842 5466
rect 58842 5414 58854 5466
rect 58854 5414 58868 5466
rect 58892 5414 58906 5466
rect 58906 5414 58918 5466
rect 58918 5414 58948 5466
rect 58972 5414 58982 5466
rect 58982 5414 59028 5466
rect 58732 5412 58788 5414
rect 58812 5412 58868 5414
rect 58892 5412 58948 5414
rect 58972 5412 59028 5414
rect 58732 4378 58788 4380
rect 58812 4378 58868 4380
rect 58892 4378 58948 4380
rect 58972 4378 59028 4380
rect 58732 4326 58778 4378
rect 58778 4326 58788 4378
rect 58812 4326 58842 4378
rect 58842 4326 58854 4378
rect 58854 4326 58868 4378
rect 58892 4326 58906 4378
rect 58906 4326 58918 4378
rect 58918 4326 58948 4378
rect 58972 4326 58982 4378
rect 58982 4326 59028 4378
rect 58732 4324 58788 4326
rect 58812 4324 58868 4326
rect 58892 4324 58948 4326
rect 58972 4324 59028 4326
rect 58732 3290 58788 3292
rect 58812 3290 58868 3292
rect 58892 3290 58948 3292
rect 58972 3290 59028 3292
rect 58732 3238 58778 3290
rect 58778 3238 58788 3290
rect 58812 3238 58842 3290
rect 58842 3238 58854 3290
rect 58854 3238 58868 3290
rect 58892 3238 58906 3290
rect 58906 3238 58918 3290
rect 58918 3238 58948 3290
rect 58972 3238 58982 3290
rect 58982 3238 59028 3290
rect 58732 3236 58788 3238
rect 58812 3236 58868 3238
rect 58892 3236 58948 3238
rect 58972 3236 59028 3238
rect 58732 2202 58788 2204
rect 58812 2202 58868 2204
rect 58892 2202 58948 2204
rect 58972 2202 59028 2204
rect 58732 2150 58778 2202
rect 58778 2150 58788 2202
rect 58812 2150 58842 2202
rect 58842 2150 58854 2202
rect 58854 2150 58868 2202
rect 58892 2150 58906 2202
rect 58906 2150 58918 2202
rect 58918 2150 58948 2202
rect 58972 2150 58982 2202
rect 58982 2150 59028 2202
rect 58732 2148 58788 2150
rect 58812 2148 58868 2150
rect 58892 2148 58948 2150
rect 58972 2148 59028 2150
<< metal3 >>
rect 15390 21792 15706 21793
rect 15390 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15706 21792
rect 15390 21727 15706 21728
rect 29834 21792 30150 21793
rect 29834 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30150 21792
rect 29834 21727 30150 21728
rect 44278 21792 44594 21793
rect 44278 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44594 21792
rect 44278 21727 44594 21728
rect 58722 21792 59038 21793
rect 58722 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59038 21792
rect 58722 21727 59038 21728
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 22612 21248 22928 21249
rect 22612 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22928 21248
rect 22612 21183 22928 21184
rect 37056 21248 37372 21249
rect 37056 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37372 21248
rect 37056 21183 37372 21184
rect 51500 21248 51816 21249
rect 51500 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51816 21248
rect 51500 21183 51816 21184
rect 15390 20704 15706 20705
rect 15390 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15706 20704
rect 15390 20639 15706 20640
rect 29834 20704 30150 20705
rect 29834 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30150 20704
rect 29834 20639 30150 20640
rect 44278 20704 44594 20705
rect 44278 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44594 20704
rect 44278 20639 44594 20640
rect 58722 20704 59038 20705
rect 58722 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59038 20704
rect 58722 20639 59038 20640
rect 24669 20498 24735 20501
rect 52821 20498 52887 20501
rect 24669 20496 52887 20498
rect 24669 20440 24674 20496
rect 24730 20440 52826 20496
rect 52882 20440 52887 20496
rect 24669 20438 52887 20440
rect 24669 20435 24735 20438
rect 52821 20435 52887 20438
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 22612 20160 22928 20161
rect 22612 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22928 20160
rect 22612 20095 22928 20096
rect 37056 20160 37372 20161
rect 37056 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37372 20160
rect 37056 20095 37372 20096
rect 51500 20160 51816 20161
rect 51500 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51816 20160
rect 51500 20095 51816 20096
rect 40033 19818 40099 19821
rect 43713 19818 43779 19821
rect 40033 19816 43779 19818
rect 40033 19760 40038 19816
rect 40094 19760 43718 19816
rect 43774 19760 43779 19816
rect 40033 19758 43779 19760
rect 40033 19755 40099 19758
rect 43713 19755 43779 19758
rect 15390 19616 15706 19617
rect 15390 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15706 19616
rect 15390 19551 15706 19552
rect 29834 19616 30150 19617
rect 29834 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30150 19616
rect 29834 19551 30150 19552
rect 44278 19616 44594 19617
rect 44278 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44594 19616
rect 44278 19551 44594 19552
rect 58722 19616 59038 19617
rect 58722 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59038 19616
rect 58722 19551 59038 19552
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 22612 19072 22928 19073
rect 22612 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22928 19072
rect 22612 19007 22928 19008
rect 37056 19072 37372 19073
rect 37056 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37372 19072
rect 37056 19007 37372 19008
rect 51500 19072 51816 19073
rect 51500 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51816 19072
rect 51500 19007 51816 19008
rect 15390 18528 15706 18529
rect 15390 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15706 18528
rect 15390 18463 15706 18464
rect 29834 18528 30150 18529
rect 29834 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30150 18528
rect 29834 18463 30150 18464
rect 44278 18528 44594 18529
rect 44278 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44594 18528
rect 44278 18463 44594 18464
rect 58722 18528 59038 18529
rect 58722 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59038 18528
rect 58722 18463 59038 18464
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 22612 17984 22928 17985
rect 22612 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22928 17984
rect 22612 17919 22928 17920
rect 37056 17984 37372 17985
rect 37056 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37372 17984
rect 37056 17919 37372 17920
rect 51500 17984 51816 17985
rect 51500 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51816 17984
rect 51500 17919 51816 17920
rect 15390 17440 15706 17441
rect 15390 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15706 17440
rect 15390 17375 15706 17376
rect 29834 17440 30150 17441
rect 29834 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30150 17440
rect 29834 17375 30150 17376
rect 44278 17440 44594 17441
rect 44278 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44594 17440
rect 44278 17375 44594 17376
rect 58722 17440 59038 17441
rect 58722 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59038 17440
rect 58722 17375 59038 17376
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 22612 16896 22928 16897
rect 22612 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22928 16896
rect 22612 16831 22928 16832
rect 37056 16896 37372 16897
rect 37056 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37372 16896
rect 37056 16831 37372 16832
rect 51500 16896 51816 16897
rect 51500 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51816 16896
rect 51500 16831 51816 16832
rect 35433 16690 35499 16693
rect 35566 16690 35572 16692
rect 35433 16688 35572 16690
rect 35433 16632 35438 16688
rect 35494 16632 35572 16688
rect 35433 16630 35572 16632
rect 35433 16627 35499 16630
rect 35566 16628 35572 16630
rect 35636 16628 35642 16692
rect 15390 16352 15706 16353
rect 15390 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15706 16352
rect 15390 16287 15706 16288
rect 29834 16352 30150 16353
rect 29834 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30150 16352
rect 29834 16287 30150 16288
rect 44278 16352 44594 16353
rect 44278 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44594 16352
rect 44278 16287 44594 16288
rect 58722 16352 59038 16353
rect 58722 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59038 16352
rect 58722 16287 59038 16288
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 22612 15808 22928 15809
rect 22612 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22928 15808
rect 22612 15743 22928 15744
rect 37056 15808 37372 15809
rect 37056 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37372 15808
rect 37056 15743 37372 15744
rect 51500 15808 51816 15809
rect 51500 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51816 15808
rect 51500 15743 51816 15744
rect 15390 15264 15706 15265
rect 15390 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15706 15264
rect 15390 15199 15706 15200
rect 29834 15264 30150 15265
rect 29834 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30150 15264
rect 29834 15199 30150 15200
rect 44278 15264 44594 15265
rect 44278 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44594 15264
rect 44278 15199 44594 15200
rect 58722 15264 59038 15265
rect 58722 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59038 15264
rect 58722 15199 59038 15200
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 22612 14720 22928 14721
rect 22612 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22928 14720
rect 22612 14655 22928 14656
rect 37056 14720 37372 14721
rect 37056 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37372 14720
rect 37056 14655 37372 14656
rect 51500 14720 51816 14721
rect 51500 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51816 14720
rect 51500 14655 51816 14656
rect 15390 14176 15706 14177
rect 15390 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15706 14176
rect 15390 14111 15706 14112
rect 29834 14176 30150 14177
rect 29834 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30150 14176
rect 29834 14111 30150 14112
rect 44278 14176 44594 14177
rect 44278 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44594 14176
rect 44278 14111 44594 14112
rect 58722 14176 59038 14177
rect 58722 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59038 14176
rect 58722 14111 59038 14112
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 22612 13632 22928 13633
rect 22612 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22928 13632
rect 22612 13567 22928 13568
rect 37056 13632 37372 13633
rect 37056 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37372 13632
rect 37056 13567 37372 13568
rect 51500 13632 51816 13633
rect 51500 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51816 13632
rect 51500 13567 51816 13568
rect 35801 13426 35867 13429
rect 38837 13426 38903 13429
rect 35801 13424 38903 13426
rect 35801 13368 35806 13424
rect 35862 13368 38842 13424
rect 38898 13368 38903 13424
rect 35801 13366 38903 13368
rect 35801 13363 35867 13366
rect 38837 13363 38903 13366
rect 52269 13290 52335 13293
rect 56685 13290 56751 13293
rect 52269 13288 56751 13290
rect 52269 13232 52274 13288
rect 52330 13232 56690 13288
rect 56746 13232 56751 13288
rect 52269 13230 56751 13232
rect 52269 13227 52335 13230
rect 56685 13227 56751 13230
rect 15390 13088 15706 13089
rect 15390 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15706 13088
rect 15390 13023 15706 13024
rect 29834 13088 30150 13089
rect 29834 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30150 13088
rect 29834 13023 30150 13024
rect 44278 13088 44594 13089
rect 44278 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44594 13088
rect 44278 13023 44594 13024
rect 58722 13088 59038 13089
rect 58722 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59038 13088
rect 58722 13023 59038 13024
rect 31109 13018 31175 13021
rect 41045 13018 41111 13021
rect 31109 13016 41111 13018
rect 31109 12960 31114 13016
rect 31170 12960 41050 13016
rect 41106 12960 41111 13016
rect 31109 12958 41111 12960
rect 31109 12955 31175 12958
rect 41045 12955 41111 12958
rect 35525 12746 35591 12749
rect 40033 12746 40099 12749
rect 35525 12744 40099 12746
rect 35525 12688 35530 12744
rect 35586 12688 40038 12744
rect 40094 12688 40099 12744
rect 35525 12686 40099 12688
rect 35525 12683 35591 12686
rect 40033 12683 40099 12686
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 22612 12544 22928 12545
rect 22612 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22928 12544
rect 22612 12479 22928 12480
rect 37056 12544 37372 12545
rect 37056 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37372 12544
rect 37056 12479 37372 12480
rect 51500 12544 51816 12545
rect 51500 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51816 12544
rect 51500 12479 51816 12480
rect 15390 12000 15706 12001
rect 15390 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15706 12000
rect 15390 11935 15706 11936
rect 29834 12000 30150 12001
rect 29834 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30150 12000
rect 29834 11935 30150 11936
rect 44278 12000 44594 12001
rect 44278 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44594 12000
rect 44278 11935 44594 11936
rect 58722 12000 59038 12001
rect 58722 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59038 12000
rect 58722 11935 59038 11936
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 22612 11456 22928 11457
rect 22612 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22928 11456
rect 22612 11391 22928 11392
rect 37056 11456 37372 11457
rect 37056 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37372 11456
rect 37056 11391 37372 11392
rect 51500 11456 51816 11457
rect 51500 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51816 11456
rect 51500 11391 51816 11392
rect 15390 10912 15706 10913
rect 15390 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15706 10912
rect 15390 10847 15706 10848
rect 29834 10912 30150 10913
rect 29834 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30150 10912
rect 29834 10847 30150 10848
rect 44278 10912 44594 10913
rect 44278 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44594 10912
rect 44278 10847 44594 10848
rect 58722 10912 59038 10913
rect 58722 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59038 10912
rect 58722 10847 59038 10848
rect 19977 10706 20043 10709
rect 30649 10706 30715 10709
rect 19977 10704 30715 10706
rect 19977 10648 19982 10704
rect 20038 10648 30654 10704
rect 30710 10648 30715 10704
rect 19977 10646 30715 10648
rect 19977 10643 20043 10646
rect 30649 10643 30715 10646
rect 12985 10570 13051 10573
rect 52821 10570 52887 10573
rect 12985 10568 52887 10570
rect 12985 10512 12990 10568
rect 13046 10512 52826 10568
rect 52882 10512 52887 10568
rect 12985 10510 52887 10512
rect 12985 10507 13051 10510
rect 52821 10507 52887 10510
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 22612 10368 22928 10369
rect 22612 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22928 10368
rect 22612 10303 22928 10304
rect 37056 10368 37372 10369
rect 37056 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37372 10368
rect 37056 10303 37372 10304
rect 51500 10368 51816 10369
rect 51500 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51816 10368
rect 51500 10303 51816 10304
rect 22001 9890 22067 9893
rect 22185 9890 22251 9893
rect 27705 9890 27771 9893
rect 22001 9888 27771 9890
rect 22001 9832 22006 9888
rect 22062 9832 22190 9888
rect 22246 9832 27710 9888
rect 27766 9832 27771 9888
rect 22001 9830 27771 9832
rect 22001 9827 22067 9830
rect 22185 9827 22251 9830
rect 27705 9827 27771 9830
rect 15390 9824 15706 9825
rect 15390 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15706 9824
rect 15390 9759 15706 9760
rect 29834 9824 30150 9825
rect 29834 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30150 9824
rect 29834 9759 30150 9760
rect 44278 9824 44594 9825
rect 44278 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44594 9824
rect 44278 9759 44594 9760
rect 58722 9824 59038 9825
rect 58722 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59038 9824
rect 58722 9759 59038 9760
rect 9489 9482 9555 9485
rect 15285 9482 15351 9485
rect 9489 9480 15351 9482
rect 9489 9424 9494 9480
rect 9550 9424 15290 9480
rect 15346 9424 15351 9480
rect 9489 9422 15351 9424
rect 9489 9419 9555 9422
rect 15285 9419 15351 9422
rect 30741 9482 30807 9485
rect 38285 9482 38351 9485
rect 30741 9480 38351 9482
rect 30741 9424 30746 9480
rect 30802 9424 38290 9480
rect 38346 9424 38351 9480
rect 30741 9422 38351 9424
rect 30741 9419 30807 9422
rect 38285 9419 38351 9422
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 22612 9280 22928 9281
rect 22612 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22928 9280
rect 22612 9215 22928 9216
rect 37056 9280 37372 9281
rect 37056 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37372 9280
rect 37056 9215 37372 9216
rect 51500 9280 51816 9281
rect 51500 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51816 9280
rect 51500 9215 51816 9216
rect 10133 9074 10199 9077
rect 56041 9074 56107 9077
rect 10133 9072 56107 9074
rect 10133 9016 10138 9072
rect 10194 9016 56046 9072
rect 56102 9016 56107 9072
rect 10133 9014 56107 9016
rect 10133 9011 10199 9014
rect 56041 9011 56107 9014
rect 9213 8938 9279 8941
rect 56869 8938 56935 8941
rect 9213 8936 56935 8938
rect 9213 8880 9218 8936
rect 9274 8880 56874 8936
rect 56930 8880 56935 8936
rect 9213 8878 56935 8880
rect 9213 8875 9279 8878
rect 56869 8875 56935 8878
rect 53741 8802 53807 8805
rect 56869 8802 56935 8805
rect 53741 8800 56935 8802
rect 53741 8744 53746 8800
rect 53802 8744 56874 8800
rect 56930 8744 56935 8800
rect 53741 8742 56935 8744
rect 53741 8739 53807 8742
rect 56869 8739 56935 8742
rect 15390 8736 15706 8737
rect 15390 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15706 8736
rect 15390 8671 15706 8672
rect 29834 8736 30150 8737
rect 29834 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30150 8736
rect 29834 8671 30150 8672
rect 44278 8736 44594 8737
rect 44278 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44594 8736
rect 44278 8671 44594 8672
rect 58722 8736 59038 8737
rect 58722 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59038 8736
rect 58722 8671 59038 8672
rect 13353 8530 13419 8533
rect 52085 8530 52151 8533
rect 13353 8528 52151 8530
rect 13353 8472 13358 8528
rect 13414 8472 52090 8528
rect 52146 8472 52151 8528
rect 13353 8470 52151 8472
rect 13353 8467 13419 8470
rect 52085 8467 52151 8470
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 22612 8192 22928 8193
rect 22612 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22928 8192
rect 22612 8127 22928 8128
rect 37056 8192 37372 8193
rect 37056 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37372 8192
rect 37056 8127 37372 8128
rect 51500 8192 51816 8193
rect 51500 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51816 8192
rect 51500 8127 51816 8128
rect 15390 7648 15706 7649
rect 15390 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15706 7648
rect 15390 7583 15706 7584
rect 29834 7648 30150 7649
rect 29834 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30150 7648
rect 29834 7583 30150 7584
rect 44278 7648 44594 7649
rect 44278 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44594 7648
rect 44278 7583 44594 7584
rect 58722 7648 59038 7649
rect 58722 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59038 7648
rect 58722 7583 59038 7584
rect 35709 7442 35775 7445
rect 38469 7442 38535 7445
rect 35709 7440 38535 7442
rect 35709 7384 35714 7440
rect 35770 7384 38474 7440
rect 38530 7384 38535 7440
rect 35709 7382 38535 7384
rect 35709 7379 35775 7382
rect 38469 7379 38535 7382
rect 40677 7442 40743 7445
rect 44081 7442 44147 7445
rect 40677 7440 44147 7442
rect 40677 7384 40682 7440
rect 40738 7384 44086 7440
rect 44142 7384 44147 7440
rect 40677 7382 44147 7384
rect 40677 7379 40743 7382
rect 44081 7379 44147 7382
rect 7230 7244 7236 7308
rect 7300 7306 7306 7308
rect 8109 7306 8175 7309
rect 54201 7306 54267 7309
rect 7300 7304 54267 7306
rect 7300 7248 8114 7304
rect 8170 7248 54206 7304
rect 54262 7248 54267 7304
rect 7300 7246 54267 7248
rect 7300 7244 7306 7246
rect 8109 7243 8175 7246
rect 54201 7243 54267 7246
rect 40125 7170 40191 7173
rect 44817 7170 44883 7173
rect 40125 7168 44883 7170
rect 40125 7112 40130 7168
rect 40186 7112 44822 7168
rect 44878 7112 44883 7168
rect 40125 7110 44883 7112
rect 40125 7107 40191 7110
rect 44817 7107 44883 7110
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 22612 7104 22928 7105
rect 22612 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22928 7104
rect 22612 7039 22928 7040
rect 37056 7104 37372 7105
rect 37056 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37372 7104
rect 37056 7039 37372 7040
rect 51500 7104 51816 7105
rect 51500 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51816 7104
rect 51500 7039 51816 7040
rect 39849 7034 39915 7037
rect 44909 7034 44975 7037
rect 39849 7032 44975 7034
rect 39849 6976 39854 7032
rect 39910 6976 44914 7032
rect 44970 6976 44975 7032
rect 39849 6974 44975 6976
rect 39849 6971 39915 6974
rect 44909 6971 44975 6974
rect 55857 7034 55923 7037
rect 55990 7034 55996 7036
rect 55857 7032 55996 7034
rect 55857 6976 55862 7032
rect 55918 6976 55996 7032
rect 55857 6974 55996 6976
rect 55857 6971 55923 6974
rect 55990 6972 55996 6974
rect 56060 6972 56066 7036
rect 30189 6898 30255 6901
rect 31293 6898 31359 6901
rect 34973 6898 35039 6901
rect 30189 6896 35039 6898
rect 30189 6840 30194 6896
rect 30250 6840 31298 6896
rect 31354 6840 34978 6896
rect 35034 6840 35039 6896
rect 30189 6838 35039 6840
rect 30189 6835 30255 6838
rect 31293 6835 31359 6838
rect 34973 6835 35039 6838
rect 48773 6898 48839 6901
rect 55489 6898 55555 6901
rect 48773 6896 55555 6898
rect 48773 6840 48778 6896
rect 48834 6840 55494 6896
rect 55550 6840 55555 6896
rect 48773 6838 55555 6840
rect 48773 6835 48839 6838
rect 55489 6835 55555 6838
rect 15390 6560 15706 6561
rect 15390 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15706 6560
rect 15390 6495 15706 6496
rect 29834 6560 30150 6561
rect 29834 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30150 6560
rect 29834 6495 30150 6496
rect 44278 6560 44594 6561
rect 44278 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44594 6560
rect 44278 6495 44594 6496
rect 58722 6560 59038 6561
rect 58722 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59038 6560
rect 58722 6495 59038 6496
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 22612 6016 22928 6017
rect 22612 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22928 6016
rect 22612 5951 22928 5952
rect 37056 6016 37372 6017
rect 37056 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37372 6016
rect 37056 5951 37372 5952
rect 51500 6016 51816 6017
rect 51500 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51816 6016
rect 51500 5951 51816 5952
rect 44173 5674 44239 5677
rect 52729 5674 52795 5677
rect 44173 5672 52795 5674
rect 44173 5616 44178 5672
rect 44234 5616 52734 5672
rect 52790 5616 52795 5672
rect 44173 5614 52795 5616
rect 44173 5611 44239 5614
rect 52729 5611 52795 5614
rect 6177 5538 6243 5541
rect 7230 5538 7236 5540
rect 6177 5536 7236 5538
rect 6177 5480 6182 5536
rect 6238 5480 7236 5536
rect 6177 5478 7236 5480
rect 6177 5475 6243 5478
rect 7230 5476 7236 5478
rect 7300 5476 7306 5540
rect 15390 5472 15706 5473
rect 15390 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15706 5472
rect 15390 5407 15706 5408
rect 29834 5472 30150 5473
rect 29834 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30150 5472
rect 29834 5407 30150 5408
rect 44278 5472 44594 5473
rect 44278 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44594 5472
rect 44278 5407 44594 5408
rect 58722 5472 59038 5473
rect 58722 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59038 5472
rect 58722 5407 59038 5408
rect 5165 5266 5231 5269
rect 8753 5266 8819 5269
rect 5165 5264 8819 5266
rect 5165 5208 5170 5264
rect 5226 5208 8758 5264
rect 8814 5208 8819 5264
rect 5165 5206 8819 5208
rect 5165 5203 5231 5206
rect 8753 5203 8819 5206
rect 31477 5266 31543 5269
rect 34881 5266 34947 5269
rect 31477 5264 34947 5266
rect 31477 5208 31482 5264
rect 31538 5208 34886 5264
rect 34942 5208 34947 5264
rect 31477 5206 34947 5208
rect 31477 5203 31543 5206
rect 34881 5203 34947 5206
rect 6177 5130 6243 5133
rect 8845 5130 8911 5133
rect 6177 5128 8911 5130
rect 6177 5072 6182 5128
rect 6238 5072 8850 5128
rect 8906 5072 8911 5128
rect 6177 5070 8911 5072
rect 6177 5067 6243 5070
rect 8845 5067 8911 5070
rect 32305 4994 32371 4997
rect 32765 4994 32831 4997
rect 32305 4992 32831 4994
rect 32305 4936 32310 4992
rect 32366 4936 32770 4992
rect 32826 4936 32831 4992
rect 32305 4934 32831 4936
rect 32305 4931 32371 4934
rect 32765 4931 32831 4934
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 22612 4928 22928 4929
rect 22612 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22928 4928
rect 22612 4863 22928 4864
rect 37056 4928 37372 4929
rect 37056 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37372 4928
rect 37056 4863 37372 4864
rect 51500 4928 51816 4929
rect 51500 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51816 4928
rect 51500 4863 51816 4864
rect 35157 4586 35223 4589
rect 42885 4586 42951 4589
rect 35157 4584 42951 4586
rect 35157 4528 35162 4584
rect 35218 4528 42890 4584
rect 42946 4528 42951 4584
rect 35157 4526 42951 4528
rect 35157 4523 35223 4526
rect 42885 4523 42951 4526
rect 4245 4450 4311 4453
rect 9213 4450 9279 4453
rect 4245 4448 9279 4450
rect 4245 4392 4250 4448
rect 4306 4392 9218 4448
rect 9274 4392 9279 4448
rect 4245 4390 9279 4392
rect 4245 4387 4311 4390
rect 9213 4387 9279 4390
rect 15390 4384 15706 4385
rect 15390 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15706 4384
rect 15390 4319 15706 4320
rect 29834 4384 30150 4385
rect 29834 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30150 4384
rect 29834 4319 30150 4320
rect 44278 4384 44594 4385
rect 44278 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44594 4384
rect 44278 4319 44594 4320
rect 58722 4384 59038 4385
rect 58722 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59038 4384
rect 58722 4319 59038 4320
rect 10593 4178 10659 4181
rect 9630 4176 10659 4178
rect 9630 4120 10598 4176
rect 10654 4120 10659 4176
rect 9630 4118 10659 4120
rect 3785 4042 3851 4045
rect 9630 4042 9690 4118
rect 10593 4115 10659 4118
rect 30373 4178 30439 4181
rect 33225 4178 33291 4181
rect 30373 4176 33291 4178
rect 30373 4120 30378 4176
rect 30434 4120 33230 4176
rect 33286 4120 33291 4176
rect 30373 4118 33291 4120
rect 30373 4115 30439 4118
rect 33225 4115 33291 4118
rect 3785 4040 9690 4042
rect 3785 3984 3790 4040
rect 3846 3984 9690 4040
rect 3785 3982 9690 3984
rect 30281 4042 30347 4045
rect 35341 4042 35407 4045
rect 39941 4042 40007 4045
rect 41045 4042 41111 4045
rect 45093 4042 45159 4045
rect 30281 4040 45159 4042
rect 30281 3984 30286 4040
rect 30342 3984 35346 4040
rect 35402 3984 39946 4040
rect 40002 3984 41050 4040
rect 41106 3984 45098 4040
rect 45154 3984 45159 4040
rect 30281 3982 45159 3984
rect 3785 3979 3851 3982
rect 30281 3979 30347 3982
rect 35341 3979 35407 3982
rect 39941 3979 40007 3982
rect 41045 3979 41111 3982
rect 45093 3979 45159 3982
rect 55990 3980 55996 4044
rect 56060 4042 56066 4044
rect 56685 4042 56751 4045
rect 56060 4040 56751 4042
rect 56060 3984 56690 4040
rect 56746 3984 56751 4040
rect 56060 3982 56751 3984
rect 56060 3980 56066 3982
rect 56685 3979 56751 3982
rect 35566 3844 35572 3908
rect 35636 3906 35642 3908
rect 36813 3906 36879 3909
rect 35636 3904 36879 3906
rect 35636 3848 36818 3904
rect 36874 3848 36879 3904
rect 35636 3846 36879 3848
rect 35636 3844 35642 3846
rect 36813 3843 36879 3846
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 22612 3840 22928 3841
rect 22612 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22928 3840
rect 22612 3775 22928 3776
rect 37056 3840 37372 3841
rect 37056 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37372 3840
rect 37056 3775 37372 3776
rect 51500 3840 51816 3841
rect 51500 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51816 3840
rect 51500 3775 51816 3776
rect 4705 3770 4771 3773
rect 6729 3770 6795 3773
rect 4705 3768 6795 3770
rect 4705 3712 4710 3768
rect 4766 3712 6734 3768
rect 6790 3712 6795 3768
rect 4705 3710 6795 3712
rect 4705 3707 4771 3710
rect 6729 3707 6795 3710
rect 2129 3634 2195 3637
rect 4889 3634 4955 3637
rect 2129 3632 4955 3634
rect 2129 3576 2134 3632
rect 2190 3576 4894 3632
rect 4950 3576 4955 3632
rect 2129 3574 4955 3576
rect 2129 3571 2195 3574
rect 4889 3571 4955 3574
rect 7281 3634 7347 3637
rect 46933 3634 46999 3637
rect 7281 3632 46999 3634
rect 7281 3576 7286 3632
rect 7342 3576 46938 3632
rect 46994 3576 46999 3632
rect 7281 3574 46999 3576
rect 7281 3571 7347 3574
rect 46933 3571 46999 3574
rect 933 3498 999 3501
rect 29545 3498 29611 3501
rect 933 3496 29611 3498
rect 933 3440 938 3496
rect 994 3440 29550 3496
rect 29606 3440 29611 3496
rect 933 3438 29611 3440
rect 933 3435 999 3438
rect 29545 3435 29611 3438
rect 1669 3362 1735 3365
rect 6637 3362 6703 3365
rect 1669 3360 6703 3362
rect 1669 3304 1674 3360
rect 1730 3304 6642 3360
rect 6698 3304 6703 3360
rect 1669 3302 6703 3304
rect 1669 3299 1735 3302
rect 6637 3299 6703 3302
rect 16021 3362 16087 3365
rect 27337 3362 27403 3365
rect 16021 3360 27403 3362
rect 16021 3304 16026 3360
rect 16082 3304 27342 3360
rect 27398 3304 27403 3360
rect 16021 3302 27403 3304
rect 16021 3299 16087 3302
rect 27337 3299 27403 3302
rect 15390 3296 15706 3297
rect 15390 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15706 3296
rect 15390 3231 15706 3232
rect 29834 3296 30150 3297
rect 29834 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30150 3296
rect 29834 3231 30150 3232
rect 44278 3296 44594 3297
rect 44278 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44594 3296
rect 44278 3231 44594 3232
rect 58722 3296 59038 3297
rect 58722 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59038 3296
rect 58722 3231 59038 3232
rect 1853 3226 1919 3229
rect 6913 3226 6979 3229
rect 1853 3224 6979 3226
rect 1853 3168 1858 3224
rect 1914 3168 6918 3224
rect 6974 3168 6979 3224
rect 1853 3166 6979 3168
rect 1853 3163 1919 3166
rect 6913 3163 6979 3166
rect 27797 2954 27863 2957
rect 42885 2954 42951 2957
rect 27797 2952 42951 2954
rect 27797 2896 27802 2952
rect 27858 2896 42890 2952
rect 42946 2896 42951 2952
rect 27797 2894 42951 2896
rect 27797 2891 27863 2894
rect 42885 2891 42951 2894
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 22612 2752 22928 2753
rect 22612 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22928 2752
rect 22612 2687 22928 2688
rect 37056 2752 37372 2753
rect 37056 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37372 2752
rect 37056 2687 37372 2688
rect 51500 2752 51816 2753
rect 51500 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51816 2752
rect 51500 2687 51816 2688
rect 15390 2208 15706 2209
rect 15390 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15706 2208
rect 15390 2143 15706 2144
rect 29834 2208 30150 2209
rect 29834 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30150 2208
rect 29834 2143 30150 2144
rect 44278 2208 44594 2209
rect 44278 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44594 2208
rect 44278 2143 44594 2144
rect 58722 2208 59038 2209
rect 58722 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59038 2208
rect 58722 2143 59038 2144
<< via3 >>
rect 15396 21788 15460 21792
rect 15396 21732 15400 21788
rect 15400 21732 15456 21788
rect 15456 21732 15460 21788
rect 15396 21728 15460 21732
rect 15476 21788 15540 21792
rect 15476 21732 15480 21788
rect 15480 21732 15536 21788
rect 15536 21732 15540 21788
rect 15476 21728 15540 21732
rect 15556 21788 15620 21792
rect 15556 21732 15560 21788
rect 15560 21732 15616 21788
rect 15616 21732 15620 21788
rect 15556 21728 15620 21732
rect 15636 21788 15700 21792
rect 15636 21732 15640 21788
rect 15640 21732 15696 21788
rect 15696 21732 15700 21788
rect 15636 21728 15700 21732
rect 29840 21788 29904 21792
rect 29840 21732 29844 21788
rect 29844 21732 29900 21788
rect 29900 21732 29904 21788
rect 29840 21728 29904 21732
rect 29920 21788 29984 21792
rect 29920 21732 29924 21788
rect 29924 21732 29980 21788
rect 29980 21732 29984 21788
rect 29920 21728 29984 21732
rect 30000 21788 30064 21792
rect 30000 21732 30004 21788
rect 30004 21732 30060 21788
rect 30060 21732 30064 21788
rect 30000 21728 30064 21732
rect 30080 21788 30144 21792
rect 30080 21732 30084 21788
rect 30084 21732 30140 21788
rect 30140 21732 30144 21788
rect 30080 21728 30144 21732
rect 44284 21788 44348 21792
rect 44284 21732 44288 21788
rect 44288 21732 44344 21788
rect 44344 21732 44348 21788
rect 44284 21728 44348 21732
rect 44364 21788 44428 21792
rect 44364 21732 44368 21788
rect 44368 21732 44424 21788
rect 44424 21732 44428 21788
rect 44364 21728 44428 21732
rect 44444 21788 44508 21792
rect 44444 21732 44448 21788
rect 44448 21732 44504 21788
rect 44504 21732 44508 21788
rect 44444 21728 44508 21732
rect 44524 21788 44588 21792
rect 44524 21732 44528 21788
rect 44528 21732 44584 21788
rect 44584 21732 44588 21788
rect 44524 21728 44588 21732
rect 58728 21788 58792 21792
rect 58728 21732 58732 21788
rect 58732 21732 58788 21788
rect 58788 21732 58792 21788
rect 58728 21728 58792 21732
rect 58808 21788 58872 21792
rect 58808 21732 58812 21788
rect 58812 21732 58868 21788
rect 58868 21732 58872 21788
rect 58808 21728 58872 21732
rect 58888 21788 58952 21792
rect 58888 21732 58892 21788
rect 58892 21732 58948 21788
rect 58948 21732 58952 21788
rect 58888 21728 58952 21732
rect 58968 21788 59032 21792
rect 58968 21732 58972 21788
rect 58972 21732 59028 21788
rect 59028 21732 59032 21788
rect 58968 21728 59032 21732
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 22618 21244 22682 21248
rect 22618 21188 22622 21244
rect 22622 21188 22678 21244
rect 22678 21188 22682 21244
rect 22618 21184 22682 21188
rect 22698 21244 22762 21248
rect 22698 21188 22702 21244
rect 22702 21188 22758 21244
rect 22758 21188 22762 21244
rect 22698 21184 22762 21188
rect 22778 21244 22842 21248
rect 22778 21188 22782 21244
rect 22782 21188 22838 21244
rect 22838 21188 22842 21244
rect 22778 21184 22842 21188
rect 22858 21244 22922 21248
rect 22858 21188 22862 21244
rect 22862 21188 22918 21244
rect 22918 21188 22922 21244
rect 22858 21184 22922 21188
rect 37062 21244 37126 21248
rect 37062 21188 37066 21244
rect 37066 21188 37122 21244
rect 37122 21188 37126 21244
rect 37062 21184 37126 21188
rect 37142 21244 37206 21248
rect 37142 21188 37146 21244
rect 37146 21188 37202 21244
rect 37202 21188 37206 21244
rect 37142 21184 37206 21188
rect 37222 21244 37286 21248
rect 37222 21188 37226 21244
rect 37226 21188 37282 21244
rect 37282 21188 37286 21244
rect 37222 21184 37286 21188
rect 37302 21244 37366 21248
rect 37302 21188 37306 21244
rect 37306 21188 37362 21244
rect 37362 21188 37366 21244
rect 37302 21184 37366 21188
rect 51506 21244 51570 21248
rect 51506 21188 51510 21244
rect 51510 21188 51566 21244
rect 51566 21188 51570 21244
rect 51506 21184 51570 21188
rect 51586 21244 51650 21248
rect 51586 21188 51590 21244
rect 51590 21188 51646 21244
rect 51646 21188 51650 21244
rect 51586 21184 51650 21188
rect 51666 21244 51730 21248
rect 51666 21188 51670 21244
rect 51670 21188 51726 21244
rect 51726 21188 51730 21244
rect 51666 21184 51730 21188
rect 51746 21244 51810 21248
rect 51746 21188 51750 21244
rect 51750 21188 51806 21244
rect 51806 21188 51810 21244
rect 51746 21184 51810 21188
rect 15396 20700 15460 20704
rect 15396 20644 15400 20700
rect 15400 20644 15456 20700
rect 15456 20644 15460 20700
rect 15396 20640 15460 20644
rect 15476 20700 15540 20704
rect 15476 20644 15480 20700
rect 15480 20644 15536 20700
rect 15536 20644 15540 20700
rect 15476 20640 15540 20644
rect 15556 20700 15620 20704
rect 15556 20644 15560 20700
rect 15560 20644 15616 20700
rect 15616 20644 15620 20700
rect 15556 20640 15620 20644
rect 15636 20700 15700 20704
rect 15636 20644 15640 20700
rect 15640 20644 15696 20700
rect 15696 20644 15700 20700
rect 15636 20640 15700 20644
rect 29840 20700 29904 20704
rect 29840 20644 29844 20700
rect 29844 20644 29900 20700
rect 29900 20644 29904 20700
rect 29840 20640 29904 20644
rect 29920 20700 29984 20704
rect 29920 20644 29924 20700
rect 29924 20644 29980 20700
rect 29980 20644 29984 20700
rect 29920 20640 29984 20644
rect 30000 20700 30064 20704
rect 30000 20644 30004 20700
rect 30004 20644 30060 20700
rect 30060 20644 30064 20700
rect 30000 20640 30064 20644
rect 30080 20700 30144 20704
rect 30080 20644 30084 20700
rect 30084 20644 30140 20700
rect 30140 20644 30144 20700
rect 30080 20640 30144 20644
rect 44284 20700 44348 20704
rect 44284 20644 44288 20700
rect 44288 20644 44344 20700
rect 44344 20644 44348 20700
rect 44284 20640 44348 20644
rect 44364 20700 44428 20704
rect 44364 20644 44368 20700
rect 44368 20644 44424 20700
rect 44424 20644 44428 20700
rect 44364 20640 44428 20644
rect 44444 20700 44508 20704
rect 44444 20644 44448 20700
rect 44448 20644 44504 20700
rect 44504 20644 44508 20700
rect 44444 20640 44508 20644
rect 44524 20700 44588 20704
rect 44524 20644 44528 20700
rect 44528 20644 44584 20700
rect 44584 20644 44588 20700
rect 44524 20640 44588 20644
rect 58728 20700 58792 20704
rect 58728 20644 58732 20700
rect 58732 20644 58788 20700
rect 58788 20644 58792 20700
rect 58728 20640 58792 20644
rect 58808 20700 58872 20704
rect 58808 20644 58812 20700
rect 58812 20644 58868 20700
rect 58868 20644 58872 20700
rect 58808 20640 58872 20644
rect 58888 20700 58952 20704
rect 58888 20644 58892 20700
rect 58892 20644 58948 20700
rect 58948 20644 58952 20700
rect 58888 20640 58952 20644
rect 58968 20700 59032 20704
rect 58968 20644 58972 20700
rect 58972 20644 59028 20700
rect 59028 20644 59032 20700
rect 58968 20640 59032 20644
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 22618 20156 22682 20160
rect 22618 20100 22622 20156
rect 22622 20100 22678 20156
rect 22678 20100 22682 20156
rect 22618 20096 22682 20100
rect 22698 20156 22762 20160
rect 22698 20100 22702 20156
rect 22702 20100 22758 20156
rect 22758 20100 22762 20156
rect 22698 20096 22762 20100
rect 22778 20156 22842 20160
rect 22778 20100 22782 20156
rect 22782 20100 22838 20156
rect 22838 20100 22842 20156
rect 22778 20096 22842 20100
rect 22858 20156 22922 20160
rect 22858 20100 22862 20156
rect 22862 20100 22918 20156
rect 22918 20100 22922 20156
rect 22858 20096 22922 20100
rect 37062 20156 37126 20160
rect 37062 20100 37066 20156
rect 37066 20100 37122 20156
rect 37122 20100 37126 20156
rect 37062 20096 37126 20100
rect 37142 20156 37206 20160
rect 37142 20100 37146 20156
rect 37146 20100 37202 20156
rect 37202 20100 37206 20156
rect 37142 20096 37206 20100
rect 37222 20156 37286 20160
rect 37222 20100 37226 20156
rect 37226 20100 37282 20156
rect 37282 20100 37286 20156
rect 37222 20096 37286 20100
rect 37302 20156 37366 20160
rect 37302 20100 37306 20156
rect 37306 20100 37362 20156
rect 37362 20100 37366 20156
rect 37302 20096 37366 20100
rect 51506 20156 51570 20160
rect 51506 20100 51510 20156
rect 51510 20100 51566 20156
rect 51566 20100 51570 20156
rect 51506 20096 51570 20100
rect 51586 20156 51650 20160
rect 51586 20100 51590 20156
rect 51590 20100 51646 20156
rect 51646 20100 51650 20156
rect 51586 20096 51650 20100
rect 51666 20156 51730 20160
rect 51666 20100 51670 20156
rect 51670 20100 51726 20156
rect 51726 20100 51730 20156
rect 51666 20096 51730 20100
rect 51746 20156 51810 20160
rect 51746 20100 51750 20156
rect 51750 20100 51806 20156
rect 51806 20100 51810 20156
rect 51746 20096 51810 20100
rect 15396 19612 15460 19616
rect 15396 19556 15400 19612
rect 15400 19556 15456 19612
rect 15456 19556 15460 19612
rect 15396 19552 15460 19556
rect 15476 19612 15540 19616
rect 15476 19556 15480 19612
rect 15480 19556 15536 19612
rect 15536 19556 15540 19612
rect 15476 19552 15540 19556
rect 15556 19612 15620 19616
rect 15556 19556 15560 19612
rect 15560 19556 15616 19612
rect 15616 19556 15620 19612
rect 15556 19552 15620 19556
rect 15636 19612 15700 19616
rect 15636 19556 15640 19612
rect 15640 19556 15696 19612
rect 15696 19556 15700 19612
rect 15636 19552 15700 19556
rect 29840 19612 29904 19616
rect 29840 19556 29844 19612
rect 29844 19556 29900 19612
rect 29900 19556 29904 19612
rect 29840 19552 29904 19556
rect 29920 19612 29984 19616
rect 29920 19556 29924 19612
rect 29924 19556 29980 19612
rect 29980 19556 29984 19612
rect 29920 19552 29984 19556
rect 30000 19612 30064 19616
rect 30000 19556 30004 19612
rect 30004 19556 30060 19612
rect 30060 19556 30064 19612
rect 30000 19552 30064 19556
rect 30080 19612 30144 19616
rect 30080 19556 30084 19612
rect 30084 19556 30140 19612
rect 30140 19556 30144 19612
rect 30080 19552 30144 19556
rect 44284 19612 44348 19616
rect 44284 19556 44288 19612
rect 44288 19556 44344 19612
rect 44344 19556 44348 19612
rect 44284 19552 44348 19556
rect 44364 19612 44428 19616
rect 44364 19556 44368 19612
rect 44368 19556 44424 19612
rect 44424 19556 44428 19612
rect 44364 19552 44428 19556
rect 44444 19612 44508 19616
rect 44444 19556 44448 19612
rect 44448 19556 44504 19612
rect 44504 19556 44508 19612
rect 44444 19552 44508 19556
rect 44524 19612 44588 19616
rect 44524 19556 44528 19612
rect 44528 19556 44584 19612
rect 44584 19556 44588 19612
rect 44524 19552 44588 19556
rect 58728 19612 58792 19616
rect 58728 19556 58732 19612
rect 58732 19556 58788 19612
rect 58788 19556 58792 19612
rect 58728 19552 58792 19556
rect 58808 19612 58872 19616
rect 58808 19556 58812 19612
rect 58812 19556 58868 19612
rect 58868 19556 58872 19612
rect 58808 19552 58872 19556
rect 58888 19612 58952 19616
rect 58888 19556 58892 19612
rect 58892 19556 58948 19612
rect 58948 19556 58952 19612
rect 58888 19552 58952 19556
rect 58968 19612 59032 19616
rect 58968 19556 58972 19612
rect 58972 19556 59028 19612
rect 59028 19556 59032 19612
rect 58968 19552 59032 19556
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 22618 19068 22682 19072
rect 22618 19012 22622 19068
rect 22622 19012 22678 19068
rect 22678 19012 22682 19068
rect 22618 19008 22682 19012
rect 22698 19068 22762 19072
rect 22698 19012 22702 19068
rect 22702 19012 22758 19068
rect 22758 19012 22762 19068
rect 22698 19008 22762 19012
rect 22778 19068 22842 19072
rect 22778 19012 22782 19068
rect 22782 19012 22838 19068
rect 22838 19012 22842 19068
rect 22778 19008 22842 19012
rect 22858 19068 22922 19072
rect 22858 19012 22862 19068
rect 22862 19012 22918 19068
rect 22918 19012 22922 19068
rect 22858 19008 22922 19012
rect 37062 19068 37126 19072
rect 37062 19012 37066 19068
rect 37066 19012 37122 19068
rect 37122 19012 37126 19068
rect 37062 19008 37126 19012
rect 37142 19068 37206 19072
rect 37142 19012 37146 19068
rect 37146 19012 37202 19068
rect 37202 19012 37206 19068
rect 37142 19008 37206 19012
rect 37222 19068 37286 19072
rect 37222 19012 37226 19068
rect 37226 19012 37282 19068
rect 37282 19012 37286 19068
rect 37222 19008 37286 19012
rect 37302 19068 37366 19072
rect 37302 19012 37306 19068
rect 37306 19012 37362 19068
rect 37362 19012 37366 19068
rect 37302 19008 37366 19012
rect 51506 19068 51570 19072
rect 51506 19012 51510 19068
rect 51510 19012 51566 19068
rect 51566 19012 51570 19068
rect 51506 19008 51570 19012
rect 51586 19068 51650 19072
rect 51586 19012 51590 19068
rect 51590 19012 51646 19068
rect 51646 19012 51650 19068
rect 51586 19008 51650 19012
rect 51666 19068 51730 19072
rect 51666 19012 51670 19068
rect 51670 19012 51726 19068
rect 51726 19012 51730 19068
rect 51666 19008 51730 19012
rect 51746 19068 51810 19072
rect 51746 19012 51750 19068
rect 51750 19012 51806 19068
rect 51806 19012 51810 19068
rect 51746 19008 51810 19012
rect 15396 18524 15460 18528
rect 15396 18468 15400 18524
rect 15400 18468 15456 18524
rect 15456 18468 15460 18524
rect 15396 18464 15460 18468
rect 15476 18524 15540 18528
rect 15476 18468 15480 18524
rect 15480 18468 15536 18524
rect 15536 18468 15540 18524
rect 15476 18464 15540 18468
rect 15556 18524 15620 18528
rect 15556 18468 15560 18524
rect 15560 18468 15616 18524
rect 15616 18468 15620 18524
rect 15556 18464 15620 18468
rect 15636 18524 15700 18528
rect 15636 18468 15640 18524
rect 15640 18468 15696 18524
rect 15696 18468 15700 18524
rect 15636 18464 15700 18468
rect 29840 18524 29904 18528
rect 29840 18468 29844 18524
rect 29844 18468 29900 18524
rect 29900 18468 29904 18524
rect 29840 18464 29904 18468
rect 29920 18524 29984 18528
rect 29920 18468 29924 18524
rect 29924 18468 29980 18524
rect 29980 18468 29984 18524
rect 29920 18464 29984 18468
rect 30000 18524 30064 18528
rect 30000 18468 30004 18524
rect 30004 18468 30060 18524
rect 30060 18468 30064 18524
rect 30000 18464 30064 18468
rect 30080 18524 30144 18528
rect 30080 18468 30084 18524
rect 30084 18468 30140 18524
rect 30140 18468 30144 18524
rect 30080 18464 30144 18468
rect 44284 18524 44348 18528
rect 44284 18468 44288 18524
rect 44288 18468 44344 18524
rect 44344 18468 44348 18524
rect 44284 18464 44348 18468
rect 44364 18524 44428 18528
rect 44364 18468 44368 18524
rect 44368 18468 44424 18524
rect 44424 18468 44428 18524
rect 44364 18464 44428 18468
rect 44444 18524 44508 18528
rect 44444 18468 44448 18524
rect 44448 18468 44504 18524
rect 44504 18468 44508 18524
rect 44444 18464 44508 18468
rect 44524 18524 44588 18528
rect 44524 18468 44528 18524
rect 44528 18468 44584 18524
rect 44584 18468 44588 18524
rect 44524 18464 44588 18468
rect 58728 18524 58792 18528
rect 58728 18468 58732 18524
rect 58732 18468 58788 18524
rect 58788 18468 58792 18524
rect 58728 18464 58792 18468
rect 58808 18524 58872 18528
rect 58808 18468 58812 18524
rect 58812 18468 58868 18524
rect 58868 18468 58872 18524
rect 58808 18464 58872 18468
rect 58888 18524 58952 18528
rect 58888 18468 58892 18524
rect 58892 18468 58948 18524
rect 58948 18468 58952 18524
rect 58888 18464 58952 18468
rect 58968 18524 59032 18528
rect 58968 18468 58972 18524
rect 58972 18468 59028 18524
rect 59028 18468 59032 18524
rect 58968 18464 59032 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 22618 17980 22682 17984
rect 22618 17924 22622 17980
rect 22622 17924 22678 17980
rect 22678 17924 22682 17980
rect 22618 17920 22682 17924
rect 22698 17980 22762 17984
rect 22698 17924 22702 17980
rect 22702 17924 22758 17980
rect 22758 17924 22762 17980
rect 22698 17920 22762 17924
rect 22778 17980 22842 17984
rect 22778 17924 22782 17980
rect 22782 17924 22838 17980
rect 22838 17924 22842 17980
rect 22778 17920 22842 17924
rect 22858 17980 22922 17984
rect 22858 17924 22862 17980
rect 22862 17924 22918 17980
rect 22918 17924 22922 17980
rect 22858 17920 22922 17924
rect 37062 17980 37126 17984
rect 37062 17924 37066 17980
rect 37066 17924 37122 17980
rect 37122 17924 37126 17980
rect 37062 17920 37126 17924
rect 37142 17980 37206 17984
rect 37142 17924 37146 17980
rect 37146 17924 37202 17980
rect 37202 17924 37206 17980
rect 37142 17920 37206 17924
rect 37222 17980 37286 17984
rect 37222 17924 37226 17980
rect 37226 17924 37282 17980
rect 37282 17924 37286 17980
rect 37222 17920 37286 17924
rect 37302 17980 37366 17984
rect 37302 17924 37306 17980
rect 37306 17924 37362 17980
rect 37362 17924 37366 17980
rect 37302 17920 37366 17924
rect 51506 17980 51570 17984
rect 51506 17924 51510 17980
rect 51510 17924 51566 17980
rect 51566 17924 51570 17980
rect 51506 17920 51570 17924
rect 51586 17980 51650 17984
rect 51586 17924 51590 17980
rect 51590 17924 51646 17980
rect 51646 17924 51650 17980
rect 51586 17920 51650 17924
rect 51666 17980 51730 17984
rect 51666 17924 51670 17980
rect 51670 17924 51726 17980
rect 51726 17924 51730 17980
rect 51666 17920 51730 17924
rect 51746 17980 51810 17984
rect 51746 17924 51750 17980
rect 51750 17924 51806 17980
rect 51806 17924 51810 17980
rect 51746 17920 51810 17924
rect 15396 17436 15460 17440
rect 15396 17380 15400 17436
rect 15400 17380 15456 17436
rect 15456 17380 15460 17436
rect 15396 17376 15460 17380
rect 15476 17436 15540 17440
rect 15476 17380 15480 17436
rect 15480 17380 15536 17436
rect 15536 17380 15540 17436
rect 15476 17376 15540 17380
rect 15556 17436 15620 17440
rect 15556 17380 15560 17436
rect 15560 17380 15616 17436
rect 15616 17380 15620 17436
rect 15556 17376 15620 17380
rect 15636 17436 15700 17440
rect 15636 17380 15640 17436
rect 15640 17380 15696 17436
rect 15696 17380 15700 17436
rect 15636 17376 15700 17380
rect 29840 17436 29904 17440
rect 29840 17380 29844 17436
rect 29844 17380 29900 17436
rect 29900 17380 29904 17436
rect 29840 17376 29904 17380
rect 29920 17436 29984 17440
rect 29920 17380 29924 17436
rect 29924 17380 29980 17436
rect 29980 17380 29984 17436
rect 29920 17376 29984 17380
rect 30000 17436 30064 17440
rect 30000 17380 30004 17436
rect 30004 17380 30060 17436
rect 30060 17380 30064 17436
rect 30000 17376 30064 17380
rect 30080 17436 30144 17440
rect 30080 17380 30084 17436
rect 30084 17380 30140 17436
rect 30140 17380 30144 17436
rect 30080 17376 30144 17380
rect 44284 17436 44348 17440
rect 44284 17380 44288 17436
rect 44288 17380 44344 17436
rect 44344 17380 44348 17436
rect 44284 17376 44348 17380
rect 44364 17436 44428 17440
rect 44364 17380 44368 17436
rect 44368 17380 44424 17436
rect 44424 17380 44428 17436
rect 44364 17376 44428 17380
rect 44444 17436 44508 17440
rect 44444 17380 44448 17436
rect 44448 17380 44504 17436
rect 44504 17380 44508 17436
rect 44444 17376 44508 17380
rect 44524 17436 44588 17440
rect 44524 17380 44528 17436
rect 44528 17380 44584 17436
rect 44584 17380 44588 17436
rect 44524 17376 44588 17380
rect 58728 17436 58792 17440
rect 58728 17380 58732 17436
rect 58732 17380 58788 17436
rect 58788 17380 58792 17436
rect 58728 17376 58792 17380
rect 58808 17436 58872 17440
rect 58808 17380 58812 17436
rect 58812 17380 58868 17436
rect 58868 17380 58872 17436
rect 58808 17376 58872 17380
rect 58888 17436 58952 17440
rect 58888 17380 58892 17436
rect 58892 17380 58948 17436
rect 58948 17380 58952 17436
rect 58888 17376 58952 17380
rect 58968 17436 59032 17440
rect 58968 17380 58972 17436
rect 58972 17380 59028 17436
rect 59028 17380 59032 17436
rect 58968 17376 59032 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 22618 16892 22682 16896
rect 22618 16836 22622 16892
rect 22622 16836 22678 16892
rect 22678 16836 22682 16892
rect 22618 16832 22682 16836
rect 22698 16892 22762 16896
rect 22698 16836 22702 16892
rect 22702 16836 22758 16892
rect 22758 16836 22762 16892
rect 22698 16832 22762 16836
rect 22778 16892 22842 16896
rect 22778 16836 22782 16892
rect 22782 16836 22838 16892
rect 22838 16836 22842 16892
rect 22778 16832 22842 16836
rect 22858 16892 22922 16896
rect 22858 16836 22862 16892
rect 22862 16836 22918 16892
rect 22918 16836 22922 16892
rect 22858 16832 22922 16836
rect 37062 16892 37126 16896
rect 37062 16836 37066 16892
rect 37066 16836 37122 16892
rect 37122 16836 37126 16892
rect 37062 16832 37126 16836
rect 37142 16892 37206 16896
rect 37142 16836 37146 16892
rect 37146 16836 37202 16892
rect 37202 16836 37206 16892
rect 37142 16832 37206 16836
rect 37222 16892 37286 16896
rect 37222 16836 37226 16892
rect 37226 16836 37282 16892
rect 37282 16836 37286 16892
rect 37222 16832 37286 16836
rect 37302 16892 37366 16896
rect 37302 16836 37306 16892
rect 37306 16836 37362 16892
rect 37362 16836 37366 16892
rect 37302 16832 37366 16836
rect 51506 16892 51570 16896
rect 51506 16836 51510 16892
rect 51510 16836 51566 16892
rect 51566 16836 51570 16892
rect 51506 16832 51570 16836
rect 51586 16892 51650 16896
rect 51586 16836 51590 16892
rect 51590 16836 51646 16892
rect 51646 16836 51650 16892
rect 51586 16832 51650 16836
rect 51666 16892 51730 16896
rect 51666 16836 51670 16892
rect 51670 16836 51726 16892
rect 51726 16836 51730 16892
rect 51666 16832 51730 16836
rect 51746 16892 51810 16896
rect 51746 16836 51750 16892
rect 51750 16836 51806 16892
rect 51806 16836 51810 16892
rect 51746 16832 51810 16836
rect 35572 16628 35636 16692
rect 15396 16348 15460 16352
rect 15396 16292 15400 16348
rect 15400 16292 15456 16348
rect 15456 16292 15460 16348
rect 15396 16288 15460 16292
rect 15476 16348 15540 16352
rect 15476 16292 15480 16348
rect 15480 16292 15536 16348
rect 15536 16292 15540 16348
rect 15476 16288 15540 16292
rect 15556 16348 15620 16352
rect 15556 16292 15560 16348
rect 15560 16292 15616 16348
rect 15616 16292 15620 16348
rect 15556 16288 15620 16292
rect 15636 16348 15700 16352
rect 15636 16292 15640 16348
rect 15640 16292 15696 16348
rect 15696 16292 15700 16348
rect 15636 16288 15700 16292
rect 29840 16348 29904 16352
rect 29840 16292 29844 16348
rect 29844 16292 29900 16348
rect 29900 16292 29904 16348
rect 29840 16288 29904 16292
rect 29920 16348 29984 16352
rect 29920 16292 29924 16348
rect 29924 16292 29980 16348
rect 29980 16292 29984 16348
rect 29920 16288 29984 16292
rect 30000 16348 30064 16352
rect 30000 16292 30004 16348
rect 30004 16292 30060 16348
rect 30060 16292 30064 16348
rect 30000 16288 30064 16292
rect 30080 16348 30144 16352
rect 30080 16292 30084 16348
rect 30084 16292 30140 16348
rect 30140 16292 30144 16348
rect 30080 16288 30144 16292
rect 44284 16348 44348 16352
rect 44284 16292 44288 16348
rect 44288 16292 44344 16348
rect 44344 16292 44348 16348
rect 44284 16288 44348 16292
rect 44364 16348 44428 16352
rect 44364 16292 44368 16348
rect 44368 16292 44424 16348
rect 44424 16292 44428 16348
rect 44364 16288 44428 16292
rect 44444 16348 44508 16352
rect 44444 16292 44448 16348
rect 44448 16292 44504 16348
rect 44504 16292 44508 16348
rect 44444 16288 44508 16292
rect 44524 16348 44588 16352
rect 44524 16292 44528 16348
rect 44528 16292 44584 16348
rect 44584 16292 44588 16348
rect 44524 16288 44588 16292
rect 58728 16348 58792 16352
rect 58728 16292 58732 16348
rect 58732 16292 58788 16348
rect 58788 16292 58792 16348
rect 58728 16288 58792 16292
rect 58808 16348 58872 16352
rect 58808 16292 58812 16348
rect 58812 16292 58868 16348
rect 58868 16292 58872 16348
rect 58808 16288 58872 16292
rect 58888 16348 58952 16352
rect 58888 16292 58892 16348
rect 58892 16292 58948 16348
rect 58948 16292 58952 16348
rect 58888 16288 58952 16292
rect 58968 16348 59032 16352
rect 58968 16292 58972 16348
rect 58972 16292 59028 16348
rect 59028 16292 59032 16348
rect 58968 16288 59032 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 22618 15804 22682 15808
rect 22618 15748 22622 15804
rect 22622 15748 22678 15804
rect 22678 15748 22682 15804
rect 22618 15744 22682 15748
rect 22698 15804 22762 15808
rect 22698 15748 22702 15804
rect 22702 15748 22758 15804
rect 22758 15748 22762 15804
rect 22698 15744 22762 15748
rect 22778 15804 22842 15808
rect 22778 15748 22782 15804
rect 22782 15748 22838 15804
rect 22838 15748 22842 15804
rect 22778 15744 22842 15748
rect 22858 15804 22922 15808
rect 22858 15748 22862 15804
rect 22862 15748 22918 15804
rect 22918 15748 22922 15804
rect 22858 15744 22922 15748
rect 37062 15804 37126 15808
rect 37062 15748 37066 15804
rect 37066 15748 37122 15804
rect 37122 15748 37126 15804
rect 37062 15744 37126 15748
rect 37142 15804 37206 15808
rect 37142 15748 37146 15804
rect 37146 15748 37202 15804
rect 37202 15748 37206 15804
rect 37142 15744 37206 15748
rect 37222 15804 37286 15808
rect 37222 15748 37226 15804
rect 37226 15748 37282 15804
rect 37282 15748 37286 15804
rect 37222 15744 37286 15748
rect 37302 15804 37366 15808
rect 37302 15748 37306 15804
rect 37306 15748 37362 15804
rect 37362 15748 37366 15804
rect 37302 15744 37366 15748
rect 51506 15804 51570 15808
rect 51506 15748 51510 15804
rect 51510 15748 51566 15804
rect 51566 15748 51570 15804
rect 51506 15744 51570 15748
rect 51586 15804 51650 15808
rect 51586 15748 51590 15804
rect 51590 15748 51646 15804
rect 51646 15748 51650 15804
rect 51586 15744 51650 15748
rect 51666 15804 51730 15808
rect 51666 15748 51670 15804
rect 51670 15748 51726 15804
rect 51726 15748 51730 15804
rect 51666 15744 51730 15748
rect 51746 15804 51810 15808
rect 51746 15748 51750 15804
rect 51750 15748 51806 15804
rect 51806 15748 51810 15804
rect 51746 15744 51810 15748
rect 15396 15260 15460 15264
rect 15396 15204 15400 15260
rect 15400 15204 15456 15260
rect 15456 15204 15460 15260
rect 15396 15200 15460 15204
rect 15476 15260 15540 15264
rect 15476 15204 15480 15260
rect 15480 15204 15536 15260
rect 15536 15204 15540 15260
rect 15476 15200 15540 15204
rect 15556 15260 15620 15264
rect 15556 15204 15560 15260
rect 15560 15204 15616 15260
rect 15616 15204 15620 15260
rect 15556 15200 15620 15204
rect 15636 15260 15700 15264
rect 15636 15204 15640 15260
rect 15640 15204 15696 15260
rect 15696 15204 15700 15260
rect 15636 15200 15700 15204
rect 29840 15260 29904 15264
rect 29840 15204 29844 15260
rect 29844 15204 29900 15260
rect 29900 15204 29904 15260
rect 29840 15200 29904 15204
rect 29920 15260 29984 15264
rect 29920 15204 29924 15260
rect 29924 15204 29980 15260
rect 29980 15204 29984 15260
rect 29920 15200 29984 15204
rect 30000 15260 30064 15264
rect 30000 15204 30004 15260
rect 30004 15204 30060 15260
rect 30060 15204 30064 15260
rect 30000 15200 30064 15204
rect 30080 15260 30144 15264
rect 30080 15204 30084 15260
rect 30084 15204 30140 15260
rect 30140 15204 30144 15260
rect 30080 15200 30144 15204
rect 44284 15260 44348 15264
rect 44284 15204 44288 15260
rect 44288 15204 44344 15260
rect 44344 15204 44348 15260
rect 44284 15200 44348 15204
rect 44364 15260 44428 15264
rect 44364 15204 44368 15260
rect 44368 15204 44424 15260
rect 44424 15204 44428 15260
rect 44364 15200 44428 15204
rect 44444 15260 44508 15264
rect 44444 15204 44448 15260
rect 44448 15204 44504 15260
rect 44504 15204 44508 15260
rect 44444 15200 44508 15204
rect 44524 15260 44588 15264
rect 44524 15204 44528 15260
rect 44528 15204 44584 15260
rect 44584 15204 44588 15260
rect 44524 15200 44588 15204
rect 58728 15260 58792 15264
rect 58728 15204 58732 15260
rect 58732 15204 58788 15260
rect 58788 15204 58792 15260
rect 58728 15200 58792 15204
rect 58808 15260 58872 15264
rect 58808 15204 58812 15260
rect 58812 15204 58868 15260
rect 58868 15204 58872 15260
rect 58808 15200 58872 15204
rect 58888 15260 58952 15264
rect 58888 15204 58892 15260
rect 58892 15204 58948 15260
rect 58948 15204 58952 15260
rect 58888 15200 58952 15204
rect 58968 15260 59032 15264
rect 58968 15204 58972 15260
rect 58972 15204 59028 15260
rect 59028 15204 59032 15260
rect 58968 15200 59032 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 22618 14716 22682 14720
rect 22618 14660 22622 14716
rect 22622 14660 22678 14716
rect 22678 14660 22682 14716
rect 22618 14656 22682 14660
rect 22698 14716 22762 14720
rect 22698 14660 22702 14716
rect 22702 14660 22758 14716
rect 22758 14660 22762 14716
rect 22698 14656 22762 14660
rect 22778 14716 22842 14720
rect 22778 14660 22782 14716
rect 22782 14660 22838 14716
rect 22838 14660 22842 14716
rect 22778 14656 22842 14660
rect 22858 14716 22922 14720
rect 22858 14660 22862 14716
rect 22862 14660 22918 14716
rect 22918 14660 22922 14716
rect 22858 14656 22922 14660
rect 37062 14716 37126 14720
rect 37062 14660 37066 14716
rect 37066 14660 37122 14716
rect 37122 14660 37126 14716
rect 37062 14656 37126 14660
rect 37142 14716 37206 14720
rect 37142 14660 37146 14716
rect 37146 14660 37202 14716
rect 37202 14660 37206 14716
rect 37142 14656 37206 14660
rect 37222 14716 37286 14720
rect 37222 14660 37226 14716
rect 37226 14660 37282 14716
rect 37282 14660 37286 14716
rect 37222 14656 37286 14660
rect 37302 14716 37366 14720
rect 37302 14660 37306 14716
rect 37306 14660 37362 14716
rect 37362 14660 37366 14716
rect 37302 14656 37366 14660
rect 51506 14716 51570 14720
rect 51506 14660 51510 14716
rect 51510 14660 51566 14716
rect 51566 14660 51570 14716
rect 51506 14656 51570 14660
rect 51586 14716 51650 14720
rect 51586 14660 51590 14716
rect 51590 14660 51646 14716
rect 51646 14660 51650 14716
rect 51586 14656 51650 14660
rect 51666 14716 51730 14720
rect 51666 14660 51670 14716
rect 51670 14660 51726 14716
rect 51726 14660 51730 14716
rect 51666 14656 51730 14660
rect 51746 14716 51810 14720
rect 51746 14660 51750 14716
rect 51750 14660 51806 14716
rect 51806 14660 51810 14716
rect 51746 14656 51810 14660
rect 15396 14172 15460 14176
rect 15396 14116 15400 14172
rect 15400 14116 15456 14172
rect 15456 14116 15460 14172
rect 15396 14112 15460 14116
rect 15476 14172 15540 14176
rect 15476 14116 15480 14172
rect 15480 14116 15536 14172
rect 15536 14116 15540 14172
rect 15476 14112 15540 14116
rect 15556 14172 15620 14176
rect 15556 14116 15560 14172
rect 15560 14116 15616 14172
rect 15616 14116 15620 14172
rect 15556 14112 15620 14116
rect 15636 14172 15700 14176
rect 15636 14116 15640 14172
rect 15640 14116 15696 14172
rect 15696 14116 15700 14172
rect 15636 14112 15700 14116
rect 29840 14172 29904 14176
rect 29840 14116 29844 14172
rect 29844 14116 29900 14172
rect 29900 14116 29904 14172
rect 29840 14112 29904 14116
rect 29920 14172 29984 14176
rect 29920 14116 29924 14172
rect 29924 14116 29980 14172
rect 29980 14116 29984 14172
rect 29920 14112 29984 14116
rect 30000 14172 30064 14176
rect 30000 14116 30004 14172
rect 30004 14116 30060 14172
rect 30060 14116 30064 14172
rect 30000 14112 30064 14116
rect 30080 14172 30144 14176
rect 30080 14116 30084 14172
rect 30084 14116 30140 14172
rect 30140 14116 30144 14172
rect 30080 14112 30144 14116
rect 44284 14172 44348 14176
rect 44284 14116 44288 14172
rect 44288 14116 44344 14172
rect 44344 14116 44348 14172
rect 44284 14112 44348 14116
rect 44364 14172 44428 14176
rect 44364 14116 44368 14172
rect 44368 14116 44424 14172
rect 44424 14116 44428 14172
rect 44364 14112 44428 14116
rect 44444 14172 44508 14176
rect 44444 14116 44448 14172
rect 44448 14116 44504 14172
rect 44504 14116 44508 14172
rect 44444 14112 44508 14116
rect 44524 14172 44588 14176
rect 44524 14116 44528 14172
rect 44528 14116 44584 14172
rect 44584 14116 44588 14172
rect 44524 14112 44588 14116
rect 58728 14172 58792 14176
rect 58728 14116 58732 14172
rect 58732 14116 58788 14172
rect 58788 14116 58792 14172
rect 58728 14112 58792 14116
rect 58808 14172 58872 14176
rect 58808 14116 58812 14172
rect 58812 14116 58868 14172
rect 58868 14116 58872 14172
rect 58808 14112 58872 14116
rect 58888 14172 58952 14176
rect 58888 14116 58892 14172
rect 58892 14116 58948 14172
rect 58948 14116 58952 14172
rect 58888 14112 58952 14116
rect 58968 14172 59032 14176
rect 58968 14116 58972 14172
rect 58972 14116 59028 14172
rect 59028 14116 59032 14172
rect 58968 14112 59032 14116
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 22618 13628 22682 13632
rect 22618 13572 22622 13628
rect 22622 13572 22678 13628
rect 22678 13572 22682 13628
rect 22618 13568 22682 13572
rect 22698 13628 22762 13632
rect 22698 13572 22702 13628
rect 22702 13572 22758 13628
rect 22758 13572 22762 13628
rect 22698 13568 22762 13572
rect 22778 13628 22842 13632
rect 22778 13572 22782 13628
rect 22782 13572 22838 13628
rect 22838 13572 22842 13628
rect 22778 13568 22842 13572
rect 22858 13628 22922 13632
rect 22858 13572 22862 13628
rect 22862 13572 22918 13628
rect 22918 13572 22922 13628
rect 22858 13568 22922 13572
rect 37062 13628 37126 13632
rect 37062 13572 37066 13628
rect 37066 13572 37122 13628
rect 37122 13572 37126 13628
rect 37062 13568 37126 13572
rect 37142 13628 37206 13632
rect 37142 13572 37146 13628
rect 37146 13572 37202 13628
rect 37202 13572 37206 13628
rect 37142 13568 37206 13572
rect 37222 13628 37286 13632
rect 37222 13572 37226 13628
rect 37226 13572 37282 13628
rect 37282 13572 37286 13628
rect 37222 13568 37286 13572
rect 37302 13628 37366 13632
rect 37302 13572 37306 13628
rect 37306 13572 37362 13628
rect 37362 13572 37366 13628
rect 37302 13568 37366 13572
rect 51506 13628 51570 13632
rect 51506 13572 51510 13628
rect 51510 13572 51566 13628
rect 51566 13572 51570 13628
rect 51506 13568 51570 13572
rect 51586 13628 51650 13632
rect 51586 13572 51590 13628
rect 51590 13572 51646 13628
rect 51646 13572 51650 13628
rect 51586 13568 51650 13572
rect 51666 13628 51730 13632
rect 51666 13572 51670 13628
rect 51670 13572 51726 13628
rect 51726 13572 51730 13628
rect 51666 13568 51730 13572
rect 51746 13628 51810 13632
rect 51746 13572 51750 13628
rect 51750 13572 51806 13628
rect 51806 13572 51810 13628
rect 51746 13568 51810 13572
rect 15396 13084 15460 13088
rect 15396 13028 15400 13084
rect 15400 13028 15456 13084
rect 15456 13028 15460 13084
rect 15396 13024 15460 13028
rect 15476 13084 15540 13088
rect 15476 13028 15480 13084
rect 15480 13028 15536 13084
rect 15536 13028 15540 13084
rect 15476 13024 15540 13028
rect 15556 13084 15620 13088
rect 15556 13028 15560 13084
rect 15560 13028 15616 13084
rect 15616 13028 15620 13084
rect 15556 13024 15620 13028
rect 15636 13084 15700 13088
rect 15636 13028 15640 13084
rect 15640 13028 15696 13084
rect 15696 13028 15700 13084
rect 15636 13024 15700 13028
rect 29840 13084 29904 13088
rect 29840 13028 29844 13084
rect 29844 13028 29900 13084
rect 29900 13028 29904 13084
rect 29840 13024 29904 13028
rect 29920 13084 29984 13088
rect 29920 13028 29924 13084
rect 29924 13028 29980 13084
rect 29980 13028 29984 13084
rect 29920 13024 29984 13028
rect 30000 13084 30064 13088
rect 30000 13028 30004 13084
rect 30004 13028 30060 13084
rect 30060 13028 30064 13084
rect 30000 13024 30064 13028
rect 30080 13084 30144 13088
rect 30080 13028 30084 13084
rect 30084 13028 30140 13084
rect 30140 13028 30144 13084
rect 30080 13024 30144 13028
rect 44284 13084 44348 13088
rect 44284 13028 44288 13084
rect 44288 13028 44344 13084
rect 44344 13028 44348 13084
rect 44284 13024 44348 13028
rect 44364 13084 44428 13088
rect 44364 13028 44368 13084
rect 44368 13028 44424 13084
rect 44424 13028 44428 13084
rect 44364 13024 44428 13028
rect 44444 13084 44508 13088
rect 44444 13028 44448 13084
rect 44448 13028 44504 13084
rect 44504 13028 44508 13084
rect 44444 13024 44508 13028
rect 44524 13084 44588 13088
rect 44524 13028 44528 13084
rect 44528 13028 44584 13084
rect 44584 13028 44588 13084
rect 44524 13024 44588 13028
rect 58728 13084 58792 13088
rect 58728 13028 58732 13084
rect 58732 13028 58788 13084
rect 58788 13028 58792 13084
rect 58728 13024 58792 13028
rect 58808 13084 58872 13088
rect 58808 13028 58812 13084
rect 58812 13028 58868 13084
rect 58868 13028 58872 13084
rect 58808 13024 58872 13028
rect 58888 13084 58952 13088
rect 58888 13028 58892 13084
rect 58892 13028 58948 13084
rect 58948 13028 58952 13084
rect 58888 13024 58952 13028
rect 58968 13084 59032 13088
rect 58968 13028 58972 13084
rect 58972 13028 59028 13084
rect 59028 13028 59032 13084
rect 58968 13024 59032 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 22618 12540 22682 12544
rect 22618 12484 22622 12540
rect 22622 12484 22678 12540
rect 22678 12484 22682 12540
rect 22618 12480 22682 12484
rect 22698 12540 22762 12544
rect 22698 12484 22702 12540
rect 22702 12484 22758 12540
rect 22758 12484 22762 12540
rect 22698 12480 22762 12484
rect 22778 12540 22842 12544
rect 22778 12484 22782 12540
rect 22782 12484 22838 12540
rect 22838 12484 22842 12540
rect 22778 12480 22842 12484
rect 22858 12540 22922 12544
rect 22858 12484 22862 12540
rect 22862 12484 22918 12540
rect 22918 12484 22922 12540
rect 22858 12480 22922 12484
rect 37062 12540 37126 12544
rect 37062 12484 37066 12540
rect 37066 12484 37122 12540
rect 37122 12484 37126 12540
rect 37062 12480 37126 12484
rect 37142 12540 37206 12544
rect 37142 12484 37146 12540
rect 37146 12484 37202 12540
rect 37202 12484 37206 12540
rect 37142 12480 37206 12484
rect 37222 12540 37286 12544
rect 37222 12484 37226 12540
rect 37226 12484 37282 12540
rect 37282 12484 37286 12540
rect 37222 12480 37286 12484
rect 37302 12540 37366 12544
rect 37302 12484 37306 12540
rect 37306 12484 37362 12540
rect 37362 12484 37366 12540
rect 37302 12480 37366 12484
rect 51506 12540 51570 12544
rect 51506 12484 51510 12540
rect 51510 12484 51566 12540
rect 51566 12484 51570 12540
rect 51506 12480 51570 12484
rect 51586 12540 51650 12544
rect 51586 12484 51590 12540
rect 51590 12484 51646 12540
rect 51646 12484 51650 12540
rect 51586 12480 51650 12484
rect 51666 12540 51730 12544
rect 51666 12484 51670 12540
rect 51670 12484 51726 12540
rect 51726 12484 51730 12540
rect 51666 12480 51730 12484
rect 51746 12540 51810 12544
rect 51746 12484 51750 12540
rect 51750 12484 51806 12540
rect 51806 12484 51810 12540
rect 51746 12480 51810 12484
rect 15396 11996 15460 12000
rect 15396 11940 15400 11996
rect 15400 11940 15456 11996
rect 15456 11940 15460 11996
rect 15396 11936 15460 11940
rect 15476 11996 15540 12000
rect 15476 11940 15480 11996
rect 15480 11940 15536 11996
rect 15536 11940 15540 11996
rect 15476 11936 15540 11940
rect 15556 11996 15620 12000
rect 15556 11940 15560 11996
rect 15560 11940 15616 11996
rect 15616 11940 15620 11996
rect 15556 11936 15620 11940
rect 15636 11996 15700 12000
rect 15636 11940 15640 11996
rect 15640 11940 15696 11996
rect 15696 11940 15700 11996
rect 15636 11936 15700 11940
rect 29840 11996 29904 12000
rect 29840 11940 29844 11996
rect 29844 11940 29900 11996
rect 29900 11940 29904 11996
rect 29840 11936 29904 11940
rect 29920 11996 29984 12000
rect 29920 11940 29924 11996
rect 29924 11940 29980 11996
rect 29980 11940 29984 11996
rect 29920 11936 29984 11940
rect 30000 11996 30064 12000
rect 30000 11940 30004 11996
rect 30004 11940 30060 11996
rect 30060 11940 30064 11996
rect 30000 11936 30064 11940
rect 30080 11996 30144 12000
rect 30080 11940 30084 11996
rect 30084 11940 30140 11996
rect 30140 11940 30144 11996
rect 30080 11936 30144 11940
rect 44284 11996 44348 12000
rect 44284 11940 44288 11996
rect 44288 11940 44344 11996
rect 44344 11940 44348 11996
rect 44284 11936 44348 11940
rect 44364 11996 44428 12000
rect 44364 11940 44368 11996
rect 44368 11940 44424 11996
rect 44424 11940 44428 11996
rect 44364 11936 44428 11940
rect 44444 11996 44508 12000
rect 44444 11940 44448 11996
rect 44448 11940 44504 11996
rect 44504 11940 44508 11996
rect 44444 11936 44508 11940
rect 44524 11996 44588 12000
rect 44524 11940 44528 11996
rect 44528 11940 44584 11996
rect 44584 11940 44588 11996
rect 44524 11936 44588 11940
rect 58728 11996 58792 12000
rect 58728 11940 58732 11996
rect 58732 11940 58788 11996
rect 58788 11940 58792 11996
rect 58728 11936 58792 11940
rect 58808 11996 58872 12000
rect 58808 11940 58812 11996
rect 58812 11940 58868 11996
rect 58868 11940 58872 11996
rect 58808 11936 58872 11940
rect 58888 11996 58952 12000
rect 58888 11940 58892 11996
rect 58892 11940 58948 11996
rect 58948 11940 58952 11996
rect 58888 11936 58952 11940
rect 58968 11996 59032 12000
rect 58968 11940 58972 11996
rect 58972 11940 59028 11996
rect 59028 11940 59032 11996
rect 58968 11936 59032 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 22618 11452 22682 11456
rect 22618 11396 22622 11452
rect 22622 11396 22678 11452
rect 22678 11396 22682 11452
rect 22618 11392 22682 11396
rect 22698 11452 22762 11456
rect 22698 11396 22702 11452
rect 22702 11396 22758 11452
rect 22758 11396 22762 11452
rect 22698 11392 22762 11396
rect 22778 11452 22842 11456
rect 22778 11396 22782 11452
rect 22782 11396 22838 11452
rect 22838 11396 22842 11452
rect 22778 11392 22842 11396
rect 22858 11452 22922 11456
rect 22858 11396 22862 11452
rect 22862 11396 22918 11452
rect 22918 11396 22922 11452
rect 22858 11392 22922 11396
rect 37062 11452 37126 11456
rect 37062 11396 37066 11452
rect 37066 11396 37122 11452
rect 37122 11396 37126 11452
rect 37062 11392 37126 11396
rect 37142 11452 37206 11456
rect 37142 11396 37146 11452
rect 37146 11396 37202 11452
rect 37202 11396 37206 11452
rect 37142 11392 37206 11396
rect 37222 11452 37286 11456
rect 37222 11396 37226 11452
rect 37226 11396 37282 11452
rect 37282 11396 37286 11452
rect 37222 11392 37286 11396
rect 37302 11452 37366 11456
rect 37302 11396 37306 11452
rect 37306 11396 37362 11452
rect 37362 11396 37366 11452
rect 37302 11392 37366 11396
rect 51506 11452 51570 11456
rect 51506 11396 51510 11452
rect 51510 11396 51566 11452
rect 51566 11396 51570 11452
rect 51506 11392 51570 11396
rect 51586 11452 51650 11456
rect 51586 11396 51590 11452
rect 51590 11396 51646 11452
rect 51646 11396 51650 11452
rect 51586 11392 51650 11396
rect 51666 11452 51730 11456
rect 51666 11396 51670 11452
rect 51670 11396 51726 11452
rect 51726 11396 51730 11452
rect 51666 11392 51730 11396
rect 51746 11452 51810 11456
rect 51746 11396 51750 11452
rect 51750 11396 51806 11452
rect 51806 11396 51810 11452
rect 51746 11392 51810 11396
rect 15396 10908 15460 10912
rect 15396 10852 15400 10908
rect 15400 10852 15456 10908
rect 15456 10852 15460 10908
rect 15396 10848 15460 10852
rect 15476 10908 15540 10912
rect 15476 10852 15480 10908
rect 15480 10852 15536 10908
rect 15536 10852 15540 10908
rect 15476 10848 15540 10852
rect 15556 10908 15620 10912
rect 15556 10852 15560 10908
rect 15560 10852 15616 10908
rect 15616 10852 15620 10908
rect 15556 10848 15620 10852
rect 15636 10908 15700 10912
rect 15636 10852 15640 10908
rect 15640 10852 15696 10908
rect 15696 10852 15700 10908
rect 15636 10848 15700 10852
rect 29840 10908 29904 10912
rect 29840 10852 29844 10908
rect 29844 10852 29900 10908
rect 29900 10852 29904 10908
rect 29840 10848 29904 10852
rect 29920 10908 29984 10912
rect 29920 10852 29924 10908
rect 29924 10852 29980 10908
rect 29980 10852 29984 10908
rect 29920 10848 29984 10852
rect 30000 10908 30064 10912
rect 30000 10852 30004 10908
rect 30004 10852 30060 10908
rect 30060 10852 30064 10908
rect 30000 10848 30064 10852
rect 30080 10908 30144 10912
rect 30080 10852 30084 10908
rect 30084 10852 30140 10908
rect 30140 10852 30144 10908
rect 30080 10848 30144 10852
rect 44284 10908 44348 10912
rect 44284 10852 44288 10908
rect 44288 10852 44344 10908
rect 44344 10852 44348 10908
rect 44284 10848 44348 10852
rect 44364 10908 44428 10912
rect 44364 10852 44368 10908
rect 44368 10852 44424 10908
rect 44424 10852 44428 10908
rect 44364 10848 44428 10852
rect 44444 10908 44508 10912
rect 44444 10852 44448 10908
rect 44448 10852 44504 10908
rect 44504 10852 44508 10908
rect 44444 10848 44508 10852
rect 44524 10908 44588 10912
rect 44524 10852 44528 10908
rect 44528 10852 44584 10908
rect 44584 10852 44588 10908
rect 44524 10848 44588 10852
rect 58728 10908 58792 10912
rect 58728 10852 58732 10908
rect 58732 10852 58788 10908
rect 58788 10852 58792 10908
rect 58728 10848 58792 10852
rect 58808 10908 58872 10912
rect 58808 10852 58812 10908
rect 58812 10852 58868 10908
rect 58868 10852 58872 10908
rect 58808 10848 58872 10852
rect 58888 10908 58952 10912
rect 58888 10852 58892 10908
rect 58892 10852 58948 10908
rect 58948 10852 58952 10908
rect 58888 10848 58952 10852
rect 58968 10908 59032 10912
rect 58968 10852 58972 10908
rect 58972 10852 59028 10908
rect 59028 10852 59032 10908
rect 58968 10848 59032 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 22618 10364 22682 10368
rect 22618 10308 22622 10364
rect 22622 10308 22678 10364
rect 22678 10308 22682 10364
rect 22618 10304 22682 10308
rect 22698 10364 22762 10368
rect 22698 10308 22702 10364
rect 22702 10308 22758 10364
rect 22758 10308 22762 10364
rect 22698 10304 22762 10308
rect 22778 10364 22842 10368
rect 22778 10308 22782 10364
rect 22782 10308 22838 10364
rect 22838 10308 22842 10364
rect 22778 10304 22842 10308
rect 22858 10364 22922 10368
rect 22858 10308 22862 10364
rect 22862 10308 22918 10364
rect 22918 10308 22922 10364
rect 22858 10304 22922 10308
rect 37062 10364 37126 10368
rect 37062 10308 37066 10364
rect 37066 10308 37122 10364
rect 37122 10308 37126 10364
rect 37062 10304 37126 10308
rect 37142 10364 37206 10368
rect 37142 10308 37146 10364
rect 37146 10308 37202 10364
rect 37202 10308 37206 10364
rect 37142 10304 37206 10308
rect 37222 10364 37286 10368
rect 37222 10308 37226 10364
rect 37226 10308 37282 10364
rect 37282 10308 37286 10364
rect 37222 10304 37286 10308
rect 37302 10364 37366 10368
rect 37302 10308 37306 10364
rect 37306 10308 37362 10364
rect 37362 10308 37366 10364
rect 37302 10304 37366 10308
rect 51506 10364 51570 10368
rect 51506 10308 51510 10364
rect 51510 10308 51566 10364
rect 51566 10308 51570 10364
rect 51506 10304 51570 10308
rect 51586 10364 51650 10368
rect 51586 10308 51590 10364
rect 51590 10308 51646 10364
rect 51646 10308 51650 10364
rect 51586 10304 51650 10308
rect 51666 10364 51730 10368
rect 51666 10308 51670 10364
rect 51670 10308 51726 10364
rect 51726 10308 51730 10364
rect 51666 10304 51730 10308
rect 51746 10364 51810 10368
rect 51746 10308 51750 10364
rect 51750 10308 51806 10364
rect 51806 10308 51810 10364
rect 51746 10304 51810 10308
rect 15396 9820 15460 9824
rect 15396 9764 15400 9820
rect 15400 9764 15456 9820
rect 15456 9764 15460 9820
rect 15396 9760 15460 9764
rect 15476 9820 15540 9824
rect 15476 9764 15480 9820
rect 15480 9764 15536 9820
rect 15536 9764 15540 9820
rect 15476 9760 15540 9764
rect 15556 9820 15620 9824
rect 15556 9764 15560 9820
rect 15560 9764 15616 9820
rect 15616 9764 15620 9820
rect 15556 9760 15620 9764
rect 15636 9820 15700 9824
rect 15636 9764 15640 9820
rect 15640 9764 15696 9820
rect 15696 9764 15700 9820
rect 15636 9760 15700 9764
rect 29840 9820 29904 9824
rect 29840 9764 29844 9820
rect 29844 9764 29900 9820
rect 29900 9764 29904 9820
rect 29840 9760 29904 9764
rect 29920 9820 29984 9824
rect 29920 9764 29924 9820
rect 29924 9764 29980 9820
rect 29980 9764 29984 9820
rect 29920 9760 29984 9764
rect 30000 9820 30064 9824
rect 30000 9764 30004 9820
rect 30004 9764 30060 9820
rect 30060 9764 30064 9820
rect 30000 9760 30064 9764
rect 30080 9820 30144 9824
rect 30080 9764 30084 9820
rect 30084 9764 30140 9820
rect 30140 9764 30144 9820
rect 30080 9760 30144 9764
rect 44284 9820 44348 9824
rect 44284 9764 44288 9820
rect 44288 9764 44344 9820
rect 44344 9764 44348 9820
rect 44284 9760 44348 9764
rect 44364 9820 44428 9824
rect 44364 9764 44368 9820
rect 44368 9764 44424 9820
rect 44424 9764 44428 9820
rect 44364 9760 44428 9764
rect 44444 9820 44508 9824
rect 44444 9764 44448 9820
rect 44448 9764 44504 9820
rect 44504 9764 44508 9820
rect 44444 9760 44508 9764
rect 44524 9820 44588 9824
rect 44524 9764 44528 9820
rect 44528 9764 44584 9820
rect 44584 9764 44588 9820
rect 44524 9760 44588 9764
rect 58728 9820 58792 9824
rect 58728 9764 58732 9820
rect 58732 9764 58788 9820
rect 58788 9764 58792 9820
rect 58728 9760 58792 9764
rect 58808 9820 58872 9824
rect 58808 9764 58812 9820
rect 58812 9764 58868 9820
rect 58868 9764 58872 9820
rect 58808 9760 58872 9764
rect 58888 9820 58952 9824
rect 58888 9764 58892 9820
rect 58892 9764 58948 9820
rect 58948 9764 58952 9820
rect 58888 9760 58952 9764
rect 58968 9820 59032 9824
rect 58968 9764 58972 9820
rect 58972 9764 59028 9820
rect 59028 9764 59032 9820
rect 58968 9760 59032 9764
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 22618 9276 22682 9280
rect 22618 9220 22622 9276
rect 22622 9220 22678 9276
rect 22678 9220 22682 9276
rect 22618 9216 22682 9220
rect 22698 9276 22762 9280
rect 22698 9220 22702 9276
rect 22702 9220 22758 9276
rect 22758 9220 22762 9276
rect 22698 9216 22762 9220
rect 22778 9276 22842 9280
rect 22778 9220 22782 9276
rect 22782 9220 22838 9276
rect 22838 9220 22842 9276
rect 22778 9216 22842 9220
rect 22858 9276 22922 9280
rect 22858 9220 22862 9276
rect 22862 9220 22918 9276
rect 22918 9220 22922 9276
rect 22858 9216 22922 9220
rect 37062 9276 37126 9280
rect 37062 9220 37066 9276
rect 37066 9220 37122 9276
rect 37122 9220 37126 9276
rect 37062 9216 37126 9220
rect 37142 9276 37206 9280
rect 37142 9220 37146 9276
rect 37146 9220 37202 9276
rect 37202 9220 37206 9276
rect 37142 9216 37206 9220
rect 37222 9276 37286 9280
rect 37222 9220 37226 9276
rect 37226 9220 37282 9276
rect 37282 9220 37286 9276
rect 37222 9216 37286 9220
rect 37302 9276 37366 9280
rect 37302 9220 37306 9276
rect 37306 9220 37362 9276
rect 37362 9220 37366 9276
rect 37302 9216 37366 9220
rect 51506 9276 51570 9280
rect 51506 9220 51510 9276
rect 51510 9220 51566 9276
rect 51566 9220 51570 9276
rect 51506 9216 51570 9220
rect 51586 9276 51650 9280
rect 51586 9220 51590 9276
rect 51590 9220 51646 9276
rect 51646 9220 51650 9276
rect 51586 9216 51650 9220
rect 51666 9276 51730 9280
rect 51666 9220 51670 9276
rect 51670 9220 51726 9276
rect 51726 9220 51730 9276
rect 51666 9216 51730 9220
rect 51746 9276 51810 9280
rect 51746 9220 51750 9276
rect 51750 9220 51806 9276
rect 51806 9220 51810 9276
rect 51746 9216 51810 9220
rect 15396 8732 15460 8736
rect 15396 8676 15400 8732
rect 15400 8676 15456 8732
rect 15456 8676 15460 8732
rect 15396 8672 15460 8676
rect 15476 8732 15540 8736
rect 15476 8676 15480 8732
rect 15480 8676 15536 8732
rect 15536 8676 15540 8732
rect 15476 8672 15540 8676
rect 15556 8732 15620 8736
rect 15556 8676 15560 8732
rect 15560 8676 15616 8732
rect 15616 8676 15620 8732
rect 15556 8672 15620 8676
rect 15636 8732 15700 8736
rect 15636 8676 15640 8732
rect 15640 8676 15696 8732
rect 15696 8676 15700 8732
rect 15636 8672 15700 8676
rect 29840 8732 29904 8736
rect 29840 8676 29844 8732
rect 29844 8676 29900 8732
rect 29900 8676 29904 8732
rect 29840 8672 29904 8676
rect 29920 8732 29984 8736
rect 29920 8676 29924 8732
rect 29924 8676 29980 8732
rect 29980 8676 29984 8732
rect 29920 8672 29984 8676
rect 30000 8732 30064 8736
rect 30000 8676 30004 8732
rect 30004 8676 30060 8732
rect 30060 8676 30064 8732
rect 30000 8672 30064 8676
rect 30080 8732 30144 8736
rect 30080 8676 30084 8732
rect 30084 8676 30140 8732
rect 30140 8676 30144 8732
rect 30080 8672 30144 8676
rect 44284 8732 44348 8736
rect 44284 8676 44288 8732
rect 44288 8676 44344 8732
rect 44344 8676 44348 8732
rect 44284 8672 44348 8676
rect 44364 8732 44428 8736
rect 44364 8676 44368 8732
rect 44368 8676 44424 8732
rect 44424 8676 44428 8732
rect 44364 8672 44428 8676
rect 44444 8732 44508 8736
rect 44444 8676 44448 8732
rect 44448 8676 44504 8732
rect 44504 8676 44508 8732
rect 44444 8672 44508 8676
rect 44524 8732 44588 8736
rect 44524 8676 44528 8732
rect 44528 8676 44584 8732
rect 44584 8676 44588 8732
rect 44524 8672 44588 8676
rect 58728 8732 58792 8736
rect 58728 8676 58732 8732
rect 58732 8676 58788 8732
rect 58788 8676 58792 8732
rect 58728 8672 58792 8676
rect 58808 8732 58872 8736
rect 58808 8676 58812 8732
rect 58812 8676 58868 8732
rect 58868 8676 58872 8732
rect 58808 8672 58872 8676
rect 58888 8732 58952 8736
rect 58888 8676 58892 8732
rect 58892 8676 58948 8732
rect 58948 8676 58952 8732
rect 58888 8672 58952 8676
rect 58968 8732 59032 8736
rect 58968 8676 58972 8732
rect 58972 8676 59028 8732
rect 59028 8676 59032 8732
rect 58968 8672 59032 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 22618 8188 22682 8192
rect 22618 8132 22622 8188
rect 22622 8132 22678 8188
rect 22678 8132 22682 8188
rect 22618 8128 22682 8132
rect 22698 8188 22762 8192
rect 22698 8132 22702 8188
rect 22702 8132 22758 8188
rect 22758 8132 22762 8188
rect 22698 8128 22762 8132
rect 22778 8188 22842 8192
rect 22778 8132 22782 8188
rect 22782 8132 22838 8188
rect 22838 8132 22842 8188
rect 22778 8128 22842 8132
rect 22858 8188 22922 8192
rect 22858 8132 22862 8188
rect 22862 8132 22918 8188
rect 22918 8132 22922 8188
rect 22858 8128 22922 8132
rect 37062 8188 37126 8192
rect 37062 8132 37066 8188
rect 37066 8132 37122 8188
rect 37122 8132 37126 8188
rect 37062 8128 37126 8132
rect 37142 8188 37206 8192
rect 37142 8132 37146 8188
rect 37146 8132 37202 8188
rect 37202 8132 37206 8188
rect 37142 8128 37206 8132
rect 37222 8188 37286 8192
rect 37222 8132 37226 8188
rect 37226 8132 37282 8188
rect 37282 8132 37286 8188
rect 37222 8128 37286 8132
rect 37302 8188 37366 8192
rect 37302 8132 37306 8188
rect 37306 8132 37362 8188
rect 37362 8132 37366 8188
rect 37302 8128 37366 8132
rect 51506 8188 51570 8192
rect 51506 8132 51510 8188
rect 51510 8132 51566 8188
rect 51566 8132 51570 8188
rect 51506 8128 51570 8132
rect 51586 8188 51650 8192
rect 51586 8132 51590 8188
rect 51590 8132 51646 8188
rect 51646 8132 51650 8188
rect 51586 8128 51650 8132
rect 51666 8188 51730 8192
rect 51666 8132 51670 8188
rect 51670 8132 51726 8188
rect 51726 8132 51730 8188
rect 51666 8128 51730 8132
rect 51746 8188 51810 8192
rect 51746 8132 51750 8188
rect 51750 8132 51806 8188
rect 51806 8132 51810 8188
rect 51746 8128 51810 8132
rect 15396 7644 15460 7648
rect 15396 7588 15400 7644
rect 15400 7588 15456 7644
rect 15456 7588 15460 7644
rect 15396 7584 15460 7588
rect 15476 7644 15540 7648
rect 15476 7588 15480 7644
rect 15480 7588 15536 7644
rect 15536 7588 15540 7644
rect 15476 7584 15540 7588
rect 15556 7644 15620 7648
rect 15556 7588 15560 7644
rect 15560 7588 15616 7644
rect 15616 7588 15620 7644
rect 15556 7584 15620 7588
rect 15636 7644 15700 7648
rect 15636 7588 15640 7644
rect 15640 7588 15696 7644
rect 15696 7588 15700 7644
rect 15636 7584 15700 7588
rect 29840 7644 29904 7648
rect 29840 7588 29844 7644
rect 29844 7588 29900 7644
rect 29900 7588 29904 7644
rect 29840 7584 29904 7588
rect 29920 7644 29984 7648
rect 29920 7588 29924 7644
rect 29924 7588 29980 7644
rect 29980 7588 29984 7644
rect 29920 7584 29984 7588
rect 30000 7644 30064 7648
rect 30000 7588 30004 7644
rect 30004 7588 30060 7644
rect 30060 7588 30064 7644
rect 30000 7584 30064 7588
rect 30080 7644 30144 7648
rect 30080 7588 30084 7644
rect 30084 7588 30140 7644
rect 30140 7588 30144 7644
rect 30080 7584 30144 7588
rect 44284 7644 44348 7648
rect 44284 7588 44288 7644
rect 44288 7588 44344 7644
rect 44344 7588 44348 7644
rect 44284 7584 44348 7588
rect 44364 7644 44428 7648
rect 44364 7588 44368 7644
rect 44368 7588 44424 7644
rect 44424 7588 44428 7644
rect 44364 7584 44428 7588
rect 44444 7644 44508 7648
rect 44444 7588 44448 7644
rect 44448 7588 44504 7644
rect 44504 7588 44508 7644
rect 44444 7584 44508 7588
rect 44524 7644 44588 7648
rect 44524 7588 44528 7644
rect 44528 7588 44584 7644
rect 44584 7588 44588 7644
rect 44524 7584 44588 7588
rect 58728 7644 58792 7648
rect 58728 7588 58732 7644
rect 58732 7588 58788 7644
rect 58788 7588 58792 7644
rect 58728 7584 58792 7588
rect 58808 7644 58872 7648
rect 58808 7588 58812 7644
rect 58812 7588 58868 7644
rect 58868 7588 58872 7644
rect 58808 7584 58872 7588
rect 58888 7644 58952 7648
rect 58888 7588 58892 7644
rect 58892 7588 58948 7644
rect 58948 7588 58952 7644
rect 58888 7584 58952 7588
rect 58968 7644 59032 7648
rect 58968 7588 58972 7644
rect 58972 7588 59028 7644
rect 59028 7588 59032 7644
rect 58968 7584 59032 7588
rect 7236 7244 7300 7308
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 22618 7100 22682 7104
rect 22618 7044 22622 7100
rect 22622 7044 22678 7100
rect 22678 7044 22682 7100
rect 22618 7040 22682 7044
rect 22698 7100 22762 7104
rect 22698 7044 22702 7100
rect 22702 7044 22758 7100
rect 22758 7044 22762 7100
rect 22698 7040 22762 7044
rect 22778 7100 22842 7104
rect 22778 7044 22782 7100
rect 22782 7044 22838 7100
rect 22838 7044 22842 7100
rect 22778 7040 22842 7044
rect 22858 7100 22922 7104
rect 22858 7044 22862 7100
rect 22862 7044 22918 7100
rect 22918 7044 22922 7100
rect 22858 7040 22922 7044
rect 37062 7100 37126 7104
rect 37062 7044 37066 7100
rect 37066 7044 37122 7100
rect 37122 7044 37126 7100
rect 37062 7040 37126 7044
rect 37142 7100 37206 7104
rect 37142 7044 37146 7100
rect 37146 7044 37202 7100
rect 37202 7044 37206 7100
rect 37142 7040 37206 7044
rect 37222 7100 37286 7104
rect 37222 7044 37226 7100
rect 37226 7044 37282 7100
rect 37282 7044 37286 7100
rect 37222 7040 37286 7044
rect 37302 7100 37366 7104
rect 37302 7044 37306 7100
rect 37306 7044 37362 7100
rect 37362 7044 37366 7100
rect 37302 7040 37366 7044
rect 51506 7100 51570 7104
rect 51506 7044 51510 7100
rect 51510 7044 51566 7100
rect 51566 7044 51570 7100
rect 51506 7040 51570 7044
rect 51586 7100 51650 7104
rect 51586 7044 51590 7100
rect 51590 7044 51646 7100
rect 51646 7044 51650 7100
rect 51586 7040 51650 7044
rect 51666 7100 51730 7104
rect 51666 7044 51670 7100
rect 51670 7044 51726 7100
rect 51726 7044 51730 7100
rect 51666 7040 51730 7044
rect 51746 7100 51810 7104
rect 51746 7044 51750 7100
rect 51750 7044 51806 7100
rect 51806 7044 51810 7100
rect 51746 7040 51810 7044
rect 55996 6972 56060 7036
rect 15396 6556 15460 6560
rect 15396 6500 15400 6556
rect 15400 6500 15456 6556
rect 15456 6500 15460 6556
rect 15396 6496 15460 6500
rect 15476 6556 15540 6560
rect 15476 6500 15480 6556
rect 15480 6500 15536 6556
rect 15536 6500 15540 6556
rect 15476 6496 15540 6500
rect 15556 6556 15620 6560
rect 15556 6500 15560 6556
rect 15560 6500 15616 6556
rect 15616 6500 15620 6556
rect 15556 6496 15620 6500
rect 15636 6556 15700 6560
rect 15636 6500 15640 6556
rect 15640 6500 15696 6556
rect 15696 6500 15700 6556
rect 15636 6496 15700 6500
rect 29840 6556 29904 6560
rect 29840 6500 29844 6556
rect 29844 6500 29900 6556
rect 29900 6500 29904 6556
rect 29840 6496 29904 6500
rect 29920 6556 29984 6560
rect 29920 6500 29924 6556
rect 29924 6500 29980 6556
rect 29980 6500 29984 6556
rect 29920 6496 29984 6500
rect 30000 6556 30064 6560
rect 30000 6500 30004 6556
rect 30004 6500 30060 6556
rect 30060 6500 30064 6556
rect 30000 6496 30064 6500
rect 30080 6556 30144 6560
rect 30080 6500 30084 6556
rect 30084 6500 30140 6556
rect 30140 6500 30144 6556
rect 30080 6496 30144 6500
rect 44284 6556 44348 6560
rect 44284 6500 44288 6556
rect 44288 6500 44344 6556
rect 44344 6500 44348 6556
rect 44284 6496 44348 6500
rect 44364 6556 44428 6560
rect 44364 6500 44368 6556
rect 44368 6500 44424 6556
rect 44424 6500 44428 6556
rect 44364 6496 44428 6500
rect 44444 6556 44508 6560
rect 44444 6500 44448 6556
rect 44448 6500 44504 6556
rect 44504 6500 44508 6556
rect 44444 6496 44508 6500
rect 44524 6556 44588 6560
rect 44524 6500 44528 6556
rect 44528 6500 44584 6556
rect 44584 6500 44588 6556
rect 44524 6496 44588 6500
rect 58728 6556 58792 6560
rect 58728 6500 58732 6556
rect 58732 6500 58788 6556
rect 58788 6500 58792 6556
rect 58728 6496 58792 6500
rect 58808 6556 58872 6560
rect 58808 6500 58812 6556
rect 58812 6500 58868 6556
rect 58868 6500 58872 6556
rect 58808 6496 58872 6500
rect 58888 6556 58952 6560
rect 58888 6500 58892 6556
rect 58892 6500 58948 6556
rect 58948 6500 58952 6556
rect 58888 6496 58952 6500
rect 58968 6556 59032 6560
rect 58968 6500 58972 6556
rect 58972 6500 59028 6556
rect 59028 6500 59032 6556
rect 58968 6496 59032 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 22618 6012 22682 6016
rect 22618 5956 22622 6012
rect 22622 5956 22678 6012
rect 22678 5956 22682 6012
rect 22618 5952 22682 5956
rect 22698 6012 22762 6016
rect 22698 5956 22702 6012
rect 22702 5956 22758 6012
rect 22758 5956 22762 6012
rect 22698 5952 22762 5956
rect 22778 6012 22842 6016
rect 22778 5956 22782 6012
rect 22782 5956 22838 6012
rect 22838 5956 22842 6012
rect 22778 5952 22842 5956
rect 22858 6012 22922 6016
rect 22858 5956 22862 6012
rect 22862 5956 22918 6012
rect 22918 5956 22922 6012
rect 22858 5952 22922 5956
rect 37062 6012 37126 6016
rect 37062 5956 37066 6012
rect 37066 5956 37122 6012
rect 37122 5956 37126 6012
rect 37062 5952 37126 5956
rect 37142 6012 37206 6016
rect 37142 5956 37146 6012
rect 37146 5956 37202 6012
rect 37202 5956 37206 6012
rect 37142 5952 37206 5956
rect 37222 6012 37286 6016
rect 37222 5956 37226 6012
rect 37226 5956 37282 6012
rect 37282 5956 37286 6012
rect 37222 5952 37286 5956
rect 37302 6012 37366 6016
rect 37302 5956 37306 6012
rect 37306 5956 37362 6012
rect 37362 5956 37366 6012
rect 37302 5952 37366 5956
rect 51506 6012 51570 6016
rect 51506 5956 51510 6012
rect 51510 5956 51566 6012
rect 51566 5956 51570 6012
rect 51506 5952 51570 5956
rect 51586 6012 51650 6016
rect 51586 5956 51590 6012
rect 51590 5956 51646 6012
rect 51646 5956 51650 6012
rect 51586 5952 51650 5956
rect 51666 6012 51730 6016
rect 51666 5956 51670 6012
rect 51670 5956 51726 6012
rect 51726 5956 51730 6012
rect 51666 5952 51730 5956
rect 51746 6012 51810 6016
rect 51746 5956 51750 6012
rect 51750 5956 51806 6012
rect 51806 5956 51810 6012
rect 51746 5952 51810 5956
rect 7236 5476 7300 5540
rect 15396 5468 15460 5472
rect 15396 5412 15400 5468
rect 15400 5412 15456 5468
rect 15456 5412 15460 5468
rect 15396 5408 15460 5412
rect 15476 5468 15540 5472
rect 15476 5412 15480 5468
rect 15480 5412 15536 5468
rect 15536 5412 15540 5468
rect 15476 5408 15540 5412
rect 15556 5468 15620 5472
rect 15556 5412 15560 5468
rect 15560 5412 15616 5468
rect 15616 5412 15620 5468
rect 15556 5408 15620 5412
rect 15636 5468 15700 5472
rect 15636 5412 15640 5468
rect 15640 5412 15696 5468
rect 15696 5412 15700 5468
rect 15636 5408 15700 5412
rect 29840 5468 29904 5472
rect 29840 5412 29844 5468
rect 29844 5412 29900 5468
rect 29900 5412 29904 5468
rect 29840 5408 29904 5412
rect 29920 5468 29984 5472
rect 29920 5412 29924 5468
rect 29924 5412 29980 5468
rect 29980 5412 29984 5468
rect 29920 5408 29984 5412
rect 30000 5468 30064 5472
rect 30000 5412 30004 5468
rect 30004 5412 30060 5468
rect 30060 5412 30064 5468
rect 30000 5408 30064 5412
rect 30080 5468 30144 5472
rect 30080 5412 30084 5468
rect 30084 5412 30140 5468
rect 30140 5412 30144 5468
rect 30080 5408 30144 5412
rect 44284 5468 44348 5472
rect 44284 5412 44288 5468
rect 44288 5412 44344 5468
rect 44344 5412 44348 5468
rect 44284 5408 44348 5412
rect 44364 5468 44428 5472
rect 44364 5412 44368 5468
rect 44368 5412 44424 5468
rect 44424 5412 44428 5468
rect 44364 5408 44428 5412
rect 44444 5468 44508 5472
rect 44444 5412 44448 5468
rect 44448 5412 44504 5468
rect 44504 5412 44508 5468
rect 44444 5408 44508 5412
rect 44524 5468 44588 5472
rect 44524 5412 44528 5468
rect 44528 5412 44584 5468
rect 44584 5412 44588 5468
rect 44524 5408 44588 5412
rect 58728 5468 58792 5472
rect 58728 5412 58732 5468
rect 58732 5412 58788 5468
rect 58788 5412 58792 5468
rect 58728 5408 58792 5412
rect 58808 5468 58872 5472
rect 58808 5412 58812 5468
rect 58812 5412 58868 5468
rect 58868 5412 58872 5468
rect 58808 5408 58872 5412
rect 58888 5468 58952 5472
rect 58888 5412 58892 5468
rect 58892 5412 58948 5468
rect 58948 5412 58952 5468
rect 58888 5408 58952 5412
rect 58968 5468 59032 5472
rect 58968 5412 58972 5468
rect 58972 5412 59028 5468
rect 59028 5412 59032 5468
rect 58968 5408 59032 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 22618 4924 22682 4928
rect 22618 4868 22622 4924
rect 22622 4868 22678 4924
rect 22678 4868 22682 4924
rect 22618 4864 22682 4868
rect 22698 4924 22762 4928
rect 22698 4868 22702 4924
rect 22702 4868 22758 4924
rect 22758 4868 22762 4924
rect 22698 4864 22762 4868
rect 22778 4924 22842 4928
rect 22778 4868 22782 4924
rect 22782 4868 22838 4924
rect 22838 4868 22842 4924
rect 22778 4864 22842 4868
rect 22858 4924 22922 4928
rect 22858 4868 22862 4924
rect 22862 4868 22918 4924
rect 22918 4868 22922 4924
rect 22858 4864 22922 4868
rect 37062 4924 37126 4928
rect 37062 4868 37066 4924
rect 37066 4868 37122 4924
rect 37122 4868 37126 4924
rect 37062 4864 37126 4868
rect 37142 4924 37206 4928
rect 37142 4868 37146 4924
rect 37146 4868 37202 4924
rect 37202 4868 37206 4924
rect 37142 4864 37206 4868
rect 37222 4924 37286 4928
rect 37222 4868 37226 4924
rect 37226 4868 37282 4924
rect 37282 4868 37286 4924
rect 37222 4864 37286 4868
rect 37302 4924 37366 4928
rect 37302 4868 37306 4924
rect 37306 4868 37362 4924
rect 37362 4868 37366 4924
rect 37302 4864 37366 4868
rect 51506 4924 51570 4928
rect 51506 4868 51510 4924
rect 51510 4868 51566 4924
rect 51566 4868 51570 4924
rect 51506 4864 51570 4868
rect 51586 4924 51650 4928
rect 51586 4868 51590 4924
rect 51590 4868 51646 4924
rect 51646 4868 51650 4924
rect 51586 4864 51650 4868
rect 51666 4924 51730 4928
rect 51666 4868 51670 4924
rect 51670 4868 51726 4924
rect 51726 4868 51730 4924
rect 51666 4864 51730 4868
rect 51746 4924 51810 4928
rect 51746 4868 51750 4924
rect 51750 4868 51806 4924
rect 51806 4868 51810 4924
rect 51746 4864 51810 4868
rect 15396 4380 15460 4384
rect 15396 4324 15400 4380
rect 15400 4324 15456 4380
rect 15456 4324 15460 4380
rect 15396 4320 15460 4324
rect 15476 4380 15540 4384
rect 15476 4324 15480 4380
rect 15480 4324 15536 4380
rect 15536 4324 15540 4380
rect 15476 4320 15540 4324
rect 15556 4380 15620 4384
rect 15556 4324 15560 4380
rect 15560 4324 15616 4380
rect 15616 4324 15620 4380
rect 15556 4320 15620 4324
rect 15636 4380 15700 4384
rect 15636 4324 15640 4380
rect 15640 4324 15696 4380
rect 15696 4324 15700 4380
rect 15636 4320 15700 4324
rect 29840 4380 29904 4384
rect 29840 4324 29844 4380
rect 29844 4324 29900 4380
rect 29900 4324 29904 4380
rect 29840 4320 29904 4324
rect 29920 4380 29984 4384
rect 29920 4324 29924 4380
rect 29924 4324 29980 4380
rect 29980 4324 29984 4380
rect 29920 4320 29984 4324
rect 30000 4380 30064 4384
rect 30000 4324 30004 4380
rect 30004 4324 30060 4380
rect 30060 4324 30064 4380
rect 30000 4320 30064 4324
rect 30080 4380 30144 4384
rect 30080 4324 30084 4380
rect 30084 4324 30140 4380
rect 30140 4324 30144 4380
rect 30080 4320 30144 4324
rect 44284 4380 44348 4384
rect 44284 4324 44288 4380
rect 44288 4324 44344 4380
rect 44344 4324 44348 4380
rect 44284 4320 44348 4324
rect 44364 4380 44428 4384
rect 44364 4324 44368 4380
rect 44368 4324 44424 4380
rect 44424 4324 44428 4380
rect 44364 4320 44428 4324
rect 44444 4380 44508 4384
rect 44444 4324 44448 4380
rect 44448 4324 44504 4380
rect 44504 4324 44508 4380
rect 44444 4320 44508 4324
rect 44524 4380 44588 4384
rect 44524 4324 44528 4380
rect 44528 4324 44584 4380
rect 44584 4324 44588 4380
rect 44524 4320 44588 4324
rect 58728 4380 58792 4384
rect 58728 4324 58732 4380
rect 58732 4324 58788 4380
rect 58788 4324 58792 4380
rect 58728 4320 58792 4324
rect 58808 4380 58872 4384
rect 58808 4324 58812 4380
rect 58812 4324 58868 4380
rect 58868 4324 58872 4380
rect 58808 4320 58872 4324
rect 58888 4380 58952 4384
rect 58888 4324 58892 4380
rect 58892 4324 58948 4380
rect 58948 4324 58952 4380
rect 58888 4320 58952 4324
rect 58968 4380 59032 4384
rect 58968 4324 58972 4380
rect 58972 4324 59028 4380
rect 59028 4324 59032 4380
rect 58968 4320 59032 4324
rect 55996 3980 56060 4044
rect 35572 3844 35636 3908
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 22618 3836 22682 3840
rect 22618 3780 22622 3836
rect 22622 3780 22678 3836
rect 22678 3780 22682 3836
rect 22618 3776 22682 3780
rect 22698 3836 22762 3840
rect 22698 3780 22702 3836
rect 22702 3780 22758 3836
rect 22758 3780 22762 3836
rect 22698 3776 22762 3780
rect 22778 3836 22842 3840
rect 22778 3780 22782 3836
rect 22782 3780 22838 3836
rect 22838 3780 22842 3836
rect 22778 3776 22842 3780
rect 22858 3836 22922 3840
rect 22858 3780 22862 3836
rect 22862 3780 22918 3836
rect 22918 3780 22922 3836
rect 22858 3776 22922 3780
rect 37062 3836 37126 3840
rect 37062 3780 37066 3836
rect 37066 3780 37122 3836
rect 37122 3780 37126 3836
rect 37062 3776 37126 3780
rect 37142 3836 37206 3840
rect 37142 3780 37146 3836
rect 37146 3780 37202 3836
rect 37202 3780 37206 3836
rect 37142 3776 37206 3780
rect 37222 3836 37286 3840
rect 37222 3780 37226 3836
rect 37226 3780 37282 3836
rect 37282 3780 37286 3836
rect 37222 3776 37286 3780
rect 37302 3836 37366 3840
rect 37302 3780 37306 3836
rect 37306 3780 37362 3836
rect 37362 3780 37366 3836
rect 37302 3776 37366 3780
rect 51506 3836 51570 3840
rect 51506 3780 51510 3836
rect 51510 3780 51566 3836
rect 51566 3780 51570 3836
rect 51506 3776 51570 3780
rect 51586 3836 51650 3840
rect 51586 3780 51590 3836
rect 51590 3780 51646 3836
rect 51646 3780 51650 3836
rect 51586 3776 51650 3780
rect 51666 3836 51730 3840
rect 51666 3780 51670 3836
rect 51670 3780 51726 3836
rect 51726 3780 51730 3836
rect 51666 3776 51730 3780
rect 51746 3836 51810 3840
rect 51746 3780 51750 3836
rect 51750 3780 51806 3836
rect 51806 3780 51810 3836
rect 51746 3776 51810 3780
rect 15396 3292 15460 3296
rect 15396 3236 15400 3292
rect 15400 3236 15456 3292
rect 15456 3236 15460 3292
rect 15396 3232 15460 3236
rect 15476 3292 15540 3296
rect 15476 3236 15480 3292
rect 15480 3236 15536 3292
rect 15536 3236 15540 3292
rect 15476 3232 15540 3236
rect 15556 3292 15620 3296
rect 15556 3236 15560 3292
rect 15560 3236 15616 3292
rect 15616 3236 15620 3292
rect 15556 3232 15620 3236
rect 15636 3292 15700 3296
rect 15636 3236 15640 3292
rect 15640 3236 15696 3292
rect 15696 3236 15700 3292
rect 15636 3232 15700 3236
rect 29840 3292 29904 3296
rect 29840 3236 29844 3292
rect 29844 3236 29900 3292
rect 29900 3236 29904 3292
rect 29840 3232 29904 3236
rect 29920 3292 29984 3296
rect 29920 3236 29924 3292
rect 29924 3236 29980 3292
rect 29980 3236 29984 3292
rect 29920 3232 29984 3236
rect 30000 3292 30064 3296
rect 30000 3236 30004 3292
rect 30004 3236 30060 3292
rect 30060 3236 30064 3292
rect 30000 3232 30064 3236
rect 30080 3292 30144 3296
rect 30080 3236 30084 3292
rect 30084 3236 30140 3292
rect 30140 3236 30144 3292
rect 30080 3232 30144 3236
rect 44284 3292 44348 3296
rect 44284 3236 44288 3292
rect 44288 3236 44344 3292
rect 44344 3236 44348 3292
rect 44284 3232 44348 3236
rect 44364 3292 44428 3296
rect 44364 3236 44368 3292
rect 44368 3236 44424 3292
rect 44424 3236 44428 3292
rect 44364 3232 44428 3236
rect 44444 3292 44508 3296
rect 44444 3236 44448 3292
rect 44448 3236 44504 3292
rect 44504 3236 44508 3292
rect 44444 3232 44508 3236
rect 44524 3292 44588 3296
rect 44524 3236 44528 3292
rect 44528 3236 44584 3292
rect 44584 3236 44588 3292
rect 44524 3232 44588 3236
rect 58728 3292 58792 3296
rect 58728 3236 58732 3292
rect 58732 3236 58788 3292
rect 58788 3236 58792 3292
rect 58728 3232 58792 3236
rect 58808 3292 58872 3296
rect 58808 3236 58812 3292
rect 58812 3236 58868 3292
rect 58868 3236 58872 3292
rect 58808 3232 58872 3236
rect 58888 3292 58952 3296
rect 58888 3236 58892 3292
rect 58892 3236 58948 3292
rect 58948 3236 58952 3292
rect 58888 3232 58952 3236
rect 58968 3292 59032 3296
rect 58968 3236 58972 3292
rect 58972 3236 59028 3292
rect 59028 3236 59032 3292
rect 58968 3232 59032 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 22618 2748 22682 2752
rect 22618 2692 22622 2748
rect 22622 2692 22678 2748
rect 22678 2692 22682 2748
rect 22618 2688 22682 2692
rect 22698 2748 22762 2752
rect 22698 2692 22702 2748
rect 22702 2692 22758 2748
rect 22758 2692 22762 2748
rect 22698 2688 22762 2692
rect 22778 2748 22842 2752
rect 22778 2692 22782 2748
rect 22782 2692 22838 2748
rect 22838 2692 22842 2748
rect 22778 2688 22842 2692
rect 22858 2748 22922 2752
rect 22858 2692 22862 2748
rect 22862 2692 22918 2748
rect 22918 2692 22922 2748
rect 22858 2688 22922 2692
rect 37062 2748 37126 2752
rect 37062 2692 37066 2748
rect 37066 2692 37122 2748
rect 37122 2692 37126 2748
rect 37062 2688 37126 2692
rect 37142 2748 37206 2752
rect 37142 2692 37146 2748
rect 37146 2692 37202 2748
rect 37202 2692 37206 2748
rect 37142 2688 37206 2692
rect 37222 2748 37286 2752
rect 37222 2692 37226 2748
rect 37226 2692 37282 2748
rect 37282 2692 37286 2748
rect 37222 2688 37286 2692
rect 37302 2748 37366 2752
rect 37302 2692 37306 2748
rect 37306 2692 37362 2748
rect 37362 2692 37366 2748
rect 37302 2688 37366 2692
rect 51506 2748 51570 2752
rect 51506 2692 51510 2748
rect 51510 2692 51566 2748
rect 51566 2692 51570 2748
rect 51506 2688 51570 2692
rect 51586 2748 51650 2752
rect 51586 2692 51590 2748
rect 51590 2692 51646 2748
rect 51646 2692 51650 2748
rect 51586 2688 51650 2692
rect 51666 2748 51730 2752
rect 51666 2692 51670 2748
rect 51670 2692 51726 2748
rect 51726 2692 51730 2748
rect 51666 2688 51730 2692
rect 51746 2748 51810 2752
rect 51746 2692 51750 2748
rect 51750 2692 51806 2748
rect 51806 2692 51810 2748
rect 51746 2688 51810 2692
rect 15396 2204 15460 2208
rect 15396 2148 15400 2204
rect 15400 2148 15456 2204
rect 15456 2148 15460 2204
rect 15396 2144 15460 2148
rect 15476 2204 15540 2208
rect 15476 2148 15480 2204
rect 15480 2148 15536 2204
rect 15536 2148 15540 2204
rect 15476 2144 15540 2148
rect 15556 2204 15620 2208
rect 15556 2148 15560 2204
rect 15560 2148 15616 2204
rect 15616 2148 15620 2204
rect 15556 2144 15620 2148
rect 15636 2204 15700 2208
rect 15636 2148 15640 2204
rect 15640 2148 15696 2204
rect 15696 2148 15700 2204
rect 15636 2144 15700 2148
rect 29840 2204 29904 2208
rect 29840 2148 29844 2204
rect 29844 2148 29900 2204
rect 29900 2148 29904 2204
rect 29840 2144 29904 2148
rect 29920 2204 29984 2208
rect 29920 2148 29924 2204
rect 29924 2148 29980 2204
rect 29980 2148 29984 2204
rect 29920 2144 29984 2148
rect 30000 2204 30064 2208
rect 30000 2148 30004 2204
rect 30004 2148 30060 2204
rect 30060 2148 30064 2204
rect 30000 2144 30064 2148
rect 30080 2204 30144 2208
rect 30080 2148 30084 2204
rect 30084 2148 30140 2204
rect 30140 2148 30144 2204
rect 30080 2144 30144 2148
rect 44284 2204 44348 2208
rect 44284 2148 44288 2204
rect 44288 2148 44344 2204
rect 44344 2148 44348 2204
rect 44284 2144 44348 2148
rect 44364 2204 44428 2208
rect 44364 2148 44368 2204
rect 44368 2148 44424 2204
rect 44424 2148 44428 2204
rect 44364 2144 44428 2148
rect 44444 2204 44508 2208
rect 44444 2148 44448 2204
rect 44448 2148 44504 2204
rect 44504 2148 44508 2204
rect 44444 2144 44508 2148
rect 44524 2204 44588 2208
rect 44524 2148 44528 2204
rect 44528 2148 44584 2204
rect 44584 2148 44588 2204
rect 44524 2144 44588 2148
rect 58728 2204 58792 2208
rect 58728 2148 58732 2204
rect 58732 2148 58788 2204
rect 58788 2148 58792 2204
rect 58728 2144 58792 2148
rect 58808 2204 58872 2208
rect 58808 2148 58812 2204
rect 58812 2148 58868 2204
rect 58868 2148 58872 2204
rect 58808 2144 58872 2148
rect 58888 2204 58952 2208
rect 58888 2148 58892 2204
rect 58892 2148 58948 2204
rect 58948 2148 58952 2204
rect 58888 2144 58952 2148
rect 58968 2204 59032 2208
rect 58968 2148 58972 2204
rect 58972 2148 59028 2204
rect 59028 2148 59032 2204
rect 58968 2144 59032 2148
<< metal4 >>
rect 8166 21248 8486 21808
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 7235 7308 7301 7309
rect 7235 7244 7236 7308
rect 7300 7244 7301 7308
rect 7235 7243 7301 7244
rect 7238 5541 7298 7243
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 7235 5540 7301 5541
rect 7235 5476 7236 5540
rect 7300 5476 7301 5540
rect 7235 5475 7301 5476
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 2128 8486 2688
rect 15388 21792 15708 21808
rect 15388 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15708 21792
rect 15388 20704 15708 21728
rect 15388 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15708 20704
rect 15388 19616 15708 20640
rect 15388 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15708 19616
rect 15388 18528 15708 19552
rect 15388 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15708 18528
rect 15388 17440 15708 18464
rect 15388 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15708 17440
rect 15388 16352 15708 17376
rect 15388 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15708 16352
rect 15388 15264 15708 16288
rect 15388 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15708 15264
rect 15388 14176 15708 15200
rect 15388 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15708 14176
rect 15388 13088 15708 14112
rect 15388 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15708 13088
rect 15388 12000 15708 13024
rect 15388 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15708 12000
rect 15388 10912 15708 11936
rect 15388 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15708 10912
rect 15388 9824 15708 10848
rect 15388 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15708 9824
rect 15388 8736 15708 9760
rect 15388 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15708 8736
rect 15388 7648 15708 8672
rect 15388 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15708 7648
rect 15388 6560 15708 7584
rect 15388 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15708 6560
rect 15388 5472 15708 6496
rect 15388 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15708 5472
rect 15388 4384 15708 5408
rect 15388 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15708 4384
rect 15388 3296 15708 4320
rect 15388 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15708 3296
rect 15388 2208 15708 3232
rect 15388 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15708 2208
rect 15388 2128 15708 2144
rect 22610 21248 22930 21808
rect 22610 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22930 21248
rect 22610 20160 22930 21184
rect 22610 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22930 20160
rect 22610 19072 22930 20096
rect 22610 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22930 19072
rect 22610 17984 22930 19008
rect 22610 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22930 17984
rect 22610 16896 22930 17920
rect 22610 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22930 16896
rect 22610 15808 22930 16832
rect 22610 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22930 15808
rect 22610 14720 22930 15744
rect 22610 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22930 14720
rect 22610 13632 22930 14656
rect 22610 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22930 13632
rect 22610 12544 22930 13568
rect 22610 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22930 12544
rect 22610 11456 22930 12480
rect 22610 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22930 11456
rect 22610 10368 22930 11392
rect 22610 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22930 10368
rect 22610 9280 22930 10304
rect 22610 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22930 9280
rect 22610 8192 22930 9216
rect 22610 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22930 8192
rect 22610 7104 22930 8128
rect 22610 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22930 7104
rect 22610 6016 22930 7040
rect 22610 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22930 6016
rect 22610 4928 22930 5952
rect 22610 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22930 4928
rect 22610 3840 22930 4864
rect 22610 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22930 3840
rect 22610 2752 22930 3776
rect 22610 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22930 2752
rect 22610 2128 22930 2688
rect 29832 21792 30152 21808
rect 29832 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30152 21792
rect 29832 20704 30152 21728
rect 29832 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30152 20704
rect 29832 19616 30152 20640
rect 29832 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30152 19616
rect 29832 18528 30152 19552
rect 29832 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30152 18528
rect 29832 17440 30152 18464
rect 29832 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30152 17440
rect 29832 16352 30152 17376
rect 37054 21248 37374 21808
rect 37054 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37374 21248
rect 37054 20160 37374 21184
rect 37054 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37374 20160
rect 37054 19072 37374 20096
rect 37054 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37374 19072
rect 37054 17984 37374 19008
rect 37054 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37374 17984
rect 37054 16896 37374 17920
rect 37054 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37374 16896
rect 35571 16692 35637 16693
rect 35571 16628 35572 16692
rect 35636 16628 35637 16692
rect 35571 16627 35637 16628
rect 29832 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30152 16352
rect 29832 15264 30152 16288
rect 29832 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30152 15264
rect 29832 14176 30152 15200
rect 29832 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30152 14176
rect 29832 13088 30152 14112
rect 29832 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30152 13088
rect 29832 12000 30152 13024
rect 29832 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30152 12000
rect 29832 10912 30152 11936
rect 29832 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30152 10912
rect 29832 9824 30152 10848
rect 29832 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30152 9824
rect 29832 8736 30152 9760
rect 29832 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30152 8736
rect 29832 7648 30152 8672
rect 29832 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30152 7648
rect 29832 6560 30152 7584
rect 29832 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30152 6560
rect 29832 5472 30152 6496
rect 29832 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30152 5472
rect 29832 4384 30152 5408
rect 29832 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30152 4384
rect 29832 3296 30152 4320
rect 35574 3909 35634 16627
rect 37054 15808 37374 16832
rect 37054 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37374 15808
rect 37054 14720 37374 15744
rect 37054 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37374 14720
rect 37054 13632 37374 14656
rect 37054 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37374 13632
rect 37054 12544 37374 13568
rect 37054 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37374 12544
rect 37054 11456 37374 12480
rect 37054 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37374 11456
rect 37054 10368 37374 11392
rect 37054 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37374 10368
rect 37054 9280 37374 10304
rect 37054 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37374 9280
rect 37054 8192 37374 9216
rect 37054 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37374 8192
rect 37054 7104 37374 8128
rect 37054 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37374 7104
rect 37054 6016 37374 7040
rect 37054 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37374 6016
rect 37054 4928 37374 5952
rect 37054 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37374 4928
rect 35571 3908 35637 3909
rect 35571 3844 35572 3908
rect 35636 3844 35637 3908
rect 35571 3843 35637 3844
rect 29832 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30152 3296
rect 29832 2208 30152 3232
rect 29832 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30152 2208
rect 29832 2128 30152 2144
rect 37054 3840 37374 4864
rect 37054 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37374 3840
rect 37054 2752 37374 3776
rect 37054 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37374 2752
rect 37054 2128 37374 2688
rect 44276 21792 44596 21808
rect 44276 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44596 21792
rect 44276 20704 44596 21728
rect 44276 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44596 20704
rect 44276 19616 44596 20640
rect 44276 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44596 19616
rect 44276 18528 44596 19552
rect 44276 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44596 18528
rect 44276 17440 44596 18464
rect 44276 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44596 17440
rect 44276 16352 44596 17376
rect 44276 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44596 16352
rect 44276 15264 44596 16288
rect 44276 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44596 15264
rect 44276 14176 44596 15200
rect 44276 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44596 14176
rect 44276 13088 44596 14112
rect 44276 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44596 13088
rect 44276 12000 44596 13024
rect 44276 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44596 12000
rect 44276 10912 44596 11936
rect 44276 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44596 10912
rect 44276 9824 44596 10848
rect 44276 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44596 9824
rect 44276 8736 44596 9760
rect 44276 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44596 8736
rect 44276 7648 44596 8672
rect 44276 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44596 7648
rect 44276 6560 44596 7584
rect 44276 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44596 6560
rect 44276 5472 44596 6496
rect 44276 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44596 5472
rect 44276 4384 44596 5408
rect 44276 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44596 4384
rect 44276 3296 44596 4320
rect 44276 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44596 3296
rect 44276 2208 44596 3232
rect 44276 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44596 2208
rect 44276 2128 44596 2144
rect 51498 21248 51818 21808
rect 51498 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51818 21248
rect 51498 20160 51818 21184
rect 51498 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51818 20160
rect 51498 19072 51818 20096
rect 51498 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51818 19072
rect 51498 17984 51818 19008
rect 51498 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51818 17984
rect 51498 16896 51818 17920
rect 51498 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51818 16896
rect 51498 15808 51818 16832
rect 51498 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51818 15808
rect 51498 14720 51818 15744
rect 51498 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51818 14720
rect 51498 13632 51818 14656
rect 51498 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51818 13632
rect 51498 12544 51818 13568
rect 51498 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51818 12544
rect 51498 11456 51818 12480
rect 51498 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51818 11456
rect 51498 10368 51818 11392
rect 51498 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51818 10368
rect 51498 9280 51818 10304
rect 51498 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51818 9280
rect 51498 8192 51818 9216
rect 51498 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51818 8192
rect 51498 7104 51818 8128
rect 51498 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51818 7104
rect 51498 6016 51818 7040
rect 58720 21792 59040 21808
rect 58720 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59040 21792
rect 58720 20704 59040 21728
rect 58720 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59040 20704
rect 58720 19616 59040 20640
rect 58720 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59040 19616
rect 58720 18528 59040 19552
rect 58720 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59040 18528
rect 58720 17440 59040 18464
rect 58720 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59040 17440
rect 58720 16352 59040 17376
rect 58720 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59040 16352
rect 58720 15264 59040 16288
rect 58720 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59040 15264
rect 58720 14176 59040 15200
rect 58720 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59040 14176
rect 58720 13088 59040 14112
rect 58720 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59040 13088
rect 58720 12000 59040 13024
rect 58720 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59040 12000
rect 58720 10912 59040 11936
rect 58720 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59040 10912
rect 58720 9824 59040 10848
rect 58720 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59040 9824
rect 58720 8736 59040 9760
rect 58720 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59040 8736
rect 58720 7648 59040 8672
rect 58720 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59040 7648
rect 55995 7036 56061 7037
rect 55995 6972 55996 7036
rect 56060 6972 56061 7036
rect 55995 6971 56061 6972
rect 51498 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51818 6016
rect 51498 4928 51818 5952
rect 51498 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51818 4928
rect 51498 3840 51818 4864
rect 55998 4045 56058 6971
rect 58720 6560 59040 7584
rect 58720 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59040 6560
rect 58720 5472 59040 6496
rect 58720 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59040 5472
rect 58720 4384 59040 5408
rect 58720 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59040 4384
rect 55995 4044 56061 4045
rect 55995 3980 55996 4044
rect 56060 3980 56061 4044
rect 55995 3979 56061 3980
rect 51498 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51818 3840
rect 51498 2752 51818 3776
rect 51498 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51818 2752
rect 51498 2128 51818 2688
rect 58720 3296 59040 4320
rect 58720 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59040 3296
rect 58720 2208 59040 3232
rect 58720 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59040 2208
rect 58720 2128 59040 2144
use sky130_fd_sc_hd__or4bb_1  _0414_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 55108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0415_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 48944 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0416_
timestamp 1688980957
transform -1 0 43700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0417_
timestamp 1688980957
transform -1 0 23460 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0418_
timestamp 1688980957
transform -1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0419_
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0420_
timestamp 1688980957
transform -1 0 35604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0421_
timestamp 1688980957
transform 1 0 27324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0422_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42872 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0423_
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0424_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0425_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _0426_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0427_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6348 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0428_
timestamp 1688980957
transform -1 0 6440 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0429_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0430_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7176 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0431_
timestamp 1688980957
transform -1 0 6072 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0432_
timestamp 1688980957
transform -1 0 8096 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0433_
timestamp 1688980957
transform -1 0 8004 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0434_
timestamp 1688980957
transform -1 0 7820 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0435_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0436_
timestamp 1688980957
transform -1 0 8832 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0437_
timestamp 1688980957
transform -1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0438_
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0439_
timestamp 1688980957
transform -1 0 13984 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0440_
timestamp 1688980957
transform -1 0 13800 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0441_
timestamp 1688980957
transform 1 0 12880 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0442_
timestamp 1688980957
transform -1 0 12788 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0443_
timestamp 1688980957
transform -1 0 14536 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0444_
timestamp 1688980957
transform -1 0 14628 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0445_
timestamp 1688980957
transform -1 0 14904 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0446_
timestamp 1688980957
transform -1 0 15364 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0447_
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0448_
timestamp 1688980957
transform -1 0 14352 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0449_
timestamp 1688980957
transform -1 0 14904 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0450_
timestamp 1688980957
transform -1 0 15548 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0451_
timestamp 1688980957
transform -1 0 16652 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0452_
timestamp 1688980957
transform -1 0 17480 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0453_
timestamp 1688980957
transform -1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0454_
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0455_
timestamp 1688980957
transform -1 0 20240 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0456_
timestamp 1688980957
transform -1 0 21160 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0457_
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0458_
timestamp 1688980957
transform -1 0 19780 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0459_
timestamp 1688980957
transform -1 0 20240 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0460_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0461_
timestamp 1688980957
transform -1 0 21068 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0462_
timestamp 1688980957
transform -1 0 22816 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0463_
timestamp 1688980957
transform -1 0 21528 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0464_
timestamp 1688980957
transform -1 0 21620 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0465_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0466_
timestamp 1688980957
transform 1 0 21896 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0467_
timestamp 1688980957
transform -1 0 26312 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0468_
timestamp 1688980957
transform -1 0 26312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0469_
timestamp 1688980957
transform 1 0 24380 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0470_
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0471_
timestamp 1688980957
transform -1 0 24748 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0472_
timestamp 1688980957
transform -1 0 24932 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0473_
timestamp 1688980957
transform -1 0 25392 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0474_
timestamp 1688980957
transform -1 0 27232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0475_
timestamp 1688980957
transform -1 0 26864 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0476_
timestamp 1688980957
transform -1 0 26864 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0477_
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0478_
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0479_
timestamp 1688980957
transform -1 0 27784 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0480_
timestamp 1688980957
transform -1 0 27600 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0481_
timestamp 1688980957
transform -1 0 28152 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0482_
timestamp 1688980957
transform 1 0 28152 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0483_
timestamp 1688980957
transform -1 0 32016 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0484_
timestamp 1688980957
transform -1 0 31832 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0485_
timestamp 1688980957
transform -1 0 31740 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0486_
timestamp 1688980957
transform -1 0 31924 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0487_
timestamp 1688980957
transform -1 0 32016 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0488_
timestamp 1688980957
transform -1 0 32844 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0489_
timestamp 1688980957
transform -1 0 33764 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0490_
timestamp 1688980957
transform -1 0 34408 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0491_
timestamp 1688980957
transform -1 0 34224 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0492_
timestamp 1688980957
transform -1 0 34132 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1688980957
transform 1 0 34408 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0494_
timestamp 1688980957
transform 1 0 33764 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0495_
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0496_
timestamp 1688980957
transform -1 0 37904 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0497_
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0498_
timestamp 1688980957
transform 1 0 35696 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0499_
timestamp 1688980957
transform -1 0 34408 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0500_
timestamp 1688980957
transform -1 0 34224 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0501_
timestamp 1688980957
transform -1 0 35512 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0502_
timestamp 1688980957
transform 1 0 36616 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0503_
timestamp 1688980957
transform 1 0 37444 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0504_
timestamp 1688980957
transform -1 0 39652 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0505_
timestamp 1688980957
transform 1 0 39284 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0506_
timestamp 1688980957
transform 1 0 39192 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0507_
timestamp 1688980957
transform -1 0 39468 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0508_
timestamp 1688980957
transform 1 0 37812 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0509_
timestamp 1688980957
transform -1 0 40112 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0510_
timestamp 1688980957
transform -1 0 42044 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0511_
timestamp 1688980957
transform 1 0 40572 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0512_
timestamp 1688980957
transform -1 0 43332 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0513_
timestamp 1688980957
transform -1 0 43240 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0514_
timestamp 1688980957
transform -1 0 44160 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0515_
timestamp 1688980957
transform -1 0 44344 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0516_
timestamp 1688980957
transform -1 0 44344 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1688980957
transform -1 0 44160 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0518_
timestamp 1688980957
transform 1 0 43700 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0519_
timestamp 1688980957
transform -1 0 44896 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0520_
timestamp 1688980957
transform -1 0 44988 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1688980957
transform 1 0 44988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0522_
timestamp 1688980957
transform 1 0 44160 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0523_
timestamp 1688980957
transform -1 0 48116 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0524_
timestamp 1688980957
transform -1 0 48576 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1688980957
transform -1 0 48392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0526_
timestamp 1688980957
transform -1 0 48760 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0527_
timestamp 1688980957
transform -1 0 49496 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0528_
timestamp 1688980957
transform -1 0 49496 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0529_
timestamp 1688980957
transform -1 0 49496 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0530_
timestamp 1688980957
transform -1 0 50692 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0531_
timestamp 1688980957
transform -1 0 50692 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0532_
timestamp 1688980957
transform -1 0 50692 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0533_
timestamp 1688980957
transform -1 0 51796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0534_
timestamp 1688980957
transform -1 0 52624 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0535_
timestamp 1688980957
transform -1 0 50324 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0536_
timestamp 1688980957
transform -1 0 50784 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0537_
timestamp 1688980957
transform -1 0 51152 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0538_
timestamp 1688980957
transform 1 0 51428 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0539_
timestamp 1688980957
transform -1 0 56120 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0540_
timestamp 1688980957
transform -1 0 56396 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0541_
timestamp 1688980957
transform 1 0 55292 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0542_
timestamp 1688980957
transform 1 0 53636 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0543_
timestamp 1688980957
transform -1 0 56028 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0544_
timestamp 1688980957
transform -1 0 56212 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0545_
timestamp 1688980957
transform 1 0 56028 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0546_
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0547_
timestamp 1688980957
transform -1 0 57224 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0548_
timestamp 1688980957
transform -1 0 57224 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0549_
timestamp 1688980957
transform 1 0 57224 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0550_
timestamp 1688980957
transform -1 0 57592 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0551_
timestamp 1688980957
transform -1 0 55844 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0552_
timestamp 1688980957
transform -1 0 55752 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0553_
timestamp 1688980957
transform -1 0 56212 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0554_
timestamp 1688980957
transform -1 0 58420 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0555_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0556_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0557_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1688980957
transform -1 0 28336 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1688980957
transform 1 0 33580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1688980957
transform -1 0 32936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1688980957
transform -1 0 35512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1688980957
transform -1 0 36984 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1688980957
transform -1 0 33672 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1688980957
transform -1 0 39560 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1688980957
transform -1 0 39744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1688980957
transform 1 0 40020 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1688980957
transform -1 0 44160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1688980957
transform -1 0 44804 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1688980957
transform -1 0 51336 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1688980957
transform 1 0 47840 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1688980957
transform -1 0 50048 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1688980957
transform 1 0 48668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1688980957
transform 1 0 56488 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1688980957
transform -1 0 57408 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 1688980957
transform -1 0 57224 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1688980957
transform -1 0 56120 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0577_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_4  _0578_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1688980957
transform -1 0 8464 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1688980957
transform -1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 1688980957
transform -1 0 9752 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1688980957
transform -1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1688980957
transform -1 0 21528 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1688980957
transform -1 0 21528 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1688980957
transform -1 0 22264 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1688980957
transform 1 0 25208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1688980957
transform 1 0 27416 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1688980957
transform -1 0 26864 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1688980957
transform -1 0 33028 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1688980957
transform -1 0 32936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform 1 0 37628 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1688980957
transform -1 0 35512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1688980957
transform 1 0 37628 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1688980957
transform 1 0 38364 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform -1 0 43240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform -1 0 44804 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1688980957
transform 1 0 49128 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1688980957
transform -1 0 49956 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform -1 0 51520 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1688980957
transform -1 0 50968 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform -1 0 58144 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1688980957
transform -1 0 57684 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform -1 0 57316 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1688980957
transform -1 0 57500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0611_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0612_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4416 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0613_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1688980957
transform -1 0 5888 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1688980957
transform -1 0 12328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1688980957
transform 1 0 14536 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform 1 0 18032 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform 1 0 17756 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform 1 0 28152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1688980957
transform -1 0 29440 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform -1 0 32108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1688980957
transform -1 0 36524 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform 1 0 30360 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1688980957
transform -1 0 38180 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform 1 0 41032 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform 1 0 42596 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1688980957
transform 1 0 42320 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform 1 0 46460 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1688980957
transform -1 0 47564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1688980957
transform -1 0 48392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform -1 0 54924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform 1 0 51796 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform 1 0 54280 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1688980957
transform -1 0 52992 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0646_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0647_
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0648_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0649_
timestamp 1688980957
transform -1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0650_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5796 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0651_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0652_
timestamp 1688980957
transform -1 0 6532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0653_
timestamp 1688980957
transform -1 0 6992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0654_
timestamp 1688980957
transform -1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0655_
timestamp 1688980957
transform -1 0 3680 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0656_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0657_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0658_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0659_
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0660_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5244 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0661_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0662_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0663_
timestamp 1688980957
transform -1 0 4140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0664_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4968 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 1688980957
transform -1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0666_
timestamp 1688980957
transform -1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0667_
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0668_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 1688980957
transform 1 0 3220 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1688980957
transform -1 0 4600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0674_
timestamp 1688980957
transform -1 0 12328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1688980957
transform -1 0 18584 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1688980957
transform 1 0 16928 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1688980957
transform -1 0 22632 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0682_
timestamp 1688980957
transform 1 0 25392 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform -1 0 29440 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0685_
timestamp 1688980957
transform 1 0 30452 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1688980957
transform 1 0 35696 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1688980957
transform 1 0 31556 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform -1 0 37812 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1688980957
transform 1 0 36340 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1688980957
transform 1 0 38916 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 41768 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 42596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1688980957
transform 1 0 46092 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1688980957
transform 1 0 45540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform 1 0 47564 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform 1 0 46552 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1688980957
transform 1 0 53820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1688980957
transform 1 0 52716 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1688980957
transform -1 0 55016 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 52256 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_4  _0701_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1688980957
transform 1 0 4232 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1688980957
transform -1 0 11408 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform -1 0 17940 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1688980957
transform 1 0 18124 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1688980957
transform 1 0 23460 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 1688980957
transform 1 0 20424 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1688980957
transform -1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1688980957
transform 1 0 28428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform 1 0 30452 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1688980957
transform 1 0 34868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform -1 0 32016 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform 1 0 36524 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1688980957
transform -1 0 43240 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1688980957
transform 1 0 42688 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1688980957
transform 1 0 45632 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1688980957
transform 1 0 45908 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform -1 0 48392 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1688980957
transform -1 0 47932 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1688980957
transform 1 0 53268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1688980957
transform -1 0 53452 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform 1 0 53268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 1688980957
transform -1 0 53544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0734_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1688980957
transform 1 0 7912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1688980957
transform 1 0 7728 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1688980957
transform -1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1688980957
transform -1 0 15088 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1688980957
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform -1 0 19964 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform -1 0 22632 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 1688980957
transform 1 0 25576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1688980957
transform 1 0 28428 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1688980957
transform 1 0 30544 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1688980957
transform -1 0 33672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform 1 0 37904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1688980957
transform -1 0 35052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1688980957
transform 1 0 38548 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1688980957
transform -1 0 39560 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0757_
timestamp 1688980957
transform 1 0 42688 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1688980957
transform -1 0 44344 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 1688980957
transform -1 0 49772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform -1 0 49404 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform -1 0 50968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1688980957
transform -1 0 50968 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1688980957
transform -1 0 57224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1688980957
transform 1 0 55660 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1688980957
transform -1 0 58052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1688980957
transform -1 0 56120 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _0767_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1688980957
transform 1 0 8004 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1688980957
transform -1 0 9752 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1688980957
transform 1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform -1 0 15364 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1688980957
transform -1 0 15272 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1688980957
transform -1 0 21068 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1688980957
transform -1 0 20884 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1688980957
transform 1 0 25208 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1688980957
transform 1 0 25392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform -1 0 28336 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1688980957
transform -1 0 32844 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1688980957
transform -1 0 33212 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1688980957
transform 1 0 34224 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform -1 0 39560 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1688980957
transform -1 0 34132 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1688980957
transform -1 0 40480 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1688980957
transform -1 0 40664 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 42320 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1688980957
transform 1 0 43884 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1688980957
transform -1 0 45816 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1688980957
transform -1 0 50968 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform -1 0 49956 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1688980957
transform -1 0 51520 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1688980957
transform 1 0 50968 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1688980957
transform 1 0 56488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1688980957
transform -1 0 57500 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1688980957
transform -1 0 57408 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1688980957
transform 1 0 56120 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0800_
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0801_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 5152 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0803_
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1688980957
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0805_
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0806_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0807_
timestamp 1688980957
transform -1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0809_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0810_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0812_
timestamp 1688980957
transform -1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0813_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0814_
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0815_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform 1 0 2944 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform -1 0 3588 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1688980957
transform 1 0 16928 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1688980957
transform -1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 1688980957
transform 1 0 22632 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1688980957
transform -1 0 21620 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1688980957
transform -1 0 25024 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1688980957
transform 1 0 28520 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 1688980957
transform -1 0 32108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1688980957
transform 1 0 35236 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 1688980957
transform 1 0 30728 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1688980957
transform 1 0 36800 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1688980957
transform 1 0 35880 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1688980957
transform -1 0 40664 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 1688980957
transform 1 0 41768 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1688980957
transform 1 0 45264 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 1688980957
transform -1 0 47104 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp 1688980957
transform -1 0 48392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1688980957
transform 1 0 52992 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1688980957
transform -1 0 53544 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1688980957
transform 1 0 53176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0847_
timestamp 1688980957
transform -1 0 53544 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1688980957
transform -1 0 6256 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1688980957
transform 1 0 6440 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1688980957
transform -1 0 13708 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1688980957
transform 1 0 13156 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1688980957
transform -1 0 13800 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1688980957
transform -1 0 15916 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1688980957
transform -1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1688980957
transform 1 0 26312 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1688980957
transform 1 0 23276 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1688980957
transform 1 0 28612 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _0861_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29256 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1688980957
transform -1 0 33580 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1688980957
transform -1 0 32568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1688980957
transform 1 0 32936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1688980957
transform -1 0 37076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1688980957
transform 1 0 32292 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1688980957
transform -1 0 39284 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1688980957
transform -1 0 41308 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1688980957
transform 1 0 38548 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1688980957
transform -1 0 44436 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1688980957
transform 1 0 43884 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1688980957
transform -1 0 50508 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1688980957
transform 1 0 47288 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1688980957
transform 1 0 49220 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1688980957
transform 1 0 48116 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1688980957
transform 1 0 56212 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1688980957
transform -1 0 57960 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1688980957
transform 1 0 56120 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1688980957
transform 1 0 55844 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1688980957
transform -1 0 8648 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1688980957
transform -1 0 9384 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1688980957
transform -1 0 9752 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1688980957
transform -1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1688980957
transform -1 0 16100 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1688980957
transform -1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1688980957
transform -1 0 18492 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1688980957
transform -1 0 21712 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1688980957
transform -1 0 21620 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1688980957
transform -1 0 21712 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1688980957
transform -1 0 26680 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1688980957
transform -1 0 26404 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1688980957
transform 1 0 27140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1688980957
transform 1 0 26220 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1688980957
transform -1 0 33396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1688980957
transform -1 0 33580 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1688980957
transform -1 0 35420 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1688980957
transform -1 0 37628 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1688980957
transform -1 0 35880 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1688980957
transform -1 0 38732 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1688980957
transform 1 0 37536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1688980957
transform -1 0 43976 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1688980957
transform 1 0 42872 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1688980957
transform 1 0 43424 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1688980957
transform 1 0 48760 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1688980957
transform -1 0 50968 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1688980957
transform -1 0 52164 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1688980957
transform -1 0 51612 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1688980957
transform -1 0 57776 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1688980957
transform -1 0 57408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1688980957
transform 1 0 56304 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1688980957
transform 1 0 56304 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1688980957
transform 1 0 2208 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1688980957
transform 1 0 4324 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1688980957
transform 1 0 4508 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1688980957
transform 1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1688980957
transform 1 0 10856 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1688980957
transform 1 0 16836 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1688980957
transform 1 0 17112 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1688980957
transform 1 0 21988 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1688980957
transform 1 0 23460 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1688980957
transform -1 0 24196 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1688980957
transform 1 0 27416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1688980957
transform -1 0 31464 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1688980957
transform 1 0 29808 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1688980957
transform 1 0 29716 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1688980957
transform 1 0 36064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1688980957
transform 1 0 36064 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1688980957
transform 1 0 40388 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1688980957
transform 1 0 41124 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1688980957
transform 1 0 40848 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1688980957
transform 1 0 45172 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1688980957
transform 1 0 45356 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1688980957
transform 1 0 46368 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1688980957
transform 1 0 46000 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1688980957
transform 1 0 52992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1688980957
transform 1 0 51704 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1688980957
transform 1 0 52900 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1688980957
transform 1 0 51520 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1688980957
transform -1 0 7820 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1688980957
transform 1 0 10120 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1688980957
transform -1 0 11592 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1688980957
transform 1 0 11868 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1688980957
transform 1 0 16100 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1688980957
transform 1 0 16928 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1688980957
transform 1 0 22172 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1688980957
transform 1 0 23460 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1688980957
transform 1 0 27968 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1688980957
transform 1 0 35144 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1688980957
transform 1 0 30176 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1688980957
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1688980957
transform 1 0 38916 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1688980957
transform 1 0 40296 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1688980957
transform 1 0 47656 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1688980957
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1688980957
transform 1 0 52532 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1688980957
transform 1 0 52072 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1688980957
transform 1 0 52808 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1688980957
transform 1 0 51612 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1688980957
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1688980957
transform 1 0 2116 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1688980957
transform 1 0 4140 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1688980957
transform 1 0 9476 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1688980957
transform 1 0 13064 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1688980957
transform 1 0 17112 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1688980957
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1688980957
transform 1 0 19688 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1688980957
transform 1 0 23460 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1688980957
transform 1 0 23552 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1688980957
transform 1 0 28520 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1688980957
transform 1 0 29808 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1688980957
transform 1 0 34224 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1688980957
transform -1 0 31188 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1688980957
transform 1 0 35696 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1688980957
transform 1 0 35696 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1688980957
transform 1 0 38824 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1688980957
transform 1 0 40848 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1688980957
transform 1 0 41216 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1688980957
transform 1 0 45080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1688980957
transform 1 0 45908 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1688980957
transform 1 0 47840 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1688980957
transform 1 0 46460 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1688980957
transform 1 0 52900 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1688980957
transform 1 0 52808 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1688980957
transform 1 0 51152 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1688980957
transform -1 0 7912 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1688980957
transform -1 0 8464 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1688980957
transform 1 0 7268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1688980957
transform -1 0 14536 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1688980957
transform -1 0 15548 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1688980957
transform -1 0 20700 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1688980957
transform 1 0 25300 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1688980957
transform 1 0 22540 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1688980957
transform 1 0 26312 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1688980957
transform 1 0 25300 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1688980957
transform -1 0 33580 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1688980957
transform -1 0 34224 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1688980957
transform -1 0 38732 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1688980957
transform 1 0 32568 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1688980957
transform 1 0 37996 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1688980957
transform -1 0 39652 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1688980957
transform 1 0 41860 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1688980957
transform 1 0 42964 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1688980957
transform -1 0 50048 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1688980957
transform 1 0 48116 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1688980957
transform -1 0 50876 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1688980957
transform -1 0 52256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1688980957
transform -1 0 57684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1688980957
transform 1 0 56120 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1688980957
transform 1 0 55752 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1688980957
transform 1 0 7360 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1688980957
transform -1 0 9016 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1688980957
transform -1 0 10304 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1688980957
transform -1 0 14444 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1688980957
transform -1 0 16100 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1688980957
transform -1 0 15824 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1688980957
transform -1 0 18400 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1688980957
transform -1 0 21252 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1688980957
transform -1 0 21160 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1688980957
transform 1 0 24564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1688980957
transform -1 0 26680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1688980957
transform -1 0 29072 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1688980957
transform -1 0 33580 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1688980957
transform -1 0 33580 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 32936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform -1 0 39008 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform -1 0 34316 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform -1 0 41308 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform -1 0 40204 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 42320 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform -1 0 46460 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform -1 0 50324 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform -1 0 50968 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform -1 0 51612 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform -1 0 51612 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1688980957
transform 1 0 56304 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1688980957
transform -1 0 57776 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1688980957
transform 1 0 56304 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1688980957
transform -1 0 3404 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1077_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform -1 0 10948 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1080_
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform 1 0 2116 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform -1 0 3404 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 2944 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1688980957
transform 1 0 16928 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform 1 0 21988 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1688980957
transform 1 0 23368 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1688980957
transform 1 0 27876 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1688980957
transform 1 0 27692 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1688980957
transform 1 0 29808 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1688980957
transform 1 0 30084 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1688980957
transform 1 0 35696 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1688980957
transform 1 0 39100 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1688980957
transform 1 0 40296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1688980957
transform 1 0 41308 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1688980957
transform 1 0 44528 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1688980957
transform 1 0 44804 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1688980957
transform 1 0 46184 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1688980957
transform -1 0 47288 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1688980957
transform 1 0 52716 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1688980957
transform 1 0 51152 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1688980957
transform 1 0 3956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform -1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1688980957
transform -1 0 14628 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1688980957
transform 1 0 12512 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1688980957
transform -1 0 13892 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1688980957
transform 1 0 17664 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1688980957
transform 1 0 27048 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__C asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0426__B
timestamp 1688980957
transform -1 0 7728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__S0
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__S1
timestamp 1688980957
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__S0
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__S1
timestamp 1688980957
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0429__S
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__A
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__S0
timestamp 1688980957
transform -1 0 2208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__S1
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__S0
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__S1
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0433__S
timestamp 1688980957
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__A
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__S0
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__S1
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__S0
timestamp 1688980957
transform -1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__S1
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0437__S
timestamp 1688980957
transform 1 0 9936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A
timestamp 1688980957
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__S0
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__S1
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__S0
timestamp 1688980957
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__S1
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__S
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__A
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__S0
timestamp 1688980957
transform 1 0 12420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__S1
timestamp 1688980957
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__S0
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__S1
timestamp 1688980957
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__S
timestamp 1688980957
transform -1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__A
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S0
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S1
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__S0
timestamp 1688980957
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__S1
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__S
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__A
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S0
timestamp 1688980957
transform -1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S1
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__S0
timestamp 1688980957
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__S1
timestamp 1688980957
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__S
timestamp 1688980957
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__A
timestamp 1688980957
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S0
timestamp 1688980957
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S1
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__S0
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__S1
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0457__S
timestamp 1688980957
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S0
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S1
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__S0
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__S1
timestamp 1688980957
transform 1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__S
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__A
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S0
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S1
timestamp 1688980957
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__S0
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__S1
timestamp 1688980957
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__S
timestamp 1688980957
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__A
timestamp 1688980957
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S0
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S1
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__S0
timestamp 1688980957
transform 1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__S1
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__S
timestamp 1688980957
transform 1 0 21252 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__A
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S0
timestamp 1688980957
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S1
timestamp 1688980957
transform 1 0 22724 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__S0
timestamp 1688980957
transform 1 0 23184 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__S1
timestamp 1688980957
transform 1 0 22816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__S
timestamp 1688980957
transform 1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__A
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S0
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S1
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0476__S0
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0476__S1
timestamp 1688980957
transform -1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__S
timestamp 1688980957
transform 1 0 26404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__A
timestamp 1688980957
transform 1 0 28060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S0
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S1
timestamp 1688980957
transform 1 0 25760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__S0
timestamp 1688980957
transform 1 0 24748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__S1
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__S
timestamp 1688980957
transform 1 0 27140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__A
timestamp 1688980957
transform 1 0 27232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S0
timestamp 1688980957
transform 1 0 32660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S1
timestamp 1688980957
transform 1 0 31372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__S0
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__S1
timestamp 1688980957
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__S
timestamp 1688980957
transform 1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1688980957
transform 1 0 27968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S0
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S1
timestamp 1688980957
transform -1 0 31096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__S0
timestamp 1688980957
transform 1 0 35236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__S1
timestamp 1688980957
transform 1 0 34868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__S
timestamp 1688980957
transform 1 0 37904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S0
timestamp 1688980957
transform 1 0 31924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S1
timestamp 1688980957
transform 1 0 32200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__S0
timestamp 1688980957
transform 1 0 31832 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__S1
timestamp 1688980957
transform 1 0 32016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__S
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1688980957
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S0
timestamp 1688980957
transform 1 0 38548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S1
timestamp 1688980957
transform 1 0 38272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__S0
timestamp 1688980957
transform 1 0 36432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__S1
timestamp 1688980957
transform 1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__S
timestamp 1688980957
transform 1 0 41308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1688980957
transform 1 0 38640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S0
timestamp 1688980957
transform 1 0 32292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S1
timestamp 1688980957
transform 1 0 32568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__S0
timestamp 1688980957
transform -1 0 32660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__S1
timestamp 1688980957
transform -1 0 32476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__S
timestamp 1688980957
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1688980957
transform 1 0 41860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S0
timestamp 1688980957
transform 1 0 37076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S1
timestamp 1688980957
transform 1 0 36708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__S0
timestamp 1688980957
transform -1 0 38548 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__S1
timestamp 1688980957
transform -1 0 37168 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__S
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1688980957
transform 1 0 43332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S0
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S1
timestamp 1688980957
transform 1 0 38180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__S0
timestamp 1688980957
transform 1 0 38272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__S1
timestamp 1688980957
transform 1 0 37812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__S
timestamp 1688980957
transform 1 0 39100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1688980957
transform 1 0 44804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__S0
timestamp 1688980957
transform -1 0 44344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__S1
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__S0
timestamp 1688980957
transform 1 0 40480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__S1
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__S
timestamp 1688980957
transform 1 0 45264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1688980957
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__S0
timestamp 1688980957
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__S1
timestamp 1688980957
transform 1 0 41032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__S0
timestamp 1688980957
transform 1 0 42044 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__S1
timestamp 1688980957
transform 1 0 41400 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__S
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1688980957
transform 1 0 48300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__S0
timestamp 1688980957
transform 1 0 45540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__S1
timestamp 1688980957
transform 1 0 45172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__S0
timestamp 1688980957
transform 1 0 46000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__S1
timestamp 1688980957
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__S
timestamp 1688980957
transform 1 0 44160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1688980957
transform 1 0 47932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S0
timestamp 1688980957
transform 1 0 47380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S1
timestamp 1688980957
transform 1 0 46736 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__S0
timestamp 1688980957
transform 1 0 46644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__S1
timestamp 1688980957
transform 1 0 47012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__S
timestamp 1688980957
transform 1 0 47748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1688980957
transform 1 0 48116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S0
timestamp 1688980957
transform 1 0 47196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S1
timestamp 1688980957
transform 1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__S0
timestamp 1688980957
transform 1 0 47748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__S1
timestamp 1688980957
transform 1 0 46828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__S
timestamp 1688980957
transform -1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1688980957
transform 1 0 52348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__S0
timestamp 1688980957
transform 1 0 48576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__S1
timestamp 1688980957
transform 1 0 48392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__S0
timestamp 1688980957
transform 1 0 48392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__S1
timestamp 1688980957
transform 1 0 48760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__S
timestamp 1688980957
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1688980957
transform 1 0 51980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S0
timestamp 1688980957
transform 1 0 49680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S1
timestamp 1688980957
transform 1 0 49036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__S0
timestamp 1688980957
transform 1 0 48852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__S1
timestamp 1688980957
transform 1 0 48852 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__S
timestamp 1688980957
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1688980957
transform 1 0 51244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S0
timestamp 1688980957
transform 1 0 53820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S1
timestamp 1688980957
transform 1 0 54924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__S0
timestamp 1688980957
transform 1 0 54096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__S1
timestamp 1688980957
transform 1 0 54464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__S
timestamp 1688980957
transform 1 0 55108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1688980957
transform 1 0 53452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S0
timestamp 1688980957
transform 1 0 55844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S1
timestamp 1688980957
transform 1 0 52348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__S0
timestamp 1688980957
transform 1 0 55476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__S1
timestamp 1688980957
transform 1 0 54832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__S
timestamp 1688980957
transform 1 0 51612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1688980957
transform -1 0 55292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S0
timestamp 1688980957
transform 1 0 55200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S1
timestamp 1688980957
transform 1 0 55568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__S0
timestamp 1688980957
transform 1 0 55476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__S1
timestamp 1688980957
transform 1 0 55752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S
timestamp 1688980957
transform -1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1688980957
transform 1 0 51980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S0
timestamp 1688980957
transform 1 0 54004 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S1
timestamp 1688980957
transform 1 0 54004 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S0
timestamp 1688980957
transform 1 0 54280 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S1
timestamp 1688980957
transform -1 0 53912 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__S
timestamp 1688980957
transform 1 0 55016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1688980957
transform 1 0 50876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__S
timestamp 1688980957
transform 1 0 27324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__S
timestamp 1688980957
transform 1 0 34592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__S
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__S
timestamp 1688980957
transform 1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__S
timestamp 1688980957
transform 1 0 36800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__S
timestamp 1688980957
transform -1 0 33304 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__S
timestamp 1688980957
transform 1 0 39468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__S
timestamp 1688980957
transform 1 0 37812 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__S
timestamp 1688980957
transform 1 0 40020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1688980957
transform 1 0 42780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__S
timestamp 1688980957
transform -1 0 45724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1688980957
transform 1 0 51980 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__S
timestamp 1688980957
transform -1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1688980957
transform 1 0 50324 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__S
timestamp 1688980957
transform 1 0 48668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__S
timestamp 1688980957
transform 1 0 55568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1688980957
transform -1 0 58512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__S
timestamp 1688980957
transform 1 0 56212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1688980957
transform 1 0 55016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__S
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__S
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__S
timestamp 1688980957
transform 1 0 12696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__S
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1688980957
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__S
timestamp 1688980957
transform 1 0 17112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__S
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1688980957
transform -1 0 21620 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__S
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__S
timestamp 1688980957
transform -1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1688980957
transform 1 0 25852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__S
timestamp 1688980957
transform 1 0 33948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1688980957
transform 1 0 28244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1688980957
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1688980957
transform 1 0 40020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__S
timestamp 1688980957
transform 1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1688980957
transform 1 0 38180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1688980957
transform 1 0 44620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1688980957
transform 1 0 45264 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__S
timestamp 1688980957
transform 1 0 44528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1688980957
transform 1 0 48944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__S
timestamp 1688980957
transform 1 0 48944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1688980957
transform 1 0 50508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__S
timestamp 1688980957
transform 1 0 49956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1688980957
transform 1 0 57500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__S
timestamp 1688980957
transform -1 0 58236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1688980957
transform 1 0 56304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__S
timestamp 1688980957
transform -1 0 56672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__S
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__S
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1688980957
transform -1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__S
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1688980957
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__S
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__S
timestamp 1688980957
transform 1 0 16928 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__S
timestamp 1688980957
transform 1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1688980957
transform 1 0 21160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__S
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__S
timestamp 1688980957
transform 1 0 23368 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__S
timestamp 1688980957
transform 1 0 27968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1688980957
transform 1 0 29348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__S
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1688980957
transform -1 0 30360 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__S
timestamp 1688980957
transform 1 0 35604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1688980957
transform 1 0 36616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__S
timestamp 1688980957
transform 1 0 40848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1688980957
transform 1 0 42412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1688980957
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__S
timestamp 1688980957
transform 1 0 47748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1688980957
transform -1 0 47196 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__S
timestamp 1688980957
transform 1 0 47380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__S
timestamp 1688980957
transform 1 0 48576 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__S
timestamp 1688980957
transform 1 0 52716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__S
timestamp 1688980957
transform 1 0 51612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__S
timestamp 1688980957
transform 1 0 54096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__S
timestamp 1688980957
transform -1 0 52164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1688980957
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A_N
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A_N
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A_N
timestamp 1688980957
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B
timestamp 1688980957
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__S
timestamp 1688980957
transform 1 0 4600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__S
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__S
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__S
timestamp 1688980957
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__S
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__S
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__S
timestamp 1688980957
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__S
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S
timestamp 1688980957
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__S
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__S
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__S
timestamp 1688980957
transform 1 0 28704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__S
timestamp 1688980957
transform -1 0 26772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S
timestamp 1688980957
transform 1 0 38180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__S
timestamp 1688980957
transform -1 0 31648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__S
timestamp 1688980957
transform -1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S
timestamp 1688980957
transform 1 0 36800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S
timestamp 1688980957
transform 1 0 39008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__S
timestamp 1688980957
transform 1 0 41584 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__S
timestamp 1688980957
transform 1 0 41676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S
timestamp 1688980957
transform 1 0 46368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S
timestamp 1688980957
transform 1 0 45356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__S
timestamp 1688980957
transform 1 0 46920 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__S
timestamp 1688980957
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S
timestamp 1688980957
transform -1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S
timestamp 1688980957
transform 1 0 51704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__S
timestamp 1688980957
transform 1 0 54004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__S
timestamp 1688980957
transform -1 0 52256 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S
timestamp 1688980957
transform 1 0 4508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__S
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__S
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S
timestamp 1688980957
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S
timestamp 1688980957
transform 1 0 10580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__S
timestamp 1688980957
transform -1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__S
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__S
timestamp 1688980957
transform 1 0 18768 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__S
timestamp 1688980957
transform 1 0 21896 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S
timestamp 1688980957
transform 1 0 20240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S
timestamp 1688980957
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__S
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__S
timestamp 1688980957
transform -1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S
timestamp 1688980957
transform 1 0 31188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S
timestamp 1688980957
transform 1 0 29900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__S
timestamp 1688980957
transform 1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__S
timestamp 1688980957
transform 1 0 29532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S
timestamp 1688980957
transform -1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S
timestamp 1688980957
transform 1 0 37076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__S
timestamp 1688980957
transform 1 0 39652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__S
timestamp 1688980957
transform 1 0 42228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S
timestamp 1688980957
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S
timestamp 1688980957
transform 1 0 48484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__S
timestamp 1688980957
transform -1 0 45908 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1688980957
transform 1 0 47380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S
timestamp 1688980957
transform 1 0 46920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S
timestamp 1688980957
transform 1 0 53084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1688980957
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__S
timestamp 1688980957
transform -1 0 52624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S
timestamp 1688980957
transform -1 0 54096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__S
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__S
timestamp 1688980957
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S
timestamp 1688980957
transform -1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__S
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__S
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S
timestamp 1688980957
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__S
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1688980957
transform 1 0 25944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__S
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S
timestamp 1688980957
transform -1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S
timestamp 1688980957
transform 1 0 35696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__S
timestamp 1688980957
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S
timestamp 1688980957
transform 1 0 35236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S
timestamp 1688980957
transform -1 0 39100 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S
timestamp 1688980957
transform 1 0 40480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1688980957
transform 1 0 44160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S
timestamp 1688980957
transform 1 0 41676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S
timestamp 1688980957
transform 1 0 43332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S
timestamp 1688980957
transform 1 0 48760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__S
timestamp 1688980957
transform 1 0 49588 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S
timestamp 1688980957
transform 1 0 51980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S
timestamp 1688980957
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__S
timestamp 1688980957
transform 1 0 57408 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp 1688980957
transform 1 0 55476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S
timestamp 1688980957
transform -1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S
timestamp 1688980957
transform 1 0 55016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp 1688980957
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp 1688980957
transform -1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp 1688980957
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp 1688980957
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__S
timestamp 1688980957
transform 1 0 19872 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__S
timestamp 1688980957
transform -1 0 22172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S
timestamp 1688980957
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp 1688980957
transform 1 0 25208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__S
timestamp 1688980957
transform 1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__S
timestamp 1688980957
transform 1 0 27324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S
timestamp 1688980957
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S
timestamp 1688980957
transform -1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp 1688980957
transform 1 0 35236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp 1688980957
transform 1 0 40112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S
timestamp 1688980957
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S
timestamp 1688980957
transform -1 0 39744 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1688980957
transform 1 0 40020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp 1688980957
transform 1 0 44436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S
timestamp 1688980957
transform 1 0 43700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S
timestamp 1688980957
transform 1 0 46368 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1688980957
transform 1 0 50324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp 1688980957
transform 1 0 50140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S
timestamp 1688980957
transform 1 0 50508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp 1688980957
transform 1 0 50140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__S
timestamp 1688980957
transform 1 0 56304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__S
timestamp 1688980957
transform -1 0 57408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S
timestamp 1688980957
transform 1 0 56396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__S
timestamp 1688980957
transform -1 0 56028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1688980957
transform 1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1688980957
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1688980957
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__S
timestamp 1688980957
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp 1688980957
transform -1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S
timestamp 1688980957
transform 1 0 5520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S
timestamp 1688980957
transform 1 0 13064 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp 1688980957
transform -1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S
timestamp 1688980957
transform 1 0 16744 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__S
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp 1688980957
transform 1 0 18308 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__S
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp 1688980957
transform 1 0 23368 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S
timestamp 1688980957
transform 1 0 30452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S
timestamp 1688980957
transform -1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__S
timestamp 1688980957
transform 1 0 31188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__S
timestamp 1688980957
transform 1 0 41032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__S
timestamp 1688980957
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S
timestamp 1688980957
transform 1 0 36616 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp 1688980957
transform 1 0 35696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__S
timestamp 1688980957
transform 1 0 44896 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S
timestamp 1688980957
transform -1 0 42320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S
timestamp 1688980957
transform 1 0 42228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__S
timestamp 1688980957
transform 1 0 46000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__S
timestamp 1688980957
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S
timestamp 1688980957
transform 1 0 46552 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S
timestamp 1688980957
transform 1 0 48300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__S
timestamp 1688980957
transform 1 0 52900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__S
timestamp 1688980957
transform 1 0 52900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S
timestamp 1688980957
transform 1 0 52992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__S
timestamp 1688980957
transform -1 0 53912 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__S
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__S
timestamp 1688980957
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__S
timestamp 1688980957
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__S
timestamp 1688980957
transform 1 0 12972 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__S
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__S
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__S
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__S
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__S
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__S
timestamp 1688980957
transform 1 0 25760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__S
timestamp 1688980957
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__S
timestamp 1688980957
transform 1 0 28704 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__CLK
timestamp 1688980957
transform 1 0 29256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__CLK
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__CLK
timestamp 1688980957
transform 1 0 33856 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__CLK
timestamp 1688980957
transform 1 0 32752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__CLK
timestamp 1688980957
transform 1 0 38640 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__CLK
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__CLK
timestamp 1688980957
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__CLK
timestamp 1688980957
transform 1 0 41308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__CLK
timestamp 1688980957
transform 1 0 44528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__CLK
timestamp 1688980957
transform 1 0 44620 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__CLK
timestamp 1688980957
transform 1 0 46000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__CLK
timestamp 1688980957
transform -1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__CLK
timestamp 1688980957
transform 1 0 51612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__CLK
timestamp 1688980957
transform 1 0 55936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__CLK
timestamp 1688980957
transform 1 0 55660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__CLK
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__CLK
timestamp 1688980957
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__CLK
timestamp 1688980957
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__CLK
timestamp 1688980957
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__CLK
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__CLK
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__CLK
timestamp 1688980957
transform 1 0 27876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__CLK
timestamp 1688980957
transform 1 0 26588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__CLK
timestamp 1688980957
transform -1 0 26588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__CLK
timestamp 1688980957
transform 1 0 31740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__CLK
timestamp 1688980957
transform 1 0 38732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__CLK
timestamp 1688980957
transform 1 0 33764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__CLK
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__CLK
timestamp 1688980957
transform 1 0 39376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__CLK
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__CLK
timestamp 1688980957
transform 1 0 44528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__CLK
timestamp 1688980957
transform -1 0 45080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__CLK
timestamp 1688980957
transform 1 0 51060 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__CLK
timestamp 1688980957
transform 1 0 52348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__CLK
timestamp 1688980957
transform 1 0 56120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__CLK
timestamp 1688980957
transform 1 0 56120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__CLK
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__CLK
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__CLK
timestamp 1688980957
transform -1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__CLK
timestamp 1688980957
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__CLK
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__CLK
timestamp 1688980957
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__CLK
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__CLK
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__CLK
timestamp 1688980957
transform 1 0 31556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__CLK
timestamp 1688980957
transform -1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__CLK
timestamp 1688980957
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__CLK
timestamp 1688980957
transform -1 0 32292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__CLK
timestamp 1688980957
transform 1 0 37720 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__CLK
timestamp 1688980957
transform 1 0 38272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__CLK
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__CLK
timestamp 1688980957
transform 1 0 40940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__CLK
timestamp 1688980957
transform 1 0 42596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__CLK
timestamp 1688980957
transform 1 0 45264 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__CLK
timestamp 1688980957
transform 1 0 45172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__CLK
timestamp 1688980957
transform 1 0 48576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__CLK
timestamp 1688980957
transform 1 0 46644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__CLK
timestamp 1688980957
transform 1 0 52808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__CLK
timestamp 1688980957
transform 1 0 52624 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__CLK
timestamp 1688980957
transform 1 0 51336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__CLK
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__CLK
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__CLK
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__CLK
timestamp 1688980957
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__CLK
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__CLK
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__CLK
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__CLK
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__CLK
timestamp 1688980957
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__CLK
timestamp 1688980957
transform -1 0 27876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__CLK
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__CLK
timestamp 1688980957
transform 1 0 31280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__CLK
timestamp 1688980957
transform 1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__CLK
timestamp 1688980957
transform 1 0 31832 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__CLK
timestamp 1688980957
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__CLK
timestamp 1688980957
transform 1 0 37352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__CLK
timestamp 1688980957
transform 1 0 40112 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__CLK
timestamp 1688980957
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__CLK
timestamp 1688980957
transform 1 0 48668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__CLK
timestamp 1688980957
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__CLK
timestamp 1688980957
transform 1 0 49496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__CLK
timestamp 1688980957
transform 1 0 45908 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__CLK
timestamp 1688980957
transform 1 0 52900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__CLK
timestamp 1688980957
transform 1 0 53084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__CLK
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__CLK
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__CLK
timestamp 1688980957
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__CLK
timestamp 1688980957
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__CLK
timestamp 1688980957
transform -1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__CLK
timestamp 1688980957
transform 1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__CLK
timestamp 1688980957
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__CLK
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__CLK
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__CLK
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__CLK
timestamp 1688980957
transform 1 0 32108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__CLK
timestamp 1688980957
transform 1 0 38548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__CLK
timestamp 1688980957
transform 1 0 41216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__CLK
timestamp 1688980957
transform 1 0 42596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__CLK
timestamp 1688980957
transform 1 0 44436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__CLK
timestamp 1688980957
transform 1 0 45172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__CLK
timestamp 1688980957
transform 1 0 45724 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__CLK
timestamp 1688980957
transform 1 0 49312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__CLK
timestamp 1688980957
transform 1 0 46276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__CLK
timestamp 1688980957
transform 1 0 52440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__CLK
timestamp 1688980957
transform 1 0 52900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__CLK
timestamp 1688980957
transform 1 0 51796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__CLK
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__CLK
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__CLK
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__CLK
timestamp 1688980957
transform 1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__CLK
timestamp 1688980957
transform 1 0 27140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__CLK
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__CLK
timestamp 1688980957
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__CLK
timestamp 1688980957
transform 1 0 29808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__CLK
timestamp 1688980957
transform 1 0 35236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__CLK
timestamp 1688980957
transform 1 0 34224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__CLK
timestamp 1688980957
transform 1 0 40480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__CLK
timestamp 1688980957
transform -1 0 35788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__CLK
timestamp 1688980957
transform 1 0 39652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__CLK
timestamp 1688980957
transform 1 0 39652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__CLK
timestamp 1688980957
transform 1 0 42044 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__CLK
timestamp 1688980957
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__CLK
timestamp 1688980957
transform -1 0 44620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__CLK
timestamp 1688980957
transform 1 0 48392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__CLK
timestamp 1688980957
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__CLK
timestamp 1688980957
transform 1 0 52348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__CLK
timestamp 1688980957
transform 1 0 50600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__CLK
timestamp 1688980957
transform 1 0 55936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__CLK
timestamp 1688980957
transform 1 0 55568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__CLK
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__CLK
timestamp 1688980957
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__CLK
timestamp 1688980957
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__CLK
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__CLK
timestamp 1688980957
transform 1 0 21344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__CLK
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__CLK
timestamp 1688980957
transform 1 0 25024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__CLK
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__CLK
timestamp 1688980957
transform 1 0 34132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__CLK
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__CLK
timestamp 1688980957
transform -1 0 40940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__CLK
timestamp 1688980957
transform -1 0 34500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__CLK
timestamp 1688980957
transform 1 0 41308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__CLK
timestamp 1688980957
transform 1 0 40388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__CLK
timestamp 1688980957
transform 1 0 43884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__CLK
timestamp 1688980957
transform 1 0 45172 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__CLK
timestamp 1688980957
transform 1 0 46736 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__CLK
timestamp 1688980957
transform -1 0 50692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__CLK
timestamp 1688980957
transform 1 0 49772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__CLK
timestamp 1688980957
transform -1 0 51796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__CLK
timestamp 1688980957
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__CLK
timestamp 1688980957
transform 1 0 56120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__CLK
timestamp 1688980957
transform 1 0 56120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__CLK
timestamp 1688980957
transform 1 0 55016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__CLK
timestamp 1688980957
transform -1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1688980957
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1688980957
transform 1 0 23460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__CLK
timestamp 1688980957
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1688980957
transform 1 0 29900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1688980957
transform 1 0 27508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1688980957
transform 1 0 31556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1688980957
transform 1 0 42044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1688980957
transform 1 0 31740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1688980957
transform 1 0 35512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1688980957
transform 1 0 37444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1688980957
transform -1 0 41308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1688980957
transform 1 0 40112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1688980957
transform 1 0 45632 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1688980957
transform 1 0 44620 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__CLK
timestamp 1688980957
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1688980957
transform 1 0 52532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__CLK
timestamp 1688980957
transform 1 0 53452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__CLK
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__CLK
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1688980957
transform 1 0 19872 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1688980957
transform 1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1688980957
transform 1 0 27876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__CLK
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1688980957
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1688980957
transform 1 0 34132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1688980957
transform 1 0 44528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1688980957
transform 1 0 51060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1688980957
transform 1 0 43608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1688980957
transform -1 0 54188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1688980957
transform 1 0 44068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1688980957
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout1_A
timestamp 1688980957
transform -1 0 38824 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout2_A
timestamp 1688980957
transform -1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform -1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform 1 0 28336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform -1 0 35052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform -1 0 34132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1688980957
transform -1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 1688980957
transform 1 0 28612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 1688980957
transform 1 0 33120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 1688980957
transform -1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 1688980957
transform -1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 1688980957
transform -1 0 31832 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp 1688980957
transform 1 0 46184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 1688980957
transform 1 0 31004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1688980957
transform -1 0 7544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1688980957
transform -1 0 43884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp 1688980957
transform 1 0 30452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold558_A
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 20056 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 39008 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1688980957
transform -1 0 8188 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1688980957
transform -1 0 21252 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1688980957
transform -1 0 33948 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1688980957
transform -1 0 45908 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1688980957
transform 1 0 50600 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1688980957
transform 1 0 43240 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1688980957
transform 1 0 53176 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1688980957
transform 1 0 26864 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1688980957
transform -1 0 13432 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1688980957
transform 1 0 9844 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout2
timestamp 1688980957
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout102 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout103
timestamp 1688980957
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout104
timestamp 1688980957
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout105
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout106
timestamp 1688980957
transform 1 0 33580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout107
timestamp 1688980957
transform -1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout108
timestamp 1688980957
transform 1 0 32660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout109
timestamp 1688980957
transform -1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout110
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout111
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout112
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout113
timestamp 1688980957
transform 1 0 13340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout114
timestamp 1688980957
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout115
timestamp 1688980957
transform -1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout116
timestamp 1688980957
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout117
timestamp 1688980957
transform -1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout119 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout120
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout121 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout122
timestamp 1688980957
transform -1 0 10212 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout123
timestamp 1688980957
transform -1 0 46000 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout124
timestamp 1688980957
transform 1 0 31188 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout125 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout126
timestamp 1688980957
transform 1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout127
timestamp 1688980957
transform -1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout128
timestamp 1688980957
transform 1 0 43884 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout129
timestamp 1688980957
transform 1 0 30636 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout130
timestamp 1688980957
transform -1 0 8832 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_116 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_150
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_318
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_340
timestamp 1688980957
transform 1 0 32384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_362
timestamp 1688980957
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_577
timestamp 1688980957
transform 1 0 54188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_587
timestamp 1688980957
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_614
timestamp 1688980957
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_25
timestamp 1688980957
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_30
timestamp 1688980957
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_95
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_236
timestamp 1688980957
transform 1 0 22816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_321
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_375
timestamp 1688980957
transform 1 0 35604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_381
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_411
timestamp 1688980957
transform 1 0 38916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_471
timestamp 1688980957
transform 1 0 44436 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_612
timestamp 1688980957
transform 1 0 57408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_62
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1688980957
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_102
timestamp 1688980957
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_114
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_131
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_161
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_236
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_275
timestamp 1688980957
transform 1 0 26404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_354
timestamp 1688980957
transform 1 0 33672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1688980957
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_459
timestamp 1688980957
transform 1 0 43332 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1688980957
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_541
timestamp 1688980957
transform 1 0 50876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_550
timestamp 1688980957
transform 1 0 51704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_586
timestamp 1688980957
transform 1 0 55016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_589
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_80
timestamp 1688980957
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_96
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_100
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_104
timestamp 1688980957
transform 1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_108
timestamp 1688980957
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_160
timestamp 1688980957
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_164
timestamp 1688980957
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_186
timestamp 1688980957
transform 1 0 18216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_243
timestamp 1688980957
transform 1 0 23460 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_291
timestamp 1688980957
transform 1 0 27876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_311
timestamp 1688980957
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_360
timestamp 1688980957
transform 1 0 34224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_404
timestamp 1688980957
transform 1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_432
timestamp 1688980957
transform 1 0 40848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_466
timestamp 1688980957
transform 1 0 43976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_498
timestamp 1688980957
transform 1 0 46920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_502
timestamp 1688980957
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_520
timestamp 1688980957
transform 1 0 48944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_546
timestamp 1688980957
transform 1 0 51336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_570
timestamp 1688980957
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_8
timestamp 1688980957
transform 1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_51
timestamp 1688980957
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_55
timestamp 1688980957
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_62
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_73
timestamp 1688980957
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_90
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_94
timestamp 1688980957
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_150
timestamp 1688980957
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_158
timestamp 1688980957
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_179
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_222
timestamp 1688980957
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_274
timestamp 1688980957
transform 1 0 26312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_281
timestamp 1688980957
transform 1 0 26956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_286
timestamp 1688980957
transform 1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_290
timestamp 1688980957
transform 1 0 27784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_302
timestamp 1688980957
transform 1 0 28888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_375
timestamp 1688980957
transform 1 0 35604 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_398
timestamp 1688980957
transform 1 0 37720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_402
timestamp 1688980957
transform 1 0 38088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_406
timestamp 1688980957
transform 1 0 38456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_474
timestamp 1688980957
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_507
timestamp 1688980957
transform 1 0 47748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_511
timestamp 1688980957
transform 1 0 48116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_515
timestamp 1688980957
transform 1 0 48484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_519
timestamp 1688980957
transform 1 0 48852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_523
timestamp 1688980957
transform 1 0 49220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_527
timestamp 1688980957
transform 1 0 49588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_549
timestamp 1688980957
transform 1 0 51612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_578
timestamp 1688980957
transform 1 0 54280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_623
timestamp 1688980957
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_13
timestamp 1688980957
transform 1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_17
timestamp 1688980957
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_30
timestamp 1688980957
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_34
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_50
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_65
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_122
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_151
timestamp 1688980957
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_156
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_160
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_186
timestamp 1688980957
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_203
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_211
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_215
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_259
timestamp 1688980957
transform 1 0 24932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_285
timestamp 1688980957
transform 1 0 27324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_289
timestamp 1688980957
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_297
timestamp 1688980957
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_301
timestamp 1688980957
transform 1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_325
timestamp 1688980957
transform 1 0 31004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_333
timestamp 1688980957
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_365
timestamp 1688980957
transform 1 0 34684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_369
timestamp 1688980957
transform 1 0 35052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_389
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_402
timestamp 1688980957
transform 1 0 38088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_435
timestamp 1688980957
transform 1 0 41124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_439
timestamp 1688980957
transform 1 0 41492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_443
timestamp 1688980957
transform 1 0 41860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_458
timestamp 1688980957
transform 1 0 43240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_462
timestamp 1688980957
transform 1 0 43608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_466
timestamp 1688980957
transform 1 0 43976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_470
timestamp 1688980957
transform 1 0 44344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_474
timestamp 1688980957
transform 1 0 44712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_478
timestamp 1688980957
transform 1 0 45080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_482
timestamp 1688980957
transform 1 0 45448 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_502
timestamp 1688980957
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_513
timestamp 1688980957
transform 1 0 48300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_517
timestamp 1688980957
transform 1 0 48668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_535
timestamp 1688980957
transform 1 0 50324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_551
timestamp 1688980957
transform 1 0 51796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_555
timestamp 1688980957
transform 1 0 52164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1688980957
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_569
timestamp 1688980957
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_573
timestamp 1688980957
transform 1 0 53820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_577
timestamp 1688980957
transform 1 0 54188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_582
timestamp 1688980957
transform 1 0 54648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_601
timestamp 1688980957
transform 1 0 56396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1688980957
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_7
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_101
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_154
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_159
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_163
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_169
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_173
timestamp 1688980957
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_201
timestamp 1688980957
transform 1 0 19596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_223
timestamp 1688980957
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_228
timestamp 1688980957
transform 1 0 22080 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_240
timestamp 1688980957
transform 1 0 23184 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_249
timestamp 1688980957
transform 1 0 24012 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_283
timestamp 1688980957
transform 1 0 27140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_287
timestamp 1688980957
transform 1 0 27508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_291
timestamp 1688980957
transform 1 0 27876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_295
timestamp 1688980957
transform 1 0 28244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_362
timestamp 1688980957
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_373
timestamp 1688980957
transform 1 0 35420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_403
timestamp 1688980957
transform 1 0 38180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_407
timestamp 1688980957
transform 1 0 38548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_441
timestamp 1688980957
transform 1 0 41676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_465
timestamp 1688980957
transform 1 0 43884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_473
timestamp 1688980957
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_586
timestamp 1688980957
transform 1 0 55016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_624
timestamp 1688980957
transform 1 0 58512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_11
timestamp 1688980957
transform 1 0 2116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_14
timestamp 1688980957
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_34
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_92
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_122
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_218
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_233
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_251
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_255
timestamp 1688980957
transform 1 0 24564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1688980957
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_289
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_330
timestamp 1688980957
transform 1 0 31464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_365
timestamp 1688980957
transform 1 0 34684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_369
timestamp 1688980957
transform 1 0 35052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_386
timestamp 1688980957
transform 1 0 36616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_390
timestamp 1688980957
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_401
timestamp 1688980957
transform 1 0 37996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_409
timestamp 1688980957
transform 1 0 38732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_434
timestamp 1688980957
transform 1 0 41032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_438
timestamp 1688980957
transform 1 0 41400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_477
timestamp 1688980957
transform 1 0 44988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_502
timestamp 1688980957
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_505
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_509
timestamp 1688980957
transform 1 0 47932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_513
timestamp 1688980957
transform 1 0 48300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_516
timestamp 1688980957
transform 1 0 48576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_545
timestamp 1688980957
transform 1 0 51244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_577
timestamp 1688980957
transform 1 0 54188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_599
timestamp 1688980957
transform 1 0 56212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_43
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_50
timestamp 1688980957
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_54
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_58
timestamp 1688980957
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_78
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_89
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_116
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_157
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_161
timestamp 1688980957
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_218
timestamp 1688980957
transform 1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_222
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_318
timestamp 1688980957
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_335
timestamp 1688980957
transform 1 0 31924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1688980957
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_369
timestamp 1688980957
transform 1 0 35052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_398
timestamp 1688980957
transform 1 0 37720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_402
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_406
timestamp 1688980957
transform 1 0 38456 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_410
timestamp 1688980957
transform 1 0 38824 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_459
timestamp 1688980957
transform 1 0 43332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_463
timestamp 1688980957
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_467
timestamp 1688980957
transform 1 0 44068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_471
timestamp 1688980957
transform 1 0 44436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_493
timestamp 1688980957
transform 1 0 46460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_497
timestamp 1688980957
transform 1 0 46828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_501
timestamp 1688980957
transform 1 0 47196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_505
timestamp 1688980957
transform 1 0 47564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_509
timestamp 1688980957
transform 1 0 47932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_513
timestamp 1688980957
transform 1 0 48300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_519
timestamp 1688980957
transform 1 0 48852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_522
timestamp 1688980957
transform 1 0 49128 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_530
timestamp 1688980957
transform 1 0 49864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_537
timestamp 1688980957
transform 1 0 50508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_543
timestamp 1688980957
transform 1 0 51060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_547
timestamp 1688980957
transform 1 0 51428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_585
timestamp 1688980957
transform 1 0 54924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_602
timestamp 1688980957
transform 1 0 56488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_621
timestamp 1688980957
transform 1 0 58236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_46
timestamp 1688980957
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_61
timestamp 1688980957
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_97
timestamp 1688980957
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_101
timestamp 1688980957
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_173
timestamp 1688980957
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_180
timestamp 1688980957
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_184
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_195
timestamp 1688980957
transform 1 0 19044 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_215
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_245
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_254
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_258
timestamp 1688980957
transform 1 0 24840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_289
timestamp 1688980957
transform 1 0 27692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_306
timestamp 1688980957
transform 1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_314
timestamp 1688980957
transform 1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_333
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_341
timestamp 1688980957
transform 1 0 32476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_355
timestamp 1688980957
transform 1 0 33764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_363
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_382
timestamp 1688980957
transform 1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_386
timestamp 1688980957
transform 1 0 36616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_390
timestamp 1688980957
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_406
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_410
timestamp 1688980957
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_414
timestamp 1688980957
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_418
timestamp 1688980957
transform 1 0 39560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_421
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_425
timestamp 1688980957
transform 1 0 40204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_430
timestamp 1688980957
transform 1 0 40664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_443
timestamp 1688980957
transform 1 0 41860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_466
timestamp 1688980957
transform 1 0 43976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_470
timestamp 1688980957
transform 1 0 44344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_474
timestamp 1688980957
transform 1 0 44712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_478
timestamp 1688980957
transform 1 0 45080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_482
timestamp 1688980957
transform 1 0 45448 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_486
timestamp 1688980957
transform 1 0 45816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_490
timestamp 1688980957
transform 1 0 46184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_494
timestamp 1688980957
transform 1 0 46552 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_498
timestamp 1688980957
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_513
timestamp 1688980957
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_532 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 50048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_544
timestamp 1688980957
transform 1 0 51152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_548
timestamp 1688980957
transform 1 0 51520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_551
timestamp 1688980957
transform 1 0 51796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_555
timestamp 1688980957
transform 1 0 52164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_561
timestamp 1688980957
transform 1 0 52716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_565
timestamp 1688980957
transform 1 0 53084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_571
timestamp 1688980957
transform 1 0 53636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_575
timestamp 1688980957
transform 1 0 54004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_584
timestamp 1688980957
transform 1 0 54832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_589
timestamp 1688980957
transform 1 0 55292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_593
timestamp 1688980957
transform 1 0 55660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_597
timestamp 1688980957
transform 1 0 56028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_608
timestamp 1688980957
transform 1 0 57040 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_32
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_39
timestamp 1688980957
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_43
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_49
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_68
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_95
timestamp 1688980957
transform 1 0 9844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_99
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_104
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_116
timestamp 1688980957
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_134
timestamp 1688980957
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_169
timestamp 1688980957
transform 1 0 16652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_184
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_192
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_234
timestamp 1688980957
transform 1 0 22632 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_278
timestamp 1688980957
transform 1 0 26680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_330
timestamp 1688980957
transform 1 0 31464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_334
timestamp 1688980957
transform 1 0 31832 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 1688980957
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_376
timestamp 1688980957
transform 1 0 35696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_417
timestamp 1688980957
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_425
timestamp 1688980957
transform 1 0 40204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_459
timestamp 1688980957
transform 1 0 43332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_463
timestamp 1688980957
transform 1 0 43700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_485
timestamp 1688980957
transform 1 0 45724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_510
timestamp 1688980957
transform 1 0 48024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_527
timestamp 1688980957
transform 1 0 49588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_549
timestamp 1688980957
transform 1 0 51612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_555
timestamp 1688980957
transform 1 0 52164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_583
timestamp 1688980957
transform 1 0 54740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1688980957
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_598
timestamp 1688980957
transform 1 0 56120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_624
timestamp 1688980957
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_22
timestamp 1688980957
transform 1 0 3128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_36
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_76
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_99
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_103
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_109
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 1688980957
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_207
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_219
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_248
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_259
timestamp 1688980957
transform 1 0 24932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_270
timestamp 1688980957
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_310
timestamp 1688980957
transform 1 0 29624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_353
timestamp 1688980957
transform 1 0 33580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_357
timestamp 1688980957
transform 1 0 33948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_422
timestamp 1688980957
transform 1 0 39928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_426
timestamp 1688980957
transform 1 0 40296 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_430
timestamp 1688980957
transform 1 0 40664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_484
timestamp 1688980957
transform 1 0 45632 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_502
timestamp 1688980957
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_598
timestamp 1688980957
transform 1 0 56120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_46
timestamp 1688980957
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_50
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_62
timestamp 1688980957
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_71
timestamp 1688980957
transform 1 0 7636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_115
timestamp 1688980957
transform 1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_169
timestamp 1688980957
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_225
timestamp 1688980957
transform 1 0 21804 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_261
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_279
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_285
timestamp 1688980957
transform 1 0 27324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_302
timestamp 1688980957
transform 1 0 28888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_353
timestamp 1688980957
transform 1 0 33580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_361
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_395
timestamp 1688980957
transform 1 0 37444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_429
timestamp 1688980957
transform 1 0 40572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_437
timestamp 1688980957
transform 1 0 41308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_449
timestamp 1688980957
transform 1 0 42412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_461
timestamp 1688980957
transform 1 0 43516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_465
timestamp 1688980957
transform 1 0 43884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_474
timestamp 1688980957
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_481
timestamp 1688980957
transform 1 0 45356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_485
timestamp 1688980957
transform 1 0 45724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_493
timestamp 1688980957
transform 1 0 46460 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_511
timestamp 1688980957
transform 1 0 48116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_515
timestamp 1688980957
transform 1 0 48484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_526
timestamp 1688980957
transform 1 0 49496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_530
timestamp 1688980957
transform 1 0 49864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_542
timestamp 1688980957
transform 1 0 50968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_550
timestamp 1688980957
transform 1 0 51704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_582
timestamp 1688980957
transform 1 0 54648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_586
timestamp 1688980957
transform 1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_597
timestamp 1688980957
transform 1 0 56028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_620
timestamp 1688980957
transform 1 0 58144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_624
timestamp 1688980957
transform 1 0 58512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_22
timestamp 1688980957
transform 1 0 3128 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_28
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_36
timestamp 1688980957
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_62
timestamp 1688980957
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_66
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_78
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_150
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_186
timestamp 1688980957
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_190
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_198
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_234
timestamp 1688980957
transform 1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_257
timestamp 1688980957
transform 1 0 24748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_275
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_285
timestamp 1688980957
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_311
timestamp 1688980957
transform 1 0 29716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_315
timestamp 1688980957
transform 1 0 30084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_330
timestamp 1688980957
transform 1 0 31464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_355
timestamp 1688980957
transform 1 0 33764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_359
timestamp 1688980957
transform 1 0 34132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_363
timestamp 1688980957
transform 1 0 34500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_379
timestamp 1688980957
transform 1 0 35972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_401
timestamp 1688980957
transform 1 0 37996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_436
timestamp 1688980957
transform 1 0 41216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_458
timestamp 1688980957
transform 1 0 43240 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_462
timestamp 1688980957
transform 1 0 43608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_474
timestamp 1688980957
transform 1 0 44712 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_486
timestamp 1688980957
transform 1 0 45816 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_490
timestamp 1688980957
transform 1 0 46184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_500
timestamp 1688980957
transform 1 0 47104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_515
timestamp 1688980957
transform 1 0 48484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_519
timestamp 1688980957
transform 1 0 48852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_523
timestamp 1688980957
transform 1 0 49220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_533
timestamp 1688980957
transform 1 0 50140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_537
timestamp 1688980957
transform 1 0 50508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_540
timestamp 1688980957
transform 1 0 50784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_552
timestamp 1688980957
transform 1 0 51888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_561
timestamp 1688980957
transform 1 0 52716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_565
timestamp 1688980957
transform 1 0 53084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_583
timestamp 1688980957
transform 1 0 54740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_589
timestamp 1688980957
transform 1 0 55292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_611
timestamp 1688980957
transform 1 0 57316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_33
timestamp 1688980957
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_45
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_94
timestamp 1688980957
transform 1 0 9752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_98
timestamp 1688980957
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_102
timestamp 1688980957
transform 1 0 10488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_114
timestamp 1688980957
transform 1 0 11592 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_120
timestamp 1688980957
transform 1 0 12144 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_150
timestamp 1688980957
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_154
timestamp 1688980957
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_202
timestamp 1688980957
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_239
timestamp 1688980957
transform 1 0 23092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_264
timestamp 1688980957
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_268
timestamp 1688980957
transform 1 0 25760 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_274
timestamp 1688980957
transform 1 0 26312 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_279
timestamp 1688980957
transform 1 0 26772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_291
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_294
timestamp 1688980957
transform 1 0 28152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_317
timestamp 1688980957
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_331
timestamp 1688980957
transform 1 0 31556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_359
timestamp 1688980957
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_393
timestamp 1688980957
transform 1 0 37260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_414
timestamp 1688980957
transform 1 0 39192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_418
timestamp 1688980957
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_453
timestamp 1688980957
transform 1 0 42780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_488
timestamp 1688980957
transform 1 0 46000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_492
timestamp 1688980957
transform 1 0 46368 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_517
timestamp 1688980957
transform 1 0 48668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_521
timestamp 1688980957
transform 1 0 49036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_528
timestamp 1688980957
transform 1 0 49680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_557
timestamp 1688980957
transform 1 0 52348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_563
timestamp 1688980957
transform 1 0 52900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_585
timestamp 1688980957
transform 1 0 54924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_597
timestamp 1688980957
transform 1 0 56028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_623
timestamp 1688980957
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_30
timestamp 1688980957
transform 1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_48
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_61
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_163
timestamp 1688980957
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1688980957
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_206
timestamp 1688980957
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_219
timestamp 1688980957
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_259
timestamp 1688980957
transform 1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_289
timestamp 1688980957
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_362
timestamp 1688980957
transform 1 0 34408 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_366
timestamp 1688980957
transform 1 0 34776 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_386
timestamp 1688980957
transform 1 0 36616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_432
timestamp 1688980957
transform 1 0 40848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_436
timestamp 1688980957
transform 1 0 41216 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_439
timestamp 1688980957
transform 1 0 41492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_445
timestamp 1688980957
transform 1 0 42044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_481
timestamp 1688980957
transform 1 0 45356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_485
timestamp 1688980957
transform 1 0 45724 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_514
timestamp 1688980957
transform 1 0 48392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_518
timestamp 1688980957
transform 1 0 48760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_556
timestamp 1688980957
transform 1 0 52256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_561
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_579
timestamp 1688980957
transform 1 0 54372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_610
timestamp 1688980957
transform 1 0 57224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_614
timestamp 1688980957
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_42
timestamp 1688980957
transform 1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_62
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_70
timestamp 1688980957
transform 1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_99
timestamp 1688980957
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_169
timestamp 1688980957
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1688980957
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_234
timestamp 1688980957
transform 1 0 22632 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_238
timestamp 1688980957
transform 1 0 23000 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_242
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_246
timestamp 1688980957
transform 1 0 23736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1688980957
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_259
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_286
timestamp 1688980957
transform 1 0 27416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_325
timestamp 1688980957
transform 1 0 31004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 1688980957
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_392
timestamp 1688980957
transform 1 0 37168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_417
timestamp 1688980957
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_429
timestamp 1688980957
transform 1 0 40572 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_460
timestamp 1688980957
transform 1 0 43424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_464
timestamp 1688980957
transform 1 0 43792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 1688980957
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_493
timestamp 1688980957
transform 1 0 46460 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_497
timestamp 1688980957
transform 1 0 46828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_517
timestamp 1688980957
transform 1 0 48668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_521
timestamp 1688980957
transform 1 0 49036 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_529
timestamp 1688980957
transform 1 0 49772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_559
timestamp 1688980957
transform 1 0 52532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_589
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_597
timestamp 1688980957
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_624
timestamp 1688980957
transform 1 0 58512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_45
timestamp 1688980957
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_61
timestamp 1688980957
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_75
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_83
timestamp 1688980957
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_202
timestamp 1688980957
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_206
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_258
timestamp 1688980957
transform 1 0 24840 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_264
timestamp 1688980957
transform 1 0 25392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1688980957
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_289
timestamp 1688980957
transform 1 0 27692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_295
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_298
timestamp 1688980957
transform 1 0 28520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_322
timestamp 1688980957
transform 1 0 30728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_327
timestamp 1688980957
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_341
timestamp 1688980957
transform 1 0 32476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_345
timestamp 1688980957
transform 1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_364
timestamp 1688980957
transform 1 0 34592 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_387
timestamp 1688980957
transform 1 0 36708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_401
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_424
timestamp 1688980957
transform 1 0 40112 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_436
timestamp 1688980957
transform 1 0 41216 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_444
timestamp 1688980957
transform 1 0 41952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_457
timestamp 1688980957
transform 1 0 43148 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_486
timestamp 1688980957
transform 1 0 45816 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_500
timestamp 1688980957
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_505
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_515
timestamp 1688980957
transform 1 0 48484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_527
timestamp 1688980957
transform 1 0 49588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_535
timestamp 1688980957
transform 1 0 50324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_547
timestamp 1688980957
transform 1 0 51428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_551
timestamp 1688980957
transform 1 0 51796 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 1688980957
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_573
timestamp 1688980957
transform 1 0 53820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_578
timestamp 1688980957
transform 1 0 54280 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_582
timestamp 1688980957
transform 1 0 54648 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_594
timestamp 1688980957
transform 1 0 55752 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_602
timestamp 1688980957
transform 1 0 56488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_611
timestamp 1688980957
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1688980957
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_617
timestamp 1688980957
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1688980957
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1688980957
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_48
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_73
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_90
timestamp 1688980957
transform 1 0 9384 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1688980957
transform 1 0 10304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_125
timestamp 1688980957
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_214
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_218
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_222
timestamp 1688980957
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_234
timestamp 1688980957
transform 1 0 22632 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_242
timestamp 1688980957
transform 1 0 23368 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_261
timestamp 1688980957
transform 1 0 25116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_267
timestamp 1688980957
transform 1 0 25668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_271
timestamp 1688980957
transform 1 0 26036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_329
timestamp 1688980957
transform 1 0 31372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_338
timestamp 1688980957
transform 1 0 32200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_346
timestamp 1688980957
transform 1 0 32936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_350
timestamp 1688980957
transform 1 0 33304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_358
timestamp 1688980957
transform 1 0 34040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_362
timestamp 1688980957
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_373
timestamp 1688980957
transform 1 0 35420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_384
timestamp 1688980957
transform 1 0 36432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_396
timestamp 1688980957
transform 1 0 37536 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_405
timestamp 1688980957
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_409
timestamp 1688980957
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_417
timestamp 1688980957
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_425
timestamp 1688980957
transform 1 0 40204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_429
timestamp 1688980957
transform 1 0 40572 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_435
timestamp 1688980957
transform 1 0 41124 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_469
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_473
timestamp 1688980957
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_486
timestamp 1688980957
transform 1 0 45816 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_490
timestamp 1688980957
transform 1 0 46184 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_494
timestamp 1688980957
transform 1 0 46552 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_498
timestamp 1688980957
transform 1 0 46920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_502
timestamp 1688980957
transform 1 0 47288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_505
timestamp 1688980957
transform 1 0 47564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_513
timestamp 1688980957
transform 1 0 48300 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_516
timestamp 1688980957
transform 1 0 48576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_520
timestamp 1688980957
transform 1 0 48944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_526
timestamp 1688980957
transform 1 0 49496 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_557
timestamp 1688980957
transform 1 0 52348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_561
timestamp 1688980957
transform 1 0 52716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_565
timestamp 1688980957
transform 1 0 53084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_573
timestamp 1688980957
transform 1 0 53820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_577
timestamp 1688980957
transform 1 0 54188 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_585
timestamp 1688980957
transform 1 0 54924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_589
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_597
timestamp 1688980957
transform 1 0 56028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_618
timestamp 1688980957
transform 1 0 57960 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_624
timestamp 1688980957
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_29
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_41
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_46
timestamp 1688980957
transform 1 0 5336 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_73
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_89
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_108
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_129
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_154
timestamp 1688980957
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_158
timestamp 1688980957
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_164
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_185
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_216
timestamp 1688980957
transform 1 0 20976 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_266
timestamp 1688980957
transform 1 0 25576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_270
timestamp 1688980957
transform 1 0 25944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_296
timestamp 1688980957
transform 1 0 28336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_307
timestamp 1688980957
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_311
timestamp 1688980957
transform 1 0 29716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_341
timestamp 1688980957
transform 1 0 32476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_369
timestamp 1688980957
transform 1 0 35052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_402
timestamp 1688980957
transform 1 0 38088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_406
timestamp 1688980957
transform 1 0 38456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_433
timestamp 1688980957
transform 1 0 40940 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_439
timestamp 1688980957
transform 1 0 41492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_453
timestamp 1688980957
transform 1 0 42780 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_514
timestamp 1688980957
transform 1 0 48392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_556
timestamp 1688980957
transform 1 0 52256 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_561
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_586
timestamp 1688980957
transform 1 0 55016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_590
timestamp 1688980957
transform 1 0 55384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_594
timestamp 1688980957
transform 1 0 55752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_614
timestamp 1688980957
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_116
timestamp 1688980957
transform 1 0 11776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_159
timestamp 1688980957
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_190
timestamp 1688980957
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_210
timestamp 1688980957
transform 1 0 20424 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_222
timestamp 1688980957
transform 1 0 21528 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_234
timestamp 1688980957
transform 1 0 22632 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_262
timestamp 1688980957
transform 1 0 25208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_266
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 1688980957
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_337
timestamp 1688980957
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_359
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_374
timestamp 1688980957
transform 1 0 35512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_378
timestamp 1688980957
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_396
timestamp 1688980957
transform 1 0 37536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_430
timestamp 1688980957
transform 1 0 40664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_457
timestamp 1688980957
transform 1 0 43148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_470
timestamp 1688980957
transform 1 0 44344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_487
timestamp 1688980957
transform 1 0 45908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_491
timestamp 1688980957
transform 1 0 46276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_551
timestamp 1688980957
transform 1 0 51796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_555
timestamp 1688980957
transform 1 0 52164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_559
timestamp 1688980957
transform 1 0 52532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_586
timestamp 1688980957
transform 1 0 55016 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_619
timestamp 1688980957
transform 1 0 58052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_623
timestamp 1688980957
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_80
timestamp 1688980957
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_84
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_108
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_145
timestamp 1688980957
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_158
timestamp 1688980957
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_199
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_245
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1688980957
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_302
timestamp 1688980957
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_308
timestamp 1688980957
transform 1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_312
timestamp 1688980957
transform 1 0 29808 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_315
timestamp 1688980957
transform 1 0 30084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_345
timestamp 1688980957
transform 1 0 32844 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_379
timestamp 1688980957
transform 1 0 35972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_383
timestamp 1688980957
transform 1 0 36340 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_402
timestamp 1688980957
transform 1 0 38088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_406
timestamp 1688980957
transform 1 0 38456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_426
timestamp 1688980957
transform 1 0 40296 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_430
timestamp 1688980957
transform 1 0 40664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_442
timestamp 1688980957
transform 1 0 41768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_479
timestamp 1688980957
transform 1 0 45172 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_491
timestamp 1688980957
transform 1 0 46276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_495
timestamp 1688980957
transform 1 0 46644 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_522
timestamp 1688980957
transform 1 0 49128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_557
timestamp 1688980957
transform 1 0 52348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_561
timestamp 1688980957
transform 1 0 52716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_591
timestamp 1688980957
transform 1 0 55476 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_597
timestamp 1688980957
transform 1 0 56028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_33
timestamp 1688980957
transform 1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_105
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_117
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_124
timestamp 1688980957
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_136
timestamp 1688980957
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_180
timestamp 1688980957
transform 1 0 17664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_205
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_225
timestamp 1688980957
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_237
timestamp 1688980957
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_257
timestamp 1688980957
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_274
timestamp 1688980957
transform 1 0 26312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_278
timestamp 1688980957
transform 1 0 26680 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_281
timestamp 1688980957
transform 1 0 26956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_293
timestamp 1688980957
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_305
timestamp 1688980957
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_325
timestamp 1688980957
transform 1 0 31004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_330
timestamp 1688980957
transform 1 0 31464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_336
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_340
timestamp 1688980957
transform 1 0 32384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_346
timestamp 1688980957
transform 1 0 32936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_350
timestamp 1688980957
transform 1 0 33304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_354
timestamp 1688980957
transform 1 0 33672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_373
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_385
timestamp 1688980957
transform 1 0 36524 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_393
timestamp 1688980957
transform 1 0 37260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_429
timestamp 1688980957
transform 1 0 40572 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_441
timestamp 1688980957
transform 1 0 41676 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_449
timestamp 1688980957
transform 1 0 42412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_458
timestamp 1688980957
transform 1 0 43240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_468
timestamp 1688980957
transform 1 0 44160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_473
timestamp 1688980957
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 1688980957
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_501
timestamp 1688980957
transform 1 0 47196 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_505
timestamp 1688980957
transform 1 0 47564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_513
timestamp 1688980957
transform 1 0 48300 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_524
timestamp 1688980957
transform 1 0 49312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_528
timestamp 1688980957
transform 1 0 49680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_533
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_564
timestamp 1688980957
transform 1 0 52992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_573
timestamp 1688980957
transform 1 0 53820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_578
timestamp 1688980957
transform 1 0 54280 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_586
timestamp 1688980957
transform 1 0 55016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_589
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_597
timestamp 1688980957
transform 1 0 56028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_619
timestamp 1688980957
transform 1 0 58052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp 1688980957
transform 1 0 2116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_37
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_45
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_66
timestamp 1688980957
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_70
timestamp 1688980957
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_74
timestamp 1688980957
transform 1 0 7912 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_83
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_95
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_130
timestamp 1688980957
transform 1 0 13064 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_151
timestamp 1688980957
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_163
timestamp 1688980957
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_191
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_195
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_233
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_241
timestamp 1688980957
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_260
timestamp 1688980957
transform 1 0 25024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_296
timestamp 1688980957
transform 1 0 28336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_306
timestamp 1688980957
transform 1 0 29256 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_379
timestamp 1688980957
transform 1 0 35972 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_385
timestamp 1688980957
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_388
timestamp 1688980957
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_397
timestamp 1688980957
transform 1 0 37628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_401
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_407
timestamp 1688980957
transform 1 0 38548 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_416
timestamp 1688980957
transform 1 0 39376 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_421
timestamp 1688980957
transform 1 0 39836 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_433
timestamp 1688980957
transform 1 0 40940 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_444
timestamp 1688980957
transform 1 0 41952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_471
timestamp 1688980957
transform 1 0 44436 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_475
timestamp 1688980957
transform 1 0 44804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_487
timestamp 1688980957
transform 1 0 45908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_493
timestamp 1688980957
transform 1 0 46460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_514
timestamp 1688980957
transform 1 0 48392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_555
timestamp 1688980957
transform 1 0 52164 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 1688980957
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_561
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_579
timestamp 1688980957
transform 1 0 54372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_589
timestamp 1688980957
transform 1 0 55292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_593
timestamp 1688980957
transform 1 0 55660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_614
timestamp 1688980957
transform 1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1688980957
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_62
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_66
timestamp 1688980957
transform 1 0 7176 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_114
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_157
timestamp 1688980957
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_262
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_266
timestamp 1688980957
transform 1 0 25576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_304
timestamp 1688980957
transform 1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_337
timestamp 1688980957
transform 1 0 32108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_360
timestamp 1688980957
transform 1 0 34224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_382
timestamp 1688980957
transform 1 0 36248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_386
timestamp 1688980957
transform 1 0 36616 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_406
timestamp 1688980957
transform 1 0 38456 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_418
timestamp 1688980957
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_489
timestamp 1688980957
transform 1 0 46092 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_522
timestamp 1688980957
transform 1 0 49128 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_537
timestamp 1688980957
transform 1 0 50508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_558
timestamp 1688980957
transform 1 0 52440 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 1688980957
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_619
timestamp 1688980957
transform 1 0 58052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_623
timestamp 1688980957
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_35
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_92
timestamp 1688980957
transform 1 0 9568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_122
timestamp 1688980957
transform 1 0 12328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_146
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_158
timestamp 1688980957
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_185
timestamp 1688980957
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_195
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_199
timestamp 1688980957
transform 1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_219
timestamp 1688980957
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_253
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_267
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_289
timestamp 1688980957
transform 1 0 27692 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_298
timestamp 1688980957
transform 1 0 28520 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_310
timestamp 1688980957
transform 1 0 29624 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_316
timestamp 1688980957
transform 1 0 30176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_373
timestamp 1688980957
transform 1 0 35420 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1688980957
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_433
timestamp 1688980957
transform 1 0 40940 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_444
timestamp 1688980957
transform 1 0 41952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_478
timestamp 1688980957
transform 1 0 45080 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_482
timestamp 1688980957
transform 1 0 45448 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_494
timestamp 1688980957
transform 1 0 46552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_500
timestamp 1688980957
transform 1 0 47104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_522
timestamp 1688980957
transform 1 0 49128 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_547
timestamp 1688980957
transform 1 0 51428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_551
timestamp 1688980957
transform 1 0 51796 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_557
timestamp 1688980957
transform 1 0 52348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_561
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_565
timestamp 1688980957
transform 1 0 53084 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_592
timestamp 1688980957
transform 1 0 55568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_596
timestamp 1688980957
transform 1 0 55936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_11
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_114
timestamp 1688980957
transform 1 0 11592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_123
timestamp 1688980957
transform 1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_128
timestamp 1688980957
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1688980957
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_169
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_213
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_222
timestamp 1688980957
transform 1 0 21528 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_234
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_261
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_267
timestamp 1688980957
transform 1 0 25668 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1688980957
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_288
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1688980957
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_325
timestamp 1688980957
transform 1 0 31004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_329
timestamp 1688980957
transform 1 0 31372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_337
timestamp 1688980957
transform 1 0 32108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_349
timestamp 1688980957
transform 1 0 33212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_361
timestamp 1688980957
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_381
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_408
timestamp 1688980957
transform 1 0 38640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_412
timestamp 1688980957
transform 1 0 39008 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_415
timestamp 1688980957
transform 1 0 39284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1688980957
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_451
timestamp 1688980957
transform 1 0 42596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_470
timestamp 1688980957
transform 1 0 44344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_474
timestamp 1688980957
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_486
timestamp 1688980957
transform 1 0 45816 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_498
timestamp 1688980957
transform 1 0 46920 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_506
timestamp 1688980957
transform 1 0 47656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_515
timestamp 1688980957
transform 1 0 48484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_524
timestamp 1688980957
transform 1 0 49312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_541
timestamp 1688980957
transform 1 0 50876 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 1688980957
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_557
timestamp 1688980957
transform 1 0 52348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_565
timestamp 1688980957
transform 1 0 53084 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_574
timestamp 1688980957
transform 1 0 53912 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_586
timestamp 1688980957
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_620
timestamp 1688980957
transform 1 0 58144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_624
timestamp 1688980957
transform 1 0 58512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_41
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_45
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_96
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_124
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_128
timestamp 1688980957
transform 1 0 12880 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_185
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_189
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_199
timestamp 1688980957
transform 1 0 19412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_207
timestamp 1688980957
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 1688980957
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_229
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_241
timestamp 1688980957
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_268
timestamp 1688980957
transform 1 0 25760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_272
timestamp 1688980957
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_333
timestamp 1688980957
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_353
timestamp 1688980957
transform 1 0 33580 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_359
timestamp 1688980957
transform 1 0 34132 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_362
timestamp 1688980957
transform 1 0 34408 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_376
timestamp 1688980957
transform 1 0 35696 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_388
timestamp 1688980957
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_397
timestamp 1688980957
transform 1 0 37628 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_424
timestamp 1688980957
transform 1 0 40112 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_436
timestamp 1688980957
transform 1 0 41216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_442
timestamp 1688980957
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_457
timestamp 1688980957
transform 1 0 43148 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_484
timestamp 1688980957
transform 1 0 45632 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_496
timestamp 1688980957
transform 1 0 46736 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_502
timestamp 1688980957
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_505
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_523
timestamp 1688980957
transform 1 0 49220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_535
timestamp 1688980957
transform 1 0 50324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_547
timestamp 1688980957
transform 1 0 51428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 1688980957
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_561
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_567
timestamp 1688980957
transform 1 0 53268 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_571
timestamp 1688980957
transform 1 0 53636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_583
timestamp 1688980957
transform 1 0 54740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_591
timestamp 1688980957
transform 1 0 55476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_595
timestamp 1688980957
transform 1 0 55844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_600
timestamp 1688980957
transform 1 0 56304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_613
timestamp 1688980957
transform 1 0 57500 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_46
timestamp 1688980957
transform 1 0 5336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_50
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_68
timestamp 1688980957
transform 1 0 7360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_76
timestamp 1688980957
transform 1 0 8096 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_79
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_118
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_166
timestamp 1688980957
transform 1 0 16376 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_232
timestamp 1688980957
transform 1 0 22448 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_244
timestamp 1688980957
transform 1 0 23552 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_248
timestamp 1688980957
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_281
timestamp 1688980957
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_298
timestamp 1688980957
transform 1 0 28520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_302
timestamp 1688980957
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_315
timestamp 1688980957
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_332
timestamp 1688980957
transform 1 0 31648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_336
timestamp 1688980957
transform 1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_355
timestamp 1688980957
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_359
timestamp 1688980957
transform 1 0 34132 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_374
timestamp 1688980957
transform 1 0 35512 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_386
timestamp 1688980957
transform 1 0 36616 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_393
timestamp 1688980957
transform 1 0 37260 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_416
timestamp 1688980957
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_449
timestamp 1688980957
transform 1 0 42412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_453
timestamp 1688980957
transform 1 0 42780 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_459
timestamp 1688980957
transform 1 0 43332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_471
timestamp 1688980957
transform 1 0 44436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_501
timestamp 1688980957
transform 1 0 47196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_518
timestamp 1688980957
transform 1 0 48760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 1688980957
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_541
timestamp 1688980957
transform 1 0 50876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_545
timestamp 1688980957
transform 1 0 51244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_573
timestamp 1688980957
transform 1 0 53820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_577
timestamp 1688980957
transform 1 0 54188 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_585
timestamp 1688980957
transform 1 0 54924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_598
timestamp 1688980957
transform 1 0 56120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_624
timestamp 1688980957
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_94
timestamp 1688980957
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_122
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_197
timestamp 1688980957
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_242
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_308
timestamp 1688980957
transform 1 0 29440 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_314
timestamp 1688980957
transform 1 0 29992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_331
timestamp 1688980957
transform 1 0 31556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_378
timestamp 1688980957
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_426
timestamp 1688980957
transform 1 0 40296 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_466
timestamp 1688980957
transform 1 0 43976 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_472
timestamp 1688980957
transform 1 0 44528 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_500
timestamp 1688980957
transform 1 0 47104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_542
timestamp 1688980957
transform 1 0 50968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_570
timestamp 1688980957
transform 1 0 53544 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_611
timestamp 1688980957
transform 1 0 57316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 1688980957
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_38
timestamp 1688980957
transform 1 0 4600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_50
timestamp 1688980957
transform 1 0 5704 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_75
timestamp 1688980957
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_79
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_94
timestamp 1688980957
transform 1 0 9752 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_98
timestamp 1688980957
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_126
timestamp 1688980957
transform 1 0 12696 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_158
timestamp 1688980957
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_170
timestamp 1688980957
transform 1 0 16744 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_176
timestamp 1688980957
transform 1 0 17296 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_238
timestamp 1688980957
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_270
timestamp 1688980957
transform 1 0 25944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_274
timestamp 1688980957
transform 1 0 26312 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_303
timestamp 1688980957
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_317
timestamp 1688980957
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_340
timestamp 1688980957
transform 1 0 32384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_344
timestamp 1688980957
transform 1 0 32752 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_415
timestamp 1688980957
transform 1 0 39284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1688980957
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_477
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_526
timestamp 1688980957
transform 1 0 49496 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_533
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_543
timestamp 1688980957
transform 1 0 51060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_547
timestamp 1688980957
transform 1 0 51428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_573
timestamp 1688980957
transform 1 0 53820 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_577
timestamp 1688980957
transform 1 0 54188 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_585
timestamp 1688980957
transform 1 0 54924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_589
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_615
timestamp 1688980957
transform 1 0 57684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_623
timestamp 1688980957
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_34
timestamp 1688980957
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_46
timestamp 1688980957
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_79
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_92
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_96
timestamp 1688980957
transform 1 0 9936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_141
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_160
timestamp 1688980957
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_177
timestamp 1688980957
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_187
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_195
timestamp 1688980957
transform 1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_219
timestamp 1688980957
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_234
timestamp 1688980957
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_238
timestamp 1688980957
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_242
timestamp 1688980957
transform 1 0 23368 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_259
timestamp 1688980957
transform 1 0 24932 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_263
timestamp 1688980957
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1688980957
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_294
timestamp 1688980957
transform 1 0 28152 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_303
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_315
timestamp 1688980957
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_319
timestamp 1688980957
transform 1 0 30452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_328
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_332
timestamp 1688980957
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_345
timestamp 1688980957
transform 1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_371
timestamp 1688980957
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_383
timestamp 1688980957
transform 1 0 36340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_387
timestamp 1688980957
transform 1 0 36708 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_390
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_417
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_421
timestamp 1688980957
transform 1 0 39836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_433
timestamp 1688980957
transform 1 0 40940 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_437
timestamp 1688980957
transform 1 0 41308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_470
timestamp 1688980957
transform 1 0 44344 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_474
timestamp 1688980957
transform 1 0 44712 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_490
timestamp 1688980957
transform 1 0 46184 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_496
timestamp 1688980957
transform 1 0 46736 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_499
timestamp 1688980957
transform 1 0 47012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 1688980957
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_505
timestamp 1688980957
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_509
timestamp 1688980957
transform 1 0 47932 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_513
timestamp 1688980957
transform 1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_517
timestamp 1688980957
transform 1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_521
timestamp 1688980957
transform 1 0 49036 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_531
timestamp 1688980957
transform 1 0 49956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_535
timestamp 1688980957
transform 1 0 50324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_547
timestamp 1688980957
transform 1 0 51428 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_553
timestamp 1688980957
transform 1 0 51980 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_556
timestamp 1688980957
transform 1 0 52256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_571
timestamp 1688980957
transform 1 0 53636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_583
timestamp 1688980957
transform 1 0 54740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_591
timestamp 1688980957
transform 1 0 55476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_594
timestamp 1688980957
transform 1 0 55752 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_603
timestamp 1688980957
transform 1 0 56580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 1688980957
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_617
timestamp 1688980957
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_57
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_94
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_122
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1688980957
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_130
timestamp 1688980957
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_173
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_190
timestamp 1688980957
transform 1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_205
timestamp 1688980957
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_225
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_234
timestamp 1688980957
transform 1 0 22632 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_270
timestamp 1688980957
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_290
timestamp 1688980957
transform 1 0 27784 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_304
timestamp 1688980957
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_335
timestamp 1688980957
transform 1 0 31924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_339
timestamp 1688980957
transform 1 0 32292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_358
timestamp 1688980957
transform 1 0 34040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 1688980957
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_373
timestamp 1688980957
transform 1 0 35420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_396
timestamp 1688980957
transform 1 0 37536 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_400
timestamp 1688980957
transform 1 0 37904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_417
timestamp 1688980957
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_429
timestamp 1688980957
transform 1 0 40572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_443
timestamp 1688980957
transform 1 0 41860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_447
timestamp 1688980957
transform 1 0 42228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_451
timestamp 1688980957
transform 1 0 42596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_461
timestamp 1688980957
transform 1 0 43516 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_474
timestamp 1688980957
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_477
timestamp 1688980957
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_505
timestamp 1688980957
transform 1 0 47564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_509
timestamp 1688980957
transform 1 0 47932 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_527
timestamp 1688980957
transform 1 0 49588 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 1688980957
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_541
timestamp 1688980957
transform 1 0 50876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_545
timestamp 1688980957
transform 1 0 51244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_572
timestamp 1688980957
transform 1 0 53728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_576
timestamp 1688980957
transform 1 0 54096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_580
timestamp 1688980957
transform 1 0 54464 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_613
timestamp 1688980957
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_100
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_122
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_173
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_199
timestamp 1688980957
transform 1 0 19412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_242
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_306
timestamp 1688980957
transform 1 0 29256 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_369
timestamp 1688980957
transform 1 0 35052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_397
timestamp 1688980957
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_428
timestamp 1688980957
transform 1 0 40480 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_436
timestamp 1688980957
transform 1 0 41216 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_439
timestamp 1688980957
transform 1 0 41492 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_465
timestamp 1688980957
transform 1 0 43884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 1688980957
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_542
timestamp 1688980957
transform 1 0 50968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_570
timestamp 1688980957
transform 1 0 53544 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_610
timestamp 1688980957
transform 1 0 57224 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_617
timestamp 1688980957
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_33
timestamp 1688980957
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_60
timestamp 1688980957
transform 1 0 6624 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_64
timestamp 1688980957
transform 1 0 6992 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_95
timestamp 1688980957
transform 1 0 9844 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1688980957
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_163
timestamp 1688980957
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_175
timestamp 1688980957
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_190
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1688980957
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_238
timestamp 1688980957
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_270
timestamp 1688980957
transform 1 0 25944 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_335
timestamp 1688980957
transform 1 0 31924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_339
timestamp 1688980957
transform 1 0 32292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_343
timestamp 1688980957
transform 1 0 32660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_361
timestamp 1688980957
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_373
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_403
timestamp 1688980957
transform 1 0 38180 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_416
timestamp 1688980957
transform 1 0 39376 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_445
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_472
timestamp 1688980957
transform 1 0 44528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_481
timestamp 1688980957
transform 1 0 45356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_513
timestamp 1688980957
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_525
timestamp 1688980957
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_529
timestamp 1688980957
transform 1 0 49772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_549
timestamp 1688980957
transform 1 0 51612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_553
timestamp 1688980957
transform 1 0 51980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_580
timestamp 1688980957
transform 1 0 54464 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_615
timestamp 1688980957
transform 1 0 57684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_623
timestamp 1688980957
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_29
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_50
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_83
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_129
timestamp 1688980957
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_141
timestamp 1688980957
transform 1 0 14076 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_157
timestamp 1688980957
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_192
timestamp 1688980957
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_197
timestamp 1688980957
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_209
timestamp 1688980957
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_229
timestamp 1688980957
transform 1 0 22172 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_241
timestamp 1688980957
transform 1 0 23276 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_253
timestamp 1688980957
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_259
timestamp 1688980957
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_271
timestamp 1688980957
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_292
timestamp 1688980957
transform 1 0 27968 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_301
timestamp 1688980957
transform 1 0 28796 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_307
timestamp 1688980957
transform 1 0 29348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_309
timestamp 1688980957
transform 1 0 29532 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_318
timestamp 1688980957
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_330
timestamp 1688980957
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_341
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_358
timestamp 1688980957
transform 1 0 34040 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_363
timestamp 1688980957
transform 1 0 34500 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_365
timestamp 1688980957
transform 1 0 34684 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_377
timestamp 1688980957
transform 1 0 35788 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_389
timestamp 1688980957
transform 1 0 36892 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_409
timestamp 1688980957
transform 1 0 38732 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_413
timestamp 1688980957
transform 1 0 39100 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_419
timestamp 1688980957
transform 1 0 39652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_421
timestamp 1688980957
transform 1 0 39836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_430
timestamp 1688980957
transform 1 0 40664 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_442
timestamp 1688980957
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_477
timestamp 1688980957
transform 1 0 44988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_487
timestamp 1688980957
transform 1 0 45908 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_497
timestamp 1688980957
transform 1 0 46828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_501
timestamp 1688980957
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_513
timestamp 1688980957
transform 1 0 48300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_523
timestamp 1688980957
transform 1 0 49220 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_531
timestamp 1688980957
transform 1 0 49956 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_533
timestamp 1688980957
transform 1 0 50140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_545
timestamp 1688980957
transform 1 0 51244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_555
timestamp 1688980957
transform 1 0 52164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 1688980957
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_561
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_570
timestamp 1688980957
transform 1 0 53544 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_574
timestamp 1688980957
transform 1 0 53912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_586
timestamp 1688980957
transform 1 0 55016 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_589
timestamp 1688980957
transform 1 0 55292 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_605
timestamp 1688980957
transform 1 0 56764 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_613
timestamp 1688980957
transform 1 0 57500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_617
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 34040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold5
timestamp 1688980957
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 24840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 35420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 33948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 24196 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 22632 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 42136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold12
timestamp 1688980957
transform -1 0 41584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 38180 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold17
timestamp 1688980957
transform -1 0 50048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 50508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold20
timestamp 1688980957
transform -1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 43976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 42320 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 43148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 41584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 27692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 26680 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 24472 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 23736 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 36892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold31
timestamp 1688980957
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 37720 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 24196 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 23184 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 31096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 29440 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 41124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 40572 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 21620 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 26772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 31924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 29440 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 47472 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 46000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 35236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 37812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform -1 0 36156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 37720 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 37996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 39008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 40572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 34684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 34408 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 48300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 46736 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 36800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 35236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 43976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 44712 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 42136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 41400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 44620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 41584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 47196 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 35420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 41400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 39744 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 39192 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 37996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 27968 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 47288 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 46460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 51796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 51704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 30728 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold86
timestamp 1688980957
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 34592 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 30728 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 29348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 31188 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 58604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold93
timestamp 1688980957
transform -1 0 55384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 54004 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 29716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 28152 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 56028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 55200 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 33764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 34132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 18216 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold104
timestamp 1688980957
transform -1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 14628 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 43148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold107
timestamp 1688980957
transform 1 0 39560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 40572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 58604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold110
timestamp 1688980957
transform -1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform 1 0 51888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 58236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 58604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 19688 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 18492 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 20792 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 19320 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 58512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 57316 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 20792 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 22264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 34316 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold127
timestamp 1688980957
transform -1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 5152 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 51612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 51980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold132
timestamp 1688980957
transform -1 0 51060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 47104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 57500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 56396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 58604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 58236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 54280 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 52624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 29440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 27048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 5796 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform -1 0 5060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 48484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform -1 0 48668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 19136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 16100 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 54924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 54188 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 51428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 51796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 48300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold159
timestamp 1688980957
transform -1 0 45724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform 1 0 41860 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 24932 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 23644 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform -1 0 16560 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold166
timestamp 1688980957
transform 1 0 17296 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform -1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 45816 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 46460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 10488 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 37260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 36524 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform -1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 44160 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 45172 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 39560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 40940 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 9752 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold185
timestamp 1688980957
transform -1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 23920 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 26772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 25208 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 25116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 24196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 58604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 55752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 38364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform -1 0 37536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 12420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 11592 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform -1 0 27416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 25484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 55016 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 54280 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform -1 0 50876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 48392 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 2024 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 58420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 58604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform -1 0 22540 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 21712 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold212
timestamp 1688980957
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 15272 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform -1 0 52348 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 51152 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 43240 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 42320 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform -1 0 45908 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 47196 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 40480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform 1 0 40480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform -1 0 22724 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 22356 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 23092 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform -1 0 48484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 48668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 55752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 58604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 40572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 38364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 50968 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold235
timestamp 1688980957
transform -1 0 51704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 50876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 49312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 47748 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 19044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 45724 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 45632 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 19872 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold244
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 19412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 56028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform 1 0 52256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform -1 0 52348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 51612 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform -1 0 22724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 21528 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform -1 0 37996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 36432 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform -1 0 21804 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 22540 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform -1 0 18676 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform -1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 44252 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform -1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform -1 0 10764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform -1 0 50048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform -1 0 47472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold269
timestamp 1688980957
transform -1 0 34500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform -1 0 32016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 43516 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 42320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform -1 0 19044 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform -1 0 18492 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 52256 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform -1 0 52348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform 1 0 54464 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold278
timestamp 1688980957
transform 1 0 57408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 57960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 49312 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform -1 0 49128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 32016 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 31004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform -1 0 18492 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform -1 0 13984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform -1 0 52256 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 52992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform -1 0 54832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform -1 0 54740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform -1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 11776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold297
timestamp 1688980957
transform 1 0 44344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 44896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform -1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 38180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform -1 0 37168 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 14904 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform -1 0 15272 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform -1 0 35972 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform -1 0 36248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 35420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 36156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform -1 0 32844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform -1 0 32016 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 58604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform -1 0 58144 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform -1 0 58604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform -1 0 58052 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform -1 0 58604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform -1 0 58604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform -1 0 11408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform 1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 49128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 47472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform -1 0 58604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 58512 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 32016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform -1 0 31004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 54740 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform -1 0 53820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform -1 0 55568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform -1 0 53912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform -1 0 55476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform -1 0 55016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform -1 0 55292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform -1 0 54832 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform -1 0 43148 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform -1 0 41952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform -1 0 50048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform -1 0 49312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform 1 0 27232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold342
timestamp 1688980957
transform -1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 28612 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform -1 0 26312 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform -1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform -1 0 35972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform -1 0 34500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform 1 0 44160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform -1 0 45632 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform -1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform -1 0 26496 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform -1 0 42044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold357 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform -1 0 38548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1688980957
transform -1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform -1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform 1 0 47288 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold362
timestamp 1688980957
transform -1 0 48300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform -1 0 43332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform -1 0 41952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1688980957
transform -1 0 28520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform 1 0 28520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform -1 0 25668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform -1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1688980957
transform -1 0 44528 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform -1 0 43424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform -1 0 51888 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform -1 0 52624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform -1 0 25576 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 1688980957
transform -1 0 24288 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 1688980957
transform 1 0 38548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform -1 0 40296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform -1 0 6164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold378
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform -1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform -1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform 1 0 37904 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform -1 0 14904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold383
timestamp 1688980957
transform -1 0 13984 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform -1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 1688980957
transform -1 0 15180 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform -1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform -1 0 11408 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform -1 0 44896 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform -1 0 42320 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 1688980957
transform -1 0 16652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 1688980957
transform -1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold393
timestamp 1688980957
transform 1 0 56304 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold394
timestamp 1688980957
transform -1 0 58604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold395
timestamp 1688980957
transform -1 0 56948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 1688980957
transform -1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 1688980957
transform -1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold399
timestamp 1688980957
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 1688980957
transform -1 0 52348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold401
timestamp 1688980957
transform 1 0 49312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold402
timestamp 1688980957
transform 1 0 50324 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 1688980957
transform -1 0 4508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold404
timestamp 1688980957
transform -1 0 2944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 1688980957
transform -1 0 39468 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold406
timestamp 1688980957
transform -1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold407
timestamp 1688980957
transform -1 0 36248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 1688980957
transform -1 0 37904 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold409
timestamp 1688980957
transform -1 0 37168 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 1688980957
transform -1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold411
timestamp 1688980957
transform -1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 1688980957
transform -1 0 34408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 1688980957
transform -1 0 33580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 1688980957
transform -1 0 31924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 1688980957
transform -1 0 30360 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 1688980957
transform -1 0 4876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold417
timestamp 1688980957
transform -1 0 3680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 1688980957
transform -1 0 58604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 1688980957
transform -1 0 58512 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 1688980957
transform -1 0 16376 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 1688980957
transform 1 0 14904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 1688980957
transform -1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 1688980957
transform -1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 1688980957
transform -1 0 43976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 1688980957
transform -1 0 44160 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 1688980957
transform -1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 1688980957
transform -1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 1688980957
transform -1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 1688980957
transform -1 0 13708 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 1688980957
transform -1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 1688980957
transform -1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold432
timestamp 1688980957
transform -1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 1688980957
transform 1 0 6624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 1688980957
transform -1 0 53820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 1688980957
transform -1 0 52256 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 1688980957
transform -1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold437
timestamp 1688980957
transform -1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 1688980957
transform -1 0 18124 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 1688980957
transform -1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 1688980957
transform -1 0 18308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 1688980957
transform -1 0 50876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 1688980957
transform -1 0 49220 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 1688980957
transform -1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 1688980957
transform -1 0 34868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 1688980957
transform -1 0 40572 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 1688980957
transform -1 0 39468 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 1688980957
transform -1 0 49220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 1688980957
transform -1 0 48484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 1688980957
transform -1 0 47196 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 1688980957
transform -1 0 46184 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 1688980957
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 1688980957
transform -1 0 3404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 1688980957
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 1688980957
transform -1 0 3312 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 1688980957
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 1688980957
transform -1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold457
timestamp 1688980957
transform -1 0 16100 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 1688980957
transform -1 0 13984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 1688980957
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold460
timestamp 1688980957
transform -1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 1688980957
transform -1 0 24288 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 1688980957
transform -1 0 48300 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 1688980957
transform 1 0 46092 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 1688980957
transform -1 0 32844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 1688980957
transform -1 0 31740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 1688980957
transform -1 0 12420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 1688980957
transform -1 0 11592 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 1688980957
transform -1 0 22448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 1688980957
transform 1 0 19504 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 1688980957
transform -1 0 28980 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 1688980957
transform -1 0 28152 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 1688980957
transform -1 0 28796 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 1688980957
transform -1 0 27968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 1688980957
transform -1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 1688980957
transform -1 0 19136 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 1688980957
transform -1 0 25944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 1688980957
transform -1 0 24288 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 1688980957
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 1688980957
transform -1 0 18768 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 1688980957
transform -1 0 57684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 1688980957
transform -1 0 56764 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 1688980957
transform -1 0 53636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 1688980957
transform -1 0 53820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 1688980957
transform -1 0 37996 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 1688980957
transform -1 0 36524 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 1688980957
transform -1 0 40664 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 1688980957
transform -1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 1688980957
transform -1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 1688980957
transform -1 0 25760 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 1688980957
transform 1 0 30728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 1688980957
transform -1 0 31924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 1688980957
transform -1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold493
timestamp 1688980957
transform 1 0 15364 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 1688980957
transform -1 0 47840 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 1688980957
transform -1 0 47104 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold496
timestamp 1688980957
transform 1 0 44160 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold497
timestamp 1688980957
transform -1 0 44160 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold498
timestamp 1688980957
transform -1 0 38732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 1688980957
transform -1 0 37996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 1688980957
transform -1 0 48300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold501
timestamp 1688980957
transform -1 0 47564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold502
timestamp 1688980957
transform -1 0 30268 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold503
timestamp 1688980957
transform -1 0 28980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 1688980957
transform -1 0 23368 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 1688980957
transform -1 0 22264 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold506
timestamp 1688980957
transform -1 0 23368 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold507
timestamp 1688980957
transform -1 0 23000 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold508
timestamp 1688980957
transform -1 0 50876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 1688980957
transform -1 0 51612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold511
timestamp 1688980957
transform -1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold512
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold513
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 1688980957
transform -1 0 23000 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 1688980957
transform -1 0 53544 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold516
timestamp 1688980957
transform -1 0 53728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold517
timestamp 1688980957
transform 1 0 28336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold518
timestamp 1688980957
transform -1 0 28796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 1688980957
transform -1 0 12696 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 1688980957
transform -1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold521
timestamp 1688980957
transform 1 0 33304 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 1688980957
transform -1 0 35420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 1688980957
transform -1 0 54464 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 1688980957
transform -1 0 53728 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 1688980957
transform -1 0 25944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 1688980957
transform -1 0 24288 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold527
timestamp 1688980957
transform -1 0 5704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold528
timestamp 1688980957
transform 1 0 4600 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold529
timestamp 1688980957
transform -1 0 57500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 1688980957
transform -1 0 56580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 1688980957
transform -1 0 6624 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 1688980957
transform -1 0 5704 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 1688980957
transform -1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 1688980957
transform -1 0 11408 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 1688980957
transform -1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 1688980957
transform -1 0 8372 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 1688980957
transform -1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 1688980957
transform -1 0 10488 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 1688980957
transform -1 0 5336 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 1688980957
transform -1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 1688980957
transform -1 0 6348 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 1688980957
transform -1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 1688980957
transform -1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold548
timestamp 1688980957
transform 1 0 5612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold550
timestamp 1688980957
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold551
timestamp 1688980957
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 1688980957
transform -1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 1688980957
transform -1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold554 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold555
timestamp 1688980957
transform -1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 1688980957
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 1688980957
transform -1 0 7636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold558
timestamp 1688980957
transform -1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 1688980957
transform -1 0 50876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 1688980957
transform 1 0 9108 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold561
timestamp 1688980957
transform -1 0 28888 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 1688980957
transform -1 0 36984 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold563
timestamp 1688980957
transform -1 0 54740 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 1688980957
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold565
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold566
timestamp 1688980957
transform -1 0 45080 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold567
timestamp 1688980957
transform -1 0 39468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold568
timestamp 1688980957
transform -1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold569
timestamp 1688980957
transform -1 0 45724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold570
timestamp 1688980957
transform -1 0 58604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold571
timestamp 1688980957
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold572
timestamp 1688980957
transform -1 0 33304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold573
timestamp 1688980957
transform -1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold574
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold575
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold576
timestamp 1688980957
transform -1 0 25944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold577
timestamp 1688980957
transform -1 0 51428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold578
timestamp 1688980957
transform -1 0 51244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold579
timestamp 1688980957
transform -1 0 57684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold580
timestamp 1688980957
transform 1 0 38640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold581
timestamp 1688980957
transform 1 0 33120 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold582
timestamp 1688980957
transform -1 0 38732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold583
timestamp 1688980957
transform -1 0 53452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 1688980957
transform -1 0 25116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold585
timestamp 1688980957
transform -1 0 32844 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold586
timestamp 1688980957
transform -1 0 19136 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold587
timestamp 1688980957
transform -1 0 48116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold588
timestamp 1688980957
transform -1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold589
timestamp 1688980957
transform -1 0 41032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold590
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 26956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 28612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 37996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 42320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 47748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 48392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 53820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 55660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 55384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 19872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform -1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 26404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 27048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform -1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform -1 0 29348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform -1 0 35604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform -1 0 39652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform -1 0 44436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 47012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 51796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform -1 0 49220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 51704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 55384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 57500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 55384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform -1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform -1 0 57684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform -1 0 58512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform -1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform -1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output69 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3588 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform 1 0 24196 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform -1 0 26864 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform -1 0 32016 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 33948 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform -1 0 42228 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform 1 0 46000 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform -1 0 49036 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform -1 0 52164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform 1 0 54188 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform 1 0 55660 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform 1 0 57132 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform -1 0 57132 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform -1 0 15732 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform -1 0 21712 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 24288 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 29440 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 34592 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 39744 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 44896 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 50048 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 55200 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire118
timestamp 1688980957
transform -1 0 35328 0 1 4352
box -38 -48 406 592
<< labels >>
flabel metal4 s 8166 2128 8486 21808 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 22610 2128 22930 21808 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 37054 2128 37374 21808 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 51498 2128 51818 21808 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 15388 2128 15708 21808 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 29832 2128 30152 21808 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 44276 2128 44596 21808 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 58720 2128 59040 21808 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal tristate
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal tristate
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 24000
<< end >>
