* NGSPICE file created from wishbone_nn.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt wishbone_nn vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold340 _1013_/X vssd1 vssd1 vccd1 vccd1 _1343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _1351_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 input43/X vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold395 _0600_/X vssd1 vssd1 vccd1 vccd1 _1097_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _1014_/X vssd1 vssd1 vccd1 vccd1 _1344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _1063_/Q vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0584__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0759__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1270_ _1334_/CLK _1270_/D vssd1 vssd1 vccd1 vccd1 _1270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0985_ hold48/X hold60/X _0994_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
Xfanout127 _0757_/S1 vssd1 vssd1 vccd1 vccd1 _0774_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout138 input1/X vssd1 vssd1 vccd1 vccd1 _0977_/C sky130_fd_sc_hd__buf_4
Xfanout105 _0776_/S vssd1 vssd1 vccd1 vccd1 _0708_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout116 _0647_/S vssd1 vssd1 vccd1 vccd1 _0630_/S sky130_fd_sc_hd__buf_8
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold192 _1128_/Q vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _0566_/X vssd1 vssd1 vccd1 vccd1 _1064_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0579__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1277__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _1109_/Q vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ hold651/X hold188/X hold99/X hold122/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0770_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1253_ _1343_/CLK _1253_/D vssd1 vssd1 vccd1 vccd1 _1253_/Q sky130_fd_sc_hd__dfxtp_1
X_1322_ _1359_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1184_ _1351_/CLK _1184_/D vssd1 vssd1 vccd1 vccd1 _1184_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0880__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0518__A _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0968_ hold101/X hold73/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0968_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout125_A _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0952__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0899_ _0907_/A _0899_/B vssd1 vssd1 vccd1 vccd1 _1237_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1023__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0862__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0772__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0822_ _0821_/A _0821_/B _0813_/X vssd1 vssd1 vccd1 vccd1 _0827_/B sky130_fd_sc_hd__a21oi_1
X_0753_ hold472/X hold501/X hold482/X hold507/X _0757_/S0 _0757_/S1 vssd1 vssd1 vccd1
+ vccd1 _0753_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0684_ hold661/X hold607/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0947__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1305_ _1337_/CLK _1305_/D vssd1 vssd1 vccd1 vccd1 _1305_/Q sky130_fd_sc_hd__dfxtp_1
X_1236_ _1272_/CLK _1236_/D vssd1 vssd1 vccd1 vccd1 _1236_/Q sky130_fd_sc_hd__dfxtp_1
X_1098_ _1333_/CLK _1098_/D vssd1 vssd1 vccd1 vccd1 _1098_/Q sky130_fd_sc_hd__dfxtp_1
X_1167_ _1363_/CLK _1167_/D vssd1 vssd1 vccd1 vccd1 _1167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1018__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1315__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0592__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0767__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1021_ hold351/X hold88/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1021_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0694__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0805_ hold107/X hold234/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0805_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 _0535_/X vssd1 vssd1 vccd1 vccd1 _1043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _1312_/Q vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_0667_ _0666_/X _0665_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0667_/X sky130_fd_sc_hd__mux2_1
Xhold725 _1157_/Q vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0736_ hold646/X hold585/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0736_/X sky130_fd_sc_hd__mux2_1
X_0598_ hold25/X hold347/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1219_ _1254_/CLK _1219_/D vssd1 vssd1 vccd1 vccd1 _1219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0685__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0587__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0521_ hold685/X hold313/X _0521_/S vssd1 vssd1 vccd1 vccd1 _0521_/X sky130_fd_sc_hd__mux2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1004_ hold399/X hold494/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0960__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold544 _0629_/X vssd1 vssd1 vccd1 vccd1 _1125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _0943_/X vssd1 vssd1 vccd1 vccd1 _1275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _1256_/Q vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _1353_/Q vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _0958_/X vssd1 vssd1 vccd1 vccd1 _1289_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1160__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0719_ _0718_/X _0717_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0719_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold555 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 input16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _0864_/Y vssd1 vssd1 vccd1 vccd1 _0865_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold599 _1172_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _0848_/Y vssd1 vssd1 vccd1 vccd1 _0849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _1174_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0658__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1031__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _1225_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 _1235_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput97 _1216_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0780__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0649__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1183__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0955__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold341 _1200_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold363 _0795_/X vssd1 vssd1 vccd1 vccd1 _1193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _1082_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _1086_/Q vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _1021_/X vssd1 vssd1 vccd1 vccd1 _1351_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold385 _0565_/X vssd1 vssd1 vccd1 vccd1 _1063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _1067_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1026__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1056__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0775__S _0775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0892__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0984_ hold137/X hold669/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout106 _1008_/S vssd1 vssd1 vccd1 vccd1 _0994_/S sky130_fd_sc_hd__buf_6
Xfanout139 input1/X vssd1 vssd1 vccd1 vccd1 _0907_/A sky130_fd_sc_hd__buf_4
Xfanout117 _0614_/S vssd1 vssd1 vccd1 vccd1 _0612_/S sky130_fd_sc_hd__buf_8
Xfanout128 _0757_/S1 vssd1 vssd1 vccd1 vccd1 _0734_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0730__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 _0632_/X vssd1 vssd1 vccd1 vccd1 _1128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _1260_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold171 _0612_/X vssd1 vssd1 vccd1 vccd1 _1109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _1069_/Q vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0595__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0874__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0721__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1321_ _1321_/CLK _1321_/D vssd1 vssd1 vccd1 vccd1 _1321_/Q sky130_fd_sc_hd__dfxtp_1
X_1252_ _1351_/CLK _1252_/D vssd1 vssd1 vccd1 vccd1 _1252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1183_ _1346_/CLK hold49/X vssd1 vssd1 vccd1 vccd1 _1183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0967_ hold54/X hold45/X _0976_/S vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__mux2_1
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0898_ _1237_/Q _0906_/A2 _0908_/B1 hold583/X vssd1 vssd1 vccd1 vccd1 _0898_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA_fanout118_A _0613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0856__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0752_ hold701/X hold573/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1169_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0821_ _0821_/A _0821_/B vssd1 vssd1 vccd1 vccd1 _0825_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0683_ _0682_/X _0681_/X _0775_/S vssd1 vssd1 vccd1 vccd1 _0683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1304_ _1337_/CLK _1304_/D vssd1 vssd1 vccd1 vccd1 _1304_/Q sky130_fd_sc_hd__dfxtp_1
X_1235_ _1272_/CLK _1235_/D vssd1 vssd1 vccd1 vccd1 _1235_/Q sky130_fd_sc_hd__dfxtp_1
X_1166_ _1272_/CLK _1166_/D vssd1 vssd1 vccd1 vccd1 _1166_/Q sky130_fd_sc_hd__dfxtp_1
X_1097_ _1358_/CLK _1097_/D vssd1 vssd1 vccd1 vccd1 _1097_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0963__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0811__A_N _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire112 wire112/A vssd1 vssd1 vccd1 vccd1 wire112/X sky130_fd_sc_hd__clkbuf_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1020_ hold648/X hold18/X _1024_/S vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__mux2_1
XANTENNA__0783__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0804_ hold399/X hold453/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0804_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold715 _1308_/Q vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 wbs_we_i vssd1 vssd1 vccd1 vccd1 input68/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0735_ _0734_/X _0733_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0735_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0958__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0666_ hold372/X _1312_/Q hold214/X hold208/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0666_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0597_ hold36/X hold463/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0597_/X sky130_fd_sc_hd__mux2_1
X_1149_ _1351_/CLK _1149_/D vssd1 vssd1 vccd1 vccd1 _1149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1218_ _1254_/CLK _1218_/D vssd1 vssd1 vccd1 vccd1 _1218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1029__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0778__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0520_ _1044_/Q _1043_/Q _0944_/C vssd1 vssd1 vccd1 vccd1 _0521_/S sky130_fd_sc_hd__nor3b_4
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1003_ hold402/X hold517/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1003_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold501 _1106_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold545 _1098_/Q vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _0924_/X vssd1 vssd1 vccd1 vccd1 _1256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _1023_/X vssd1 vssd1 vccd1 vccd1 _1353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _1285_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0718_ hold415/X hold370/X hold421/X hold682/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0718_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_25_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold567 hold718/X vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold556 input16/X vssd1 vssd1 vccd1 vccd1 _0832_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold578 _0906_/Y vssd1 vssd1 vccd1 vccd1 _0907_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0688__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0649_ hold292/X hold271/X hold310/X hold366/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0649_/X sky130_fd_sc_hd__mux4_1
Xhold589 hold720/X vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__buf_1
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput87 _1236_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput76 _1226_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput98 _1217_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XANTENNA__0598__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1328__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0971__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold353 _1051_/Q vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _0802_/X vssd1 vssd1 vccd1 vccd1 _1200_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _1041_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _0589_/X vssd1 vssd1 vccd1 vccd1 _1086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _0585_/X vssd1 vssd1 vccd1 vccd1 _1082_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold320 _0956_/X vssd1 vssd1 vccd1 vccd1 _1287_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold331 _0569_/X vssd1 vssd1 vccd1 vccd1 _1067_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold364 _1090_/Q vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0791__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1150__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0983_ hold197/X hold206/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0983_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout107 _1009_/S vssd1 vssd1 vccd1 vccd1 _1008_/S sky130_fd_sc_hd__buf_8
Xfanout129 hold712/X vssd1 vssd1 vccd1 vccd1 _0757_/S1 sky130_fd_sc_hd__buf_4
Xfanout118 _0613_/S vssd1 vssd1 vccd1 vccd1 _0614_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0966__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0730__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold183 _0928_/X vssd1 vssd1 vccd1 vccd1 _1260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _1296_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _0571_/X vssd1 vssd1 vccd1 vccd1 _1069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _1055_/Q vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _0637_/X vssd1 vssd1 vccd1 vccd1 _1133_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0721__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0905__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1320_ _1353_/CLK _1320_/D vssd1 vssd1 vccd1 vccd1 _1320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0786__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1182_ _1346_/CLK _1182_/D vssd1 vssd1 vccd1 vccd1 _1182_/Q sky130_fd_sc_hd__dfxtp_1
X_1251_ _1251_/CLK _1251_/D vssd1 vssd1 vccd1 vccd1 _1251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0966_ hold10/X hold6/X _0976_/S vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__mux2_1
X_0897_ _0907_/A _0897_/B vssd1 vssd1 vccd1 vccd1 _1236_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1046__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1196__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0696__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0751_ _0750_/X _0749_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0820_ _0539_/B _0819_/Y _0825_/A vssd1 vssd1 vccd1 vccd1 _0820_/X sky130_fd_sc_hd__a21o_1
X_0682_ hold298/X hold263/X hold286/X hold252/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0682_/X sky130_fd_sc_hd__mux4_1
X_1303_ _1363_/CLK _1303_/D vssd1 vssd1 vccd1 vccd1 _1303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1096_ _1359_/CLK _1096_/D vssd1 vssd1 vccd1 vccd1 _1096_/Q sky130_fd_sc_hd__dfxtp_1
X_1234_ _1272_/CLK _1234_/D vssd1 vssd1 vccd1 vccd1 _1234_/Q sky130_fd_sc_hd__dfxtp_1
X_1165_ _1266_/CLK _1165_/D vssd1 vssd1 vccd1 vccd1 _1165_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0697__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout130_A _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0545__A _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0949_ hold214/X hold200/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1361__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0665_ hold236/X hold226/X hold232/X hold242/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0665_/X sky130_fd_sc_hd__mux4_1
X_0803_ hold402/X hold519/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold716 _1156_/Q vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
X_0734_ hold33/X hold8/X hold10/X hold645/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0734_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 _0977_/D vssd1 vssd1 vccd1 vccd1 _0532_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0596_ hold497/X hold527/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0596_/X sky130_fd_sc_hd__mux2_1
X_1079_ _1334_/CLK _1079_/D vssd1 vssd1 vccd1 vccd1 _1079_/Q sky130_fd_sc_hd__dfxtp_1
X_1148_ _1344_/CLK _1148_/D vssd1 vssd1 vccd1 vccd1 _1148_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0974__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1217_ _1251_/CLK _1217_/D vssd1 vssd1 vccd1 vccd1 _1217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ hold313/X hold315/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0794__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 _0609_/X vssd1 vssd1 vccd1 vccd1 _1106_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _0601_/X vssd1 vssd1 vccd1 vccd1 _1098_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0717_ hold411/X hold394/X hold392/X hold433/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0717_/X sky130_fd_sc_hd__mux4_1
Xhold524 _0954_/X vssd1 vssd1 vccd1 vccd1 _1285_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0969__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 _1288_/Q vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _1349_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold579 hold722/X vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__buf_1
Xhold568 _0850_/Y vssd1 vssd1 vccd1 vccd1 _0851_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _0832_/X vssd1 vssd1 vccd1 vccd1 _0836_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0648_ _0911_/A _0648_/B vssd1 vssd1 vccd1 vccd1 _0776_/S sky130_fd_sc_hd__nand2b_4
X_0579_ hold178/X hold114/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0579_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput88 _1237_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput77 _1227_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput99 _1218_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0789__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0699__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold310 _1048_/Q vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold354 _0553_/X vssd1 vssd1 vccd1 vccd1 _1051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _1300_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _0528_/X vssd1 vssd1 vccd1 vccd1 _1041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _1356_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _1255_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _1059_/Q vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold398 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 input53/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _0593_/X vssd1 vssd1 vccd1 vccd1 _1090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0892__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0982_ hold200/X hold714/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout108 _0944_/X vssd1 vssd1 vccd1 vccd1 _0961_/S sky130_fd_sc_hd__buf_8
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout119 _0564_/S vssd1 vssd1 vccd1 vccd1 _0580_/S sky130_fd_sc_hd__buf_8
XANTENNA__0982__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold162 _1340_/Q vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _1305_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _0558_/X vssd1 vssd1 vccd1 vccd1 _1056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _0965_/X vssd1 vssd1 vccd1 vccd1 _1296_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1318__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 _0557_/X vssd1 vssd1 vccd1 vccd1 _1055_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _1081_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0874__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1181_ _1343_/CLK _1181_/D vssd1 vssd1 vccd1 vccd1 _1181_/Q sky130_fd_sc_hd__dfxtp_1
X_1250_ _1344_/CLK _1250_/D vssd1 vssd1 vccd1 vccd1 _1250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0965_ hold194/X hold156/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0965_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0896_ _1236_/Q _0906_/A2 _0908_/B1 hold573/X vssd1 vssd1 vccd1 vccd1 _0896_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0856__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1290__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0750_ hold700/X hold517/X hold539/X hold519/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0750_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0681_ _1120_/Q hold290/X hold139/X hold284/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0681_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1302_ _1339_/CLK _1302_/D vssd1 vssd1 vccd1 vccd1 _1302_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0797__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1233_ _1266_/CLK _1233_/D vssd1 vssd1 vccd1 vccd1 _1233_/Q sky130_fd_sc_hd__dfxtp_1
X_1164_ _1363_/CLK _1164_/D vssd1 vssd1 vccd1 vccd1 _1164_/Q sky130_fd_sc_hd__dfxtp_1
X_1095_ _1265_/CLK _1095_/D vssd1 vssd1 vccd1 vccd1 _1095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0697__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0948_ hold368/X hold276/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0948_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout123_A _0775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0879_ _0907_/A _0879_/B vssd1 vssd1 vccd1 vccd1 _1227_/D sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0802_ hold313/X hold341/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1186__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0664_ hold699/X hold563/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1147_/D sky130_fd_sc_hd__mux2_1
Xhold717 _1170_/Q vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold706 _0532_/X vssd1 vssd1 vccd1 vccd1 _1042_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0733_ hold149/X hold118/X hold160/X hold296/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0733_/X sky130_fd_sc_hd__mux4_1
X_0595_ hold470/X hold509/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1216_ _1251_/CLK _1216_/D vssd1 vssd1 vccd1 vccd1 _1216_/Q sky130_fd_sc_hd__dfxtp_1
X_1147_ _1344_/CLK _1147_/D vssd1 vssd1 vccd1 vccd1 _1147_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0990__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1078_ _1339_/CLK _1078_/D vssd1 vssd1 vccd1 vccd1 _1078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__clkbuf_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ hold73/X hold673/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold503 _1136_/Q vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold547 _1130_/Q vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
X_0647_ hold488/X hold326/X _0647_/S vssd1 vssd1 vccd1 vccd1 _0647_/X sky130_fd_sc_hd__mux2_1
Xhold525 _1320_/Q vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _0957_/X vssd1 vssd1 vccd1 vccd1 _1288_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _1019_/X vssd1 vssd1 vccd1 vccd1 _1349_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0716_ hold672/X hold617/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1160_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold558 _0836_/X vssd1 vssd1 vccd1 vccd1 _0847_/B sky130_fd_sc_hd__buf_1
X_0578_ hold109/X hold65/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0578_/X sky130_fd_sc_hd__mux2_1
Xhold569 _1150_/Q vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0985__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput89 _1238_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput78 _1228_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0742__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold322 _0969_/X vssd1 vssd1 vccd1 vccd1 _1300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _0550_/X vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _0923_/X vssd1 vssd1 vccd1 vccd1 _1255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _0561_/X vssd1 vssd1 vccd1 vccd1 _1059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 _1119_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _1307_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _1178_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _1026_/X vssd1 vssd1 vccd1 vccd1 _1356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _1244_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 input53/X vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0733__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0886__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0981_ hold276/X hold698/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0981_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout109 _0944_/X vssd1 vssd1 vccd1 vccd1 _0976_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0868__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold163 _1010_/X vssd1 vssd1 vccd1 vccd1 _1340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _1346_/Q vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _0974_/X vssd1 vssd1 vccd1 vccd1 _1305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _0599_/X vssd1 vssd1 vccd1 vccd1 _1096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _1134_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _0584_/X vssd1 vssd1 vccd1 vccd1 _1081_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0706__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ _1343_/CLK _1180_/D vssd1 vssd1 vccd1 vccd1 _1180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0964_ hold31/X hold13/X _0976_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
X_0895_ _0907_/A _0895_/B vssd1 vssd1 vccd1 vccd1 _1235_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0993__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0680_ hold627/X hold611/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0680_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1258_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1301_ _1333_/CLK _1301_/D vssd1 vssd1 vccd1 vccd1 _1301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1232_ _1266_/CLK _1232_/D vssd1 vssd1 vccd1 vccd1 _1232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1163_ _1266_/CLK _1163_/D vssd1 vssd1 vccd1 vccd1 _1163_/Q sky130_fd_sc_hd__dfxtp_1
X_1094_ _1258_/CLK _1094_/D vssd1 vssd1 vccd1 vccd1 _1094_/Q sky130_fd_sc_hd__dfxtp_1
X_0947_ hold425/X hold335/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1308__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0988__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0878_ _1227_/Q _0906_/A2 _0878_/B1 hold617/X vssd1 vssd1 vccd1 vccd1 _0878_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA_fanout116_A _0647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ hold73/X hold97/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0601__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0663_ _0662_/X _0661_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0663_/X sky130_fd_sc_hd__mux2_1
X_0732_ hold676/X hold581/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1164_/D sky130_fd_sc_hd__mux2_1
Xhold718 _1146_/Q vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
X_0594_ hold88/X hold663/X _0614_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
Xhold707 _1044_/Q vssd1 vssd1 vccd1 vccd1 _0537_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1146_ _1344_/CLK _1146_/D vssd1 vssd1 vccd1 vccd1 _1146_/Q sky130_fd_sc_hd__dfxtp_1
X_1215_ _1251_/CLK _1215_/D vssd1 vssd1 vccd1 vccd1 _1215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1077_ _1337_/CLK _1077_/D vssd1 vssd1 vccd1 vccd1 _1077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1000_ hold45/X hold50/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold515 _1061_/Q vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold504 _0640_/X vssd1 vssd1 vccd1 vccd1 _1136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _0990_/X vssd1 vssd1 vccd1 vccd1 _1320_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0715_ _0714_/X _0713_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold537 _1257_/Q vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold548 _0634_/X vssd1 vssd1 vccd1 vccd1 _1130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0646_ hold212/X hold91/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0646_/X sky130_fd_sc_hd__mux2_1
X_0577_ hold265/X hold107/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0577_/X sky130_fd_sc_hd__mux2_1
Xhold559 _0847_/Y vssd1 vssd1 vccd1 vccd1 wire112/A sky130_fd_sc_hd__dlygate4sd3_1
X_1129_ _1358_/CLK _1129_/D vssd1 vssd1 vccd1 vccd1 _1129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1176__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 _1229_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
XFILLER_0_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_1_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0742__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1049__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 _1115_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _1207_/Q vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _0780_/X vssd1 vssd1 vccd1 vccd1 _1178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _1342_/Q vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _0912_/X vssd1 vssd1 vccd1 vccd1 _1244_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1199__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold312 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 input51/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 _0623_/X vssd1 vssd1 vccd1 vccd1 _1119_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0629_ hold543/X hold497/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0996__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 _0976_/X vssd1 vssd1 vccd1 vccd1 _1307_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0733__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0980_ hold335/X hold680/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1341__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold186 _1110_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _1016_/X vssd1 vssd1 vccd1 vccd1 _1346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 input62/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__clkbuf_2
Xhold153 _1039_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _1038_/Q vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold142 _0638_/X vssd1 vssd1 vccd1 vccd1 _1134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _1087_/Q vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _1251_/Q vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0706__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0963_ hold443/X hold409/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0894_ _1235_/Q _0906_/A2 _0908_/B1 hold589/X vssd1 vssd1 vccd1 vccd1 _0894_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0604__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1300_ _1358_/CLK _1300_/D vssd1 vssd1 vccd1 vccd1 _1300_/Q sky130_fd_sc_hd__dfxtp_1
X_1162_ _1332_/CLK _1162_/D vssd1 vssd1 vccd1 vccd1 _1162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1231_ _1266_/CLK _1231_/D vssd1 vssd1 vccd1 vccd1 _1231_/Q sky130_fd_sc_hd__dfxtp_1
X_1093_ _1321_/CLK _1093_/D vssd1 vssd1 vccd1 vccd1 _1093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0946_ hold79/X hold70/X _0961_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__mux2_1
X_0877_ _0907_/A _0877_/B vssd1 vssd1 vccd1 vccd1 _1226_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout109_A _0944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold719 _1153_/Q vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
X_0731_ _0730_/X _0729_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__mux2_1
X_0800_ hold45/X hold639/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold708 _0911_/B vssd1 vssd1 vccd1 vccd1 _0538_/B sky130_fd_sc_hd__dlygate4sd3_1
X_0662_ hold339/X hold698/X hold368/X hold302/X _0706_/S0 _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0662_/X sky130_fd_sc_hd__mux4_1
X_0593_ hold18/X hold364/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0593_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1214_ _1251_/CLK _1214_/D vssd1 vssd1 vccd1 vccd1 _1214_/Q sky130_fd_sc_hd__dfxtp_1
X_1145_ _1251_/CLK _1145_/D vssd1 vssd1 vccd1 vccd1 _1145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0853__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1076_ _1337_/CLK _1076_/D vssd1 vssd1 vccd1 vccd1 _1076_/Q sky130_fd_sc_hd__dfxtp_1
X_0929_ hold433/X hold362/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0999__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0904__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold516 _0563_/X vssd1 vssd1 vccd1 vccd1 _1061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _1093_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _0925_/X vssd1 vssd1 vccd1 vccd1 _1257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 _1072_/Q vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
X_0714_ hold376/X hold427/X hold445/X hold467/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0714_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0612__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold549 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 input30/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0645_ hold204/X hold114/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0645_/X sky130_fd_sc_hd__mux2_1
X_0576_ hold482/X hold399/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0576_/X sky130_fd_sc_hd__mux2_1
X_1128_ _1363_/CLK _1128_/D vssd1 vssd1 vccd1 vccd1 _1128_/Q sky130_fd_sc_hd__dfxtp_1
X_1059_ _1351_/CLK _1059_/D vssd1 vssd1 vccd1 vccd1 _1059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0522__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput69 _1243_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1120__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0607__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 _0619_/X vssd1 vssd1 vccd1 vccd1 _1115_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0628_ hold490/X hold470/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0628_/X sky130_fd_sc_hd__mux2_1
Xhold302 _1179_/Q vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _1279_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _0809_/X vssd1 vssd1 vccd1 vccd1 _1207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _1012_/X vssd1 vssd1 vccd1 vccd1 _1342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _1271_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 input51/X vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__buf_2
XFILLER_0_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold335 input57/X vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__buf_2
X_0559_ hold273/X hold259/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0559_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0886__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0868__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0861__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _0578_/X vssd1 vssd1 vccd1 vccd1 _1076_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _0783_/X vssd1 vssd1 vccd1 vccd1 _1181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _0613_/X vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _1176_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _1276_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _0525_/X vssd1 vssd1 vccd1 vccd1 _1038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _0526_/X vssd1 vssd1 vccd1 vccd1 _1039_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0800__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 _0590_/X vssd1 vssd1 vccd1 vccd1 _1087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _0919_/X vssd1 vssd1 vccd1 vccd1 _1251_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ hold421/X hold362/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0893_ _0907_/A _0893_/B vssd1 vssd1 vccd1 vccd1 _1234_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0620__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1331__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1092_ _1321_/CLK _1092_/D vssd1 vssd1 vccd1 vccd1 _1092_/Q sky130_fd_sc_hd__dfxtp_1
X_1161_ _1332_/CLK _1161_/D vssd1 vssd1 vccd1 vccd1 _1161_/Q sky130_fd_sc_hd__dfxtp_1
X_1230_ _1266_/CLK _1230_/D vssd1 vssd1 vccd1 vccd1 _1230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0945_ hold143/X hold134/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0945_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0876_ _1226_/Q _0906_/A2 _0878_/B1 hold619/X vssd1 vssd1 vccd1 vccd1 _0876_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1354__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ _1359_/CLK hold23/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0525__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0661_ hold323/X hold282/X hold353/X hold406/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0661_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0730_ hold202/X hold166/X hold194/X hold675/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0730_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 _0538_/X vssd1 vssd1 vccd1 vccd1 _1044_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0592_ hold259/X hold480/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1213_ _1251_/CLK _1213_/D vssd1 vssd1 vccd1 vccd1 _1213_/Q sky130_fd_sc_hd__dfxtp_1
X_1075_ _1332_/CLK _1075_/D vssd1 vssd1 vccd1 vccd1 _1075_/Q sky130_fd_sc_hd__dfxtp_1
X_1144_ _1346_/CLK _1144_/D vssd1 vssd1 vccd1 vccd1 _1144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout121_A _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ hold182/X hold129/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0928_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0859_ _0977_/C _0859_/B vssd1 vssd1 vccd1 vccd1 _1217_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkbuf_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0754__S0 _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold528 _0596_/X vssd1 vssd1 vccd1 vccd1 _1093_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 _1333_/Q vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _1301_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 _0574_/X vssd1 vssd1 vccd1 vccd1 _1072_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0713_ hold192/X hold671/X hold180/X hold182/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0713_/X sky130_fd_sc_hd__mux4_1
X_0644_ hold111/X hold65/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0644_/X sky130_fd_sc_hd__mux2_1
X_0575_ hold455/X hold402/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0575_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0898__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0745__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1058_ _1254_/CLK _1058_/D vssd1 vssd1 vccd1 vccd1 _1058_/Q sky130_fd_sc_hd__dfxtp_1
X_1127_ _1265_/CLK _1127_/D vssd1 vssd1 vccd1 vccd1 _1127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0803__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0623__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold303 _0781_/X vssd1 vssd1 vccd1 vccd1 _1179_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _0948_/X vssd1 vssd1 vccd1 vccd1 _1279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _0521_/X vssd1 vssd1 vccd1 vccd1 _1034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _0980_/X vssd1 vssd1 vccd1 vccd1 _1310_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _0939_/X vssd1 vssd1 vccd1 vccd1 _1271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0627_ hold168/X hold88/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0627_/X sky130_fd_sc_hd__mux2_1
X_0558_ hold139/X hold104/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0558_/X sky130_fd_sc_hd__mux2_1
Xhold325 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0859__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold347 _1095_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0718__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0708__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0709__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0618__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 _1206_/Q vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 _0975_/X vssd1 vssd1 vccd1 vccd1 _1306_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _0945_/X vssd1 vssd1 vccd1 vccd1 _1276_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold133 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 _1140_/Q vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 _0778_/X vssd1 vssd1 vccd1 vccd1 _1176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _1338_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _1328_/Q vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0528__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1260__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0961_ hold445/X hold129/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__mux2_1
X_0892_ _1234_/Q _0906_/A2 _0908_/B1 hold591/X vssd1 vssd1 vccd1 vccd1 _0892_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1283__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _1359_/CLK _1160_/D vssd1 vssd1 vccd1 vccd1 _1160_/Q sky130_fd_sc_hd__dfxtp_1
X_1091_ _1359_/CLK hold89/X vssd1 vssd1 vccd1 vccd1 _1091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0944_ _1044_/Q _1043_/Q _0944_/C vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__and3b_2
X_0875_ _0977_/C _0875_/B vssd1 vssd1 vccd1 vccd1 _1225_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0631__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1358_ _1358_/CLK _1358_/D vssd1 vssd1 vccd1 vccd1 _1358_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0867__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1289_ _1321_/CLK _1289_/D vssd1 vssd1 vccd1 vccd1 _1289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0806__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0716__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0660_ hold681/X hold567/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1146_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0591_ hold104/X hold290/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0591_/X sky130_fd_sc_hd__mux2_1
X_1212_ _1251_/CLK _1212_/D vssd1 vssd1 vccd1 vccd1 _1212_/Q sky130_fd_sc_hd__dfxtp_1
X_1074_ _1334_/CLK _1074_/D vssd1 vssd1 vccd1 vccd1 _1074_/Q sky130_fd_sc_hd__dfxtp_1
X_1143_ _1334_/CLK _1143_/D vssd1 vssd1 vccd1 vccd1 _1143_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0626__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ hold382/X hold25/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0789_ hold88/X hold308/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0789_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout114_A _0809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0858_ _1217_/Q _0847_/D _0878_/B1 hold569/X vssd1 vssd1 vccd1 vccd1 _0858_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__0904__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0754__S1 _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold507 _1270_/Q vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _1003_/X vssd1 vssd1 vccd1 vccd1 _1333_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0574_ hold505/X hold313/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0574_/X sky130_fd_sc_hd__mux2_1
Xhold529 _1321_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_0643_ hold267/X hold107/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0643_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0690__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0712_ hold637/X hold619/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0712_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0745__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1332_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1126_ _1258_/CLK _1126_/D vssd1 vssd1 vccd1 vccd1 _1126_/Q sky130_fd_sc_hd__dfxtp_1
X_1057_ _1343_/CLK _1057_/D vssd1 vssd1 vccd1 vccd1 _1057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0681__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold315 _1332_/Q vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _1118_/Q vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 input59/X vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold359 _1054_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 _0598_/X vssd1 vssd1 vccd1 vccd1 _1095_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0557_ hold172/X hold48/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0557_/X sky130_fd_sc_hd__mux2_1
X_0626_ hold240/X hold18/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0626_/X sky130_fd_sc_hd__mux2_1
Xhold337 _1131_/Q vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0718__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0875__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1109_ _1337_/CLK _1109_/D vssd1 vssd1 vccd1 vccd1 _1109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0654__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0709__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0724__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0634__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 _0808_/X vssd1 vssd1 vccd1 vccd1 _1206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 _1299_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _0998_/X vssd1 vssd1 vccd1 vccd1 _1328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _1303_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold156 input47/X vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__clkbuf_2
Xhold112 _0644_/X vssd1 vssd1 vccd1 vccd1 _1140_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 input35/X vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__clkbuf_2
X_0609_ hold399/X hold501/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0609_/X sky130_fd_sc_hd__mux2_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0809__S _0809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 _1008_/X vssd1 vssd1 vccd1 vccd1 _1338_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _1077_/Q vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold690 _1181_/Q vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0719__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ hold40/X hold25/X _0976_/S vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_0_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0891_ _0907_/A _0891_/B vssd1 vssd1 vccd1 vccd1 _1233_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0629__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1090_ _1258_/CLK _1090_/D vssd1 vssd1 vccd1 vccd1 _1090_/Q sky130_fd_sc_hd__dfxtp_1
X_0943_ hold499/X hold326/X _0943_/S vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0912__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0874_ _1225_/Q _0847_/D _0878_/B1 hold593/X vssd1 vssd1 vccd1 vccd1 _0874_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1357_ _1358_/CLK _1357_/D vssd1 vssd1 vccd1 vccd1 _1357_/Q sky130_fd_sc_hd__dfxtp_1
X_1288_ _1353_/CLK _1288_/D vssd1 vssd1 vccd1 vccd1 _1288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0883__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0732__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1123__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0590_ hold48/X hold131/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0590_/X sky130_fd_sc_hd__mux2_1
X_1142_ _1339_/CLK _1142_/D vssd1 vssd1 vccd1 vccd1 _1142_/Q sky130_fd_sc_hd__dfxtp_1
X_1211_ _1251_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _1211_/Q sky130_fd_sc_hd__dfxtp_1
X_1073_ _1334_/CLK _1073_/D vssd1 vssd1 vccd1 vccd1 _1073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0642__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0857_ _0977_/C _0857_/B vssd1 vssd1 vccd1 vccd1 _1216_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0926_ hold441/X hold36/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout107_A _1009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ hold18/X hold20/X _0792_/S vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__mux2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0552__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1296__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0727__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 _0938_/X vssd1 vssd1 vccd1 vccd1 _1270_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0711_ _0710_/X _0709_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0711_/X sky130_fd_sc_hd__mux2_1
X_0642_ hold472/X hold399/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0642_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold519 _1201_/Q vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
X_0573_ hold250/X hold73/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0573_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0690__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0898__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1125_ _1333_/CLK _1125_/D vssd1 vssd1 vccd1 vccd1 _1125_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0637__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1056_ _1346_/CLK _1056_/D vssd1 vssd1 vccd1 vccd1 _1056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0681__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0909_ input1/X _0909_/B vssd1 vssd1 vccd1 vccd1 _1242_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0625_ hold541/X hold259/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0625_/X sky130_fd_sc_hd__mux2_1
Xhold327 _1009_/X vssd1 vssd1 vccd1 vccd1 _1339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _1002_/X vssd1 vssd1 vccd1 vccd1 _1332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 _0622_/X vssd1 vssd1 vccd1 vccd1 _1118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _1132_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0920__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold338 _0635_/X vssd1 vssd1 vccd1 vccd1 _1131_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0556_ hold359/X hold137/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0556_/X sky130_fd_sc_hd__mux2_1
X_1039_ _1337_/CLK _1039_/D vssd1 vssd1 vccd1 vccd1 _1039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0891__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1108_ _1337_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _1108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0654__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0740__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0915__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0608_ hold402/X hold439/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0608_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold102 _0968_/X vssd1 vssd1 vccd1 vccd1 _1299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _0798_/X vssd1 vssd1 vccd1 vccd1 _1196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _1123_/Q vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _0972_/X vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _0978_/X vssd1 vssd1 vccd1 vccd1 _1308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _0579_/X vssd1 vssd1 vccd1 vccd1 _1077_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _1304_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 input56/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0539_/A _0539_/B _0539_/C vssd1 vssd1 vccd1 vccd1 _0541_/C sky130_fd_sc_hd__or3_1
XFILLER_0_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0560__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 _0670_/X vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 _1310_/Q vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0735__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0890_ _1233_/Q _0906_/A2 _0908_/B1 hold603/X vssd1 vssd1 vccd1 vccd1 _0890_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0645__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0555__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0870__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0942_ hold218/X hold91/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0942_/X sky130_fd_sc_hd__mux2_1
X_0873_ _0977_/C _0873_/B vssd1 vssd1 vccd1 vccd1 _1224_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1356_ _1358_/CLK _1356_/D vssd1 vssd1 vccd1 vccd1 _1356_/Q sky130_fd_sc_hd__dfxtp_1
X_1287_ _1351_/CLK _1287_/D vssd1 vssd1 vccd1 vccd1 _1287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0852__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0766__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1072_ _1333_/CLK _1072_/D vssd1 vssd1 vccd1 vccd1 _1072_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0757__S0 _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1210_ _1346_/CLK _1210_/D vssd1 vssd1 vccd1 vccd1 _1210_/Q sky130_fd_sc_hd__dfxtp_1
X_1141_ _1337_/CLK _1141_/D vssd1 vssd1 vccd1 vccd1 _1141_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0923__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0925_ hold537/X hold497/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__mux2_1
X_0787_ hold259/X hold423/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0787_/X sky130_fd_sc_hd__mux2_1
X_0856_ _1216_/Q _0847_/D _0878_/B1 hold561/X vssd1 vssd1 vccd1 vccd1 _0856_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ _1339_/CLK _1339_/D vssd1 vssd1 vccd1 vccd1 _1339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0743__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0641_ hold465/X hold402/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0641_/X sky130_fd_sc_hd__mux2_1
Xhold509 _1092_/Q vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_0710_ hold42/X hold636/X hold40/X hold29/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0710_/X sky130_fd_sc_hd__mux4_1
X_0572_ hold269/X hold45/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0572_/X sky130_fd_sc_hd__mux2_1
X_1124_ _1321_/CLK _1124_/D vssd1 vssd1 vccd1 vccd1 _1124_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0918__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1055_ _1251_/CLK _1055_/D vssd1 vssd1 vccd1 vccd1 _1055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0839_ _0839_/A input4/X input3/X input6/X vssd1 vssd1 vccd1 vccd1 _0841_/C sky130_fd_sc_hd__or4_1
X_0908_ _1242_/Q _0843_/Y _0908_/B1 hold579/X vssd1 vssd1 vccd1 vccd1 _0908_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__0889__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0563__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1113__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold339 _1343_/Q vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 _1267_/Q vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _1100_/Q vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _1068_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
X_0624_ hold713/X hold104/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0624_/X sky130_fd_sc_hd__mux2_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0555_ hold222/X hold197/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0555_/X sky130_fd_sc_hd__mux2_1
X_1107_ _1332_/CLK _1107_/D vssd1 vssd1 vccd1 vccd1 _1107_/Q sky130_fd_sc_hd__dfxtp_1
X_1038_ _1337_/CLK _1038_/D vssd1 vssd1 vccd1 vccd1 _1038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1286__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0558__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0931__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0607_ hold313/X hold461/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0607_/X sky130_fd_sc_hd__mux2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold147 _1182_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _0627_/X vssd1 vssd1 vccd1 vccd1 _1123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _0973_/X vssd1 vssd1 vccd1 vccd1 _1304_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
X_0538_ _0911_/A _0538_/B _0538_/C vssd1 vssd1 vccd1 vccd1 _0538_/X sky130_fd_sc_hd__and3b_1
Xhold114 input56/X vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__clkbuf_2
Xhold158 _1273_/Q vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1002__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold692 _1189_/Q vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _0659_/X vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 _0675_/X vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0751__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0926__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0897__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0571__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1347__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0941_ hold158/X hold114/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0941_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0872_ _1224_/Q _0847_/D _0878_/B1 hold615/X vssd1 vssd1 vccd1 vccd1 _0872_/Y sky130_fd_sc_hd__a22oi_1
X_1355_ _1359_/CLK hold43/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1286_ _1359_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0656__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0766__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0566__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0757__S1 _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1071_ _1332_/CLK _1071_/D vssd1 vssd1 vccd1 vccd1 _1071_/Q sky130_fd_sc_hd__dfxtp_1
X_1140_ _1337_/CLK _1140_/D vssd1 vssd1 vccd1 vccd1 _1140_/Q sky130_fd_sc_hd__dfxtp_1
X_0924_ hold511/X hold470/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0924_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0786_ hold104/X hold252/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0693__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0855_ _0977_/C _0855_/B vssd1 vssd1 vccd1 vccd1 _1215_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1338_ _1339_/CLK _1338_/D vssd1 vssd1 vccd1 vccd1 _1338_/Q sky130_fd_sc_hd__dfxtp_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkbuf_2
X_1269_ _1334_/CLK _1269_/D vssd1 vssd1 vccd1 vccd1 _1269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1010__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0640_ hold503/X hold313/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0571_ hold160/X hold6/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ _1344_/CLK _1054_/D vssd1 vssd1 vccd1 vccd1 _1054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1123_ _1359_/CLK _1123_/D vssd1 vssd1 vccd1 vccd1 _1123_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0934__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0666__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0907_ _0907_/A _0907_/B vssd1 vssd1 vccd1 vccd1 _1241_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0769_ hold212/X hold186/X hold220/X hold218/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0769_/X sky130_fd_sc_hd__mux4_1
X_0838_ _0838_/A _0838_/B _0838_/C _0838_/D vssd1 vssd1 vccd1 vccd1 _0841_/B sky130_fd_sc_hd__or4_1
XANTENNA__1005__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0657__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0554_ hold232/X hold200/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0554_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 _0603_/X vssd1 vssd1 vccd1 vccd1 _1100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _0570_/X vssd1 vssd1 vccd1 vccd1 _1068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold307 _0935_/X vssd1 vssd1 vccd1 vccd1 _1267_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0623_ hold300/X hold48/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0623_/X sky130_fd_sc_hd__mux2_1
X_1106_ _1334_/CLK _1106_/D vssd1 vssd1 vccd1 vccd1 _1106_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0929__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0664__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1037_ _1339_/CLK _1037_/D vssd1 vssd1 vccd1 vccd1 _1037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0574__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 _1007_/X vssd1 vssd1 vccd1 vccd1 _1337_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _1363_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold104 input65/X vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__clkbuf_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0659__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ hold73/X hold230/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold148 _0784_/X vssd1 vssd1 vccd1 vccd1 _1182_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0537_ _0537_/A _0537_/B vssd1 vssd1 vccd1 vccd1 _0538_/C sky130_fd_sc_hd__or2_1
Xhold159 _0941_/X vssd1 vssd1 vccd1 vccd1 _1273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 input63/X vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__clkbuf_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 _1096_/Q vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 hold710/X vssd1 vssd1 vccd1 vccd1 _0775_/S sky130_fd_sc_hd__buf_4
Xhold693 _0703_/X vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _1193_/Q vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0569__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1276__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0942__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1013__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0870__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold490 _1124_/Q vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1299__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0940_ hold248/X hold65/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0871_ _0977_/C _0871_/B vssd1 vssd1 vccd1 vccd1 _1223_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0937__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1285_ _1353_/CLK _1285_/D vssd1 vssd1 vccd1 vccd1 _1285_/Q sky130_fd_sc_hd__dfxtp_1
X_1354_ _1359_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0852__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0672__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1008__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1314__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1272_/CLK _1070_/D vssd1 vssd1 vccd1 vccd1 _1070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0923_ hold332/X hold88/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0693__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0854_ _1215_/Q _0847_/D _0878_/B1 _1148_/Q vssd1 vssd1 vccd1 vccd1 _0854_/Y sky130_fd_sc_hd__a22oi_1
X_0785_ hold48/X hold626/X _0792_/S vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1268_ _1333_/CLK _1268_/D vssd1 vssd1 vccd1 vccd1 _1268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0667__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1337_ _1337_/CLK _1337_/D vssd1 vssd1 vccd1 vccd1 _1337_/Q sky130_fd_sc_hd__dfxtp_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1199_ _1363_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0577__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0570_ hold328/X hold156/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0570_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1122_ _1254_/CLK _1122_/D vssd1 vssd1 vccd1 vccd1 _1122_/Q sky130_fd_sc_hd__dfxtp_1
X_1053_ _1343_/CLK _1053_/D vssd1 vssd1 vccd1 vccd1 _1053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0666__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0950__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0837_ _0837_/A _0837_/B _0837_/C _0837_/D vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__or4_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0906_ _1241_/Q _0906_/A2 _0908_/B1 hold577/X vssd1 vssd1 vccd1 vccd1 _0906_/Y sky130_fd_sc_hd__a22oi_1
X_0699_ _0698_/X _0697_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0699_/X sky130_fd_sc_hd__mux2_1
X_0768_ hold655/X hold601/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0768_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout105_A _0776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1021__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0657__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 _1187_/Q vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0553_ hold353/X hold276/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0553_/X sky130_fd_sc_hd__mux2_1
X_0622_ hold304/X hold137/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0622_/X sky130_fd_sc_hd__mux2_1
Xhold319 _1287_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_1105_ _1334_/CLK _1105_/D vssd1 vssd1 vccd1 vccd1 _1105_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0945__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1036_ _1339_/CLK _1036_/D vssd1 vssd1 vccd1 vccd1 _1036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0680__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1182__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1016__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0590__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold105 _0624_/X vssd1 vssd1 vccd1 vccd1 _1120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _1033_/X vssd1 vssd1 vccd1 vccd1 _1363_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _0984_/X vssd1 vssd1 vccd1 vccd1 _1314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _1205_/Q vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold149 _1133_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0536_ _0537_/A _0537_/B vssd1 vssd1 vccd1 vccd1 _0911_/B sky130_fd_sc_hd__nand2_1
X_0605_ hold45/X hold246/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0605_/X sky130_fd_sc_hd__mux2_1
X_1019_ hold535/X hold259/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1019_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0675__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0882__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 _1339_/Q vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _0719_/X vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _0715_/X vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _0683_/X vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 _0692_/X vssd1 vssd1 vccd1 vccd1 _1154_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0585__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0864__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ _1042_/Q _0911_/A _0910_/D _0530_/B vssd1 vssd1 vccd1 vccd1 _0944_/C sky130_fd_sc_hd__and4bb_1
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0702__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold491 _0628_/X vssd1 vssd1 vccd1 vccd1 _1124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold480 _1089_/Q vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0769__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0870_ _1223_/Q _0847_/D _0878_/B1 hold597/X vssd1 vssd1 vccd1 vccd1 _0870_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1353_ _1353_/CLK _1353_/D vssd1 vssd1 vccd1 vccd1 _1353_/Q sky130_fd_sc_hd__dfxtp_1
X_1284_ _1351_/CLK _1284_/D vssd1 vssd1 vccd1 vccd1 _1284_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0953__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0999_ hold6/X hold8/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout135_A _0843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1024__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0853_ _0977_/C _0853_/B vssd1 vssd1 vccd1 vccd1 _1214_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0922_ hold210/X hold18/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0948__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0784_ hold137/X hold147/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1267_ _1332_/CLK _1267_/D vssd1 vssd1 vccd1 vccd1 _1267_/Q sky130_fd_sc_hd__dfxtp_1
X_1336_ _1337_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_1198_ _1363_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 _1198_/Q sky130_fd_sc_hd__dfxtp_1
Xinput1 wb_rst_i vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0683__S _0775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1019__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0593__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0768__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1052_ _1343_/CLK _1052_/D vssd1 vssd1 vccd1 vccd1 _1052_/Q sky130_fd_sc_hd__dfxtp_1
X_1121_ _1321_/CLK _1121_/D vssd1 vssd1 vccd1 vccd1 _1121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0836_ _0836_/A _0836_/B _0836_/C _0836_/D vssd1 vssd1 vccd1 vccd1 _0836_/X sky130_fd_sc_hd__or4_1
X_0905_ _0907_/A _0905_/B vssd1 vssd1 vccd1 vccd1 _1240_/D sky130_fd_sc_hd__nor2_1
X_0767_ _0766_/X _0765_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0767_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0698_ hold492/X hold525/X hold513/X hold679/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0698_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1319_ _1351_/CLK _1319_/D vssd1 vssd1 vccd1 vccd1 _1319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0588__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ hold254/X hold197/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold309 _0789_/X vssd1 vssd1 vccd1 vccd1 _1187_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0552_ hold449/X hold335/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0552_/X sky130_fd_sc_hd__mux2_1
X_1104_ _1333_/CLK _1104_/D vssd1 vssd1 vccd1 vccd1 _1104_/Q sky130_fd_sc_hd__dfxtp_1
X_1035_ _1339_/CLK _1035_/D vssd1 vssd1 vccd1 vccd1 _1035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0961__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0819_ _0911_/A _0825_/A _0819_/C _0827_/A vssd1 vssd1 vccd1 vccd1 _0819_/Y sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1032__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0781__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold139 _1056_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _0807_/X vssd1 vssd1 vccd1 vccd1 _1205_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold106 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 input54/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input42/A sky130_fd_sc_hd__dlygate4sd3_1
X_0604_ hold6/X hold118/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0604_/X sky130_fd_sc_hd__mux2_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0956__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0535_ _0533_/A _0533_/B _0534_/Y vssd1 vssd1 vccd1 vccd1 _0535_/X sky130_fd_sc_hd__o21a_1
X_1018_ hold298/X hold104/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1018_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0691__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold684 _1253_/Q vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _0775_/X vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1027__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 _1040_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _1331_/Q vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _0684_/X vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 _0739_/X vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0776__S _0776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0518_ _0817_/B vssd1 vssd1 vccd1 vccd1 _0518_/Y sky130_fd_sc_hd__inv_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0702__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0596__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 _0592_/X vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _1352_/Q vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0769__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1195__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 input38/X vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0846__A1 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1352_ _1353_/CLK _1352_/D vssd1 vssd1 vccd1 vccd1 _1352_/Q sky130_fd_sc_hd__dfxtp_1
X_1283_ _1346_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0998_ hold156/X hold166/X _1008_/S vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout128_A _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0921_ hold684/X hold259/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0921_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1210__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0783_ hold197/X hold690/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0783_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1360__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0678__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0852_ _1214_/Q _0847_/D _0878_/B1 hold563/X vssd1 vssd1 vccd1 vccd1 _0852_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1335_ _1363_/CLK _1335_/D vssd1 vssd1 vccd1 vccd1 _1335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0964__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1197_ _1363_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _1197_/Q sky130_fd_sc_hd__dfxtp_1
Xinput2 hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
X_1266_ _1266_/CLK _1266_/D vssd1 vssd1 vccd1 vccd1 _1266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0669__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0903__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1051_ _1343_/CLK _1051_/D vssd1 vssd1 vccd1 vccd1 _1051_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0784__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1120_ _1346_/CLK _1120_/D vssd1 vssd1 vccd1 vccd1 _1120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0904_ _1240_/Q _0906_/A2 _0908_/B1 hold601/X vssd1 vssd1 vccd1 vccd1 _0904_/Y sky130_fd_sc_hd__a22oi_1
X_0697_ hold490/X hold509/X hold486/X hold511/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0697_/X sky130_fd_sc_hd__mux4_1
X_0766_ hold153/X hold654/X hold151/X hold116/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0766_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0959__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0835_ _0835_/A _0835_/B input22/X vssd1 vssd1 vccd1 vccd1 _0836_/D sky130_fd_sc_hd__or3b_1
XFILLER_0_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ _1359_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0900__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1249_ _1343_/CLK _1249_/D vssd1 vssd1 vccd1 vccd1 _1249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0620_ hold236/X hold200/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0779__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0551_ hold81/X hold70/X _0564_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1034_ _1339_/CLK _1034_/D vssd1 vssd1 vccd1 vccd1 _1034_/Q sky130_fd_sc_hd__dfxtp_1
X_1103_ _1332_/CLK _1103_/D vssd1 vssd1 vccd1 vccd1 _1103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0749_ hold465/X hold439/X hold455/X hold484/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0749_/X sky130_fd_sc_hd__mux4_1
X_0818_ _0825_/B _0818_/B vssd1 vssd1 vccd1 vccd1 _0827_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout110_A wire112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0599__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ hold156/X hold317/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0603_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold118 _1101_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
X_0534_ _0911_/A _0537_/B vssd1 vssd1 vccd1 vccd1 _0534_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0810__B _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 input42/X vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__clkbuf_2
Xhold107 input54/X vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__clkbuf_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0972__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1017_ hold58/X hold48/X _1024_/S vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__mux2_1
XANTENNA__0882__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold630 _0727_/X vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold685 _1034_/Q vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _1148_/Q vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _0743_/X vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _1091_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _0771_/X vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _0740_/X vssd1 vssd1 vccd1 vccd1 _1166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0792__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0864__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0967__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ _1211_/Q vssd1 vssd1 vccd1 vccd1 _0517_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 _0581_/X vssd1 vssd1 vccd1 vccd1 _1079_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _0790_/X vssd1 vssd1 vccd1 vccd1 _1188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold482 _1074_/Q vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _1022_/X vssd1 vssd1 vccd1 vccd1 _1352_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0543__A1 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0787__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1351_ _1351_/CLK _1351_/D vssd1 vssd1 vccd1 vccd1 _1351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1282_ _1346_/CLK _1282_/D vssd1 vssd1 vccd1 vccd1 _1282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0997_ hold13/X hold629/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold290 _1088_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ hold284/X hold104/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0920_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0678__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0782_ hold200/X hold208/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0782_/X sky130_fd_sc_hd__mux2_1
X_0851_ _0911_/A _0851_/B vssd1 vssd1 vccd1 vccd1 _1213_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1334_ _1334_/CLK _1334_/D vssd1 vssd1 vccd1 vccd1 _1334_/Q sky130_fd_sc_hd__dfxtp_1
X_1265_ _1265_/CLK _1265_/D vssd1 vssd1 vccd1 vccd1 _1265_/Q sky130_fd_sc_hd__dfxtp_1
X_1196_ _1363_/CLK _1196_/D vssd1 vssd1 vccd1 vccd1 _1196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0669__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0980__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ _1344_/CLK _1050_/D vssd1 vssd1 vccd1 vccd1 _1050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0834_ _0834_/A _0834_/B _0834_/C input23/X vssd1 vssd1 vccd1 vccd1 _0836_/C sky130_fd_sc_hd__or4b_1
X_0903_ _0907_/A _0903_/B vssd1 vssd1 vccd1 vccd1 _1239_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0696_ hold664/X hold609/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1155_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0765_ hold204/X hold170/X hold178/X hold158/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0765_/X sky130_fd_sc_hd__mux4_1
X_1248_ _1343_/CLK _1248_/D vssd1 vssd1 vccd1 vccd1 _1248_/Q sky130_fd_sc_hd__dfxtp_1
X_1317_ _1353_/CLK _1317_/D vssd1 vssd1 vccd1 vccd1 _1317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0975__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1179_ _1343_/CLK _1179_/D vssd1 vssd1 vccd1 vccd1 _1179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1350__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0750__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0550_ hold310/X hold134/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0550_/X sky130_fd_sc_hd__mux2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0795__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0894__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1102_ _1272_/CLK _1102_/D vssd1 vssd1 vccd1 vccd1 _1102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0741__S0 _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1033_ hold126/X hold73/X _1033_/S vssd1 vssd1 vccd1 vccd1 _1033_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0817_ _1044_/Q _0817_/B vssd1 vssd1 vccd1 vccd1 _0818_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
Xinput50 hold72/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__clkbuf_1
X_0748_ hold686/X hold589/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1168_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout103_A _0943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0679_ _0678_/X _0677_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0876__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0909__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 _1005_/X vssd1 vssd1 vccd1 vccd1 _1335_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold119 _0604_/X vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0533_ _0533_/A _0533_/B vssd1 vssd1 vccd1 vccd1 _0537_/B sky130_fd_sc_hd__and2_1
X_0602_ hold13/X hold294/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0602_/X sky130_fd_sc_hd__mux2_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0714__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1016_ hold174/X hold137/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1359_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold620 _0876_/Y vssd1 vssd1 vccd1 vccd1 _0877_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _0728_/X vssd1 vssd1 vccd1 vccd1 _1163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _0772_/X vssd1 vssd1 vccd1 vccd1 _1174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _1108_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _0747_/X vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _0668_/X vssd1 vssd1 vccd1 vccd1 _1148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _1196_/Q vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _0695_/X vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0858__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0705__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0813__A_N _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0983__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold483 _0576_/X vssd1 vssd1 vccd1 vccd1 _1074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _1138_/Q vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _1104_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _1334_/Q vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _0552_/X vssd1 vssd1 vccd1 vccd1 _1050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1091__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1281_ _1343_/CLK _1281_/D vssd1 vssd1 vccd1 vccd1 _1281_/Q sky130_fd_sc_hd__dfxtp_1
X_1350_ _1359_/CLK hold19/X vssd1 vssd1 vccd1 vccd1 _1350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0996_ hold409/X hold677/X _1008_/S vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0978__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 _1319_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _0591_/X vssd1 vssd1 vccd1 vccd1 _1088_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0850_ _1213_/Q _0847_/D _0878_/B1 hold567/X vssd1 vssd1 vccd1 vccd1 _0850_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0781_ hold276/X hold302/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0781_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0798__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1333_ _1333_/CLK _1333_/D vssd1 vssd1 vccd1 vccd1 _1333_/Q sky130_fd_sc_hd__dfxtp_1
X_1264_ _1332_/CLK _1264_/D vssd1 vssd1 vccd1 vccd1 _1264_/Q sky130_fd_sc_hd__dfxtp_1
Xinput4 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1195_ _1359_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0979_ hold70/X hold95/X _0994_/S vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__mux2_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout133_A _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0902_ _1239_/Q _0906_/A2 _0908_/B1 hold599/X vssd1 vssd1 vccd1 vccd1 _0902_/Y sky130_fd_sc_hd__a22oi_1
X_0833_ input9/X _0833_/B _0833_/C _0833_/D vssd1 vssd1 vccd1 vccd1 _0836_/B sky130_fd_sc_hd__or4_1
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0695_ _0694_/X _0693_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0695_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0764_ hold643/X hold599/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1247_ _1343_/CLK _1247_/D vssd1 vssd1 vccd1 vccd1 _1247_/Q sky130_fd_sc_hd__dfxtp_1
X_1178_ _1344_/CLK _1178_/D vssd1 vssd1 vccd1 vccd1 _1178_/Q sky130_fd_sc_hd__dfxtp_1
X_1316_ _1351_/CLK _1316_/D vssd1 vssd1 vccd1 vccd1 _1316_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0900__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0991__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0750__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1032_ hold77/X hold45/X _1033_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
X_1101_ _1266_/CLK _1101_/D vssd1 vssd1 vccd1 vccd1 _1101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0741__S1 _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0747_ _0746_/X _0745_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0816_ _0817_/B _1044_/Q vssd1 vssd1 vccd1 vccd1 _0825_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 input51/A vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput40 hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0986__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0678_ hold58/X hold60/X hold62/X hold626/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0678_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1198__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0601_ hold409/X hold545/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0601_/X sky130_fd_sc_hd__mux2_1
Xhold109 _1076_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ _0911_/A _0532_/B _0532_/C vssd1 vssd1 vccd1 vccd1 _0532_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1015_ hold478/X hold197/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1015_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0714__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 _1302_/Q vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1340__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 _0731_/X vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _1210_/Q vssd1 vssd1 vccd1 vccd1 _0539_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _1337_/Q vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _1144_/Q vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _1208_/Q vssd1 vssd1 vccd1 vccd1 _0539_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold610 _0868_/Y vssd1 vssd1 vccd1 vccd1 _0869_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold643 _0763_/X vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 _1311_/Q vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0650__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0705__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1363__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold473 _0642_/X vssd1 vssd1 vccd1 vccd1 _1138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _0608_/X vssd1 vssd1 vccd1 vccd1 _1105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _1269_/Q vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _0607_/X vssd1 vssd1 vccd1 vccd1 _1104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _1004_/X vssd1 vssd1 vccd1 vccd1 _1334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _1194_/Q vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1351_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1280_ _1343_/CLK _1280_/D vssd1 vssd1 vccd1 vccd1 _1280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ hold362/X hold370/X _1008_/S vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0994__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 _0989_/X vssd1 vssd1 vccd1 vccd1 _1319_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _1112_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _0572_/X vssd1 vssd1 vccd1 vccd1 _1070_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0780_ hold335/X hold355/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0780_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1332_ _1332_/CLK _1332_/D vssd1 vssd1 vccd1 vccd1 _1332_/Q sky130_fd_sc_hd__dfxtp_1
X_1194_ _1358_/CLK _1194_/D vssd1 vssd1 vccd1 vccd1 _1194_/Q sky130_fd_sc_hd__dfxtp_1
Xinput5 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_1263_ _1265_/CLK _1263_/D vssd1 vssd1 vccd1 vccd1 _1263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0989__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0978_ hold134/X hold715/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout126_A _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0832_ _0832_/A _0832_/B _0832_/C _0832_/D vssd1 vssd1 vccd1 vccd1 _0832_/X sky130_fd_sc_hd__or4_1
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ _0907_/A _0901_/B vssd1 vssd1 vccd1 vccd1 _1238_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0602__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0763_ _0762_/X _0761_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0763_/X sky130_fd_sc_hd__mux2_1
X_0694_ hold351/X hold280/X hold319/X hold308/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0694_/X sky130_fd_sc_hd__mux4_1
X_1315_ _1346_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1246_ _1344_/CLK _1246_/D vssd1 vssd1 vccd1 vccd1 _1246_/Q sky130_fd_sc_hd__dfxtp_1
X_1177_ _1346_/CLK hold71/X vssd1 vssd1 vccd1 vccd1 _1177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _1332_/CLK _1100_/D vssd1 vssd1 vccd1 vccd1 _1100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ hold33/X hold6/X _1033_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
XANTENNA__0894__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0746_ hold685/X hold315/X hold321/X hold341/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0746_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0815_ _0821_/B vssd1 vssd1 vccd1 vccd1 _0819_/C sky130_fd_sc_hd__inv_2
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput41 hold24/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__clkbuf_1
Xinput30 input30/A vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0677_ hold300/X hold131/X hold172/X hold164/X _0810_/B _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0677_/X sky130_fd_sc_hd__mux4_1
X_1229_ _1266_/CLK _1229_/D vssd1 vssd1 vccd1 vccd1 _1229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0876__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0600_ hold362/X hold394/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0600_/X sky130_fd_sc_hd__mux2_1
X_0531_ _0530_/B _0910_/D _1042_/Q vssd1 vssd1 vccd1 vccd1 _0532_/C sky130_fd_sc_hd__a21o_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1014_ hold372/X hold200/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold688 _0754_/X vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 _0663_/X vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _1326_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
X_0729_ hold349/X hold317/X hold328/X hold380/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0729_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0650__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 _0831_/X vssd1 vssd1 vccd1 vccd1 _1210_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0997__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 _0820_/X vssd1 vssd1 vccd1 vccd1 _1208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _0652_/X vssd1 vssd1 vccd1 vccd1 _1144_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 _0902_/Y vssd1 vssd1 vccd1 vccd1 _0903_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _1151_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _0764_/X vssd1 vssd1 vccd1 vccd1 _1172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 _0767_/X vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0858__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0700__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0610__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold474 _1085_/Q vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _0937_/X vssd1 vssd1 vccd1 vccd1 _1269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold452 _0796_/X vssd1 vssd1 vccd1 vccd1 _1194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _1258_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _1094_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _0631_/X vssd1 vssd1 vccd1 vccd1 _1127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1330__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0994_ hold129/X hold427/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0994_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0605__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold260 _0921_/X vssd1 vssd1 vccd1 vccd1 _1253_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold271 _1080_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold282 _1083_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _0616_/X vssd1 vssd1 vccd1 vccd1 _1112_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1331_ _1363_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 _1331_/Q sky130_fd_sc_hd__dfxtp_1
X_1262_ _1358_/CLK _1262_/D vssd1 vssd1 vccd1 vccd1 _1262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1193_ _1358_/CLK _1193_/D vssd1 vssd1 vccd1 vccd1 _1193_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ _1044_/Q _1043_/Q _0977_/C _0977_/D vssd1 vssd1 vccd1 vccd1 _1009_/S sky130_fd_sc_hd__or4_4
XANTENNA_fanout119_A _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0762__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0753__S0 _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0900_ _1238_/Q _0906_/A2 _0908_/B1 hold605/X vssd1 vssd1 vccd1 vccd1 _0900_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0693_ hold168/X hold663/X hold343/X hold332/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0693_/X sky130_fd_sc_hd__mux4_1
X_0831_ _0539_/C _0819_/Y _0829_/Y _0830_/X vssd1 vssd1 vccd1 vccd1 _0831_/X sky130_fd_sc_hd__a22o_1
X_0762_ hold120/X hold83/X hold124/X hold67/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0762_/X sky130_fd_sc_hd__mux4_1
X_1314_ _1346_/CLK _1314_/D vssd1 vssd1 vccd1 vccd1 _1314_/Q sky130_fd_sc_hd__dfxtp_1
X_1176_ _1346_/CLK _1176_/D vssd1 vssd1 vccd1 vccd1 _1176_/Q sky130_fd_sc_hd__dfxtp_1
X_1245_ _1251_/CLK _1245_/D vssd1 vssd1 vccd1 vccd1 _1245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0888__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0703__S _0775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0816__A_N _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1030_ hold202/X hold156/X _1033_/S vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0726__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0613__S _0613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _0834_/C sky130_fd_sc_hd__clkbuf_1
Xinput31 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _0837_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0814_ _0814_/A _1043_/Q vssd1 vssd1 vccd1 vccd1 _0821_/B sky130_fd_sc_hd__xnor2_2
X_0745_ hold503/X hold461/X hold505/X hold531/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0745_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0676_ hold670/X hold569/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1150_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput53 input53/A vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput42 input42/A vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput64 hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1228_ _1266_/CLK _1228_/D vssd1 vssd1 vccd1 vccd1 _1228_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0717__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1159_ _1266_/CLK _1159_/D vssd1 vssd1 vccd1 vccd1 _1159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0523__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ _1042_/Q _0530_/B _0910_/D vssd1 vssd1 vccd1 vccd1 _0977_/D sky130_fd_sc_hd__nand3_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0608__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1013_ hold339/X hold276/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1013_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_1_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold612 _0860_/Y vssd1 vssd1 vccd1 vccd1 _0861_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 _1173_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold689 _0755_/X vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _0723_/X vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_0659_ _0658_/X _0657_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0659_/X sky130_fd_sc_hd__mux2_1
Xhold667 _1335_/Q vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _1209_/Q vssd1 vssd1 vccd1 vccd1 _0539_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 _1197_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _1190_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
X_0728_ hold630/X hold571/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__mux2_1
Xhold656 _0768_/X vssd1 vssd1 vccd1 vccd1 _1173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold453 _1202_/Q vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _1262_/Q vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold420 _0523_/X vssd1 vssd1 vccd1 vccd1 _1036_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0801__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 _0926_/X vssd1 vssd1 vccd1 vccd1 _1258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _0588_/X vssd1 vssd1 vccd1 vccd1 _1085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _1060_/Q vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 input39/X vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__clkbuf_2
Xhold464 _0597_/X vssd1 vssd1 vccd1 vccd1 _1094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1282__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0711__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0993_ hold25/X hold636/X _0994_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0621__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1155__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0857__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold283 _0586_/X vssd1 vssd1 vccd1 vccd1 _1083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _1107_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _0583_/X vssd1 vssd1 vccd1 vccd1 _1080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 _1071_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold294 _1099_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1261_ _1358_/CLK _1261_/D vssd1 vssd1 vccd1 vccd1 _1261_/Q sky130_fd_sc_hd__dfxtp_1
X_1330_ _1363_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1192_ _1353_/CLK _1192_/D vssd1 vssd1 vccd1 vccd1 _1192_/Q sky130_fd_sc_hd__dfxtp_1
Xinput7 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ hold388/X hold326/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0616__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0526__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0762__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0753__S1 _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0830_ _0825_/D _0829_/A _0829_/B vssd1 vssd1 vccd1 vccd1 _0830_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0692_ hold649/X hold613/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0692_/X sky130_fd_sc_hd__mux2_1
X_0761_ hold111/X hold642/X hold109/X hold248/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0761_/X sky130_fd_sc_hd__mux4_1
X_1313_ _1343_/CLK _1313_/D vssd1 vssd1 vccd1 vccd1 _1313_/Q sky130_fd_sc_hd__dfxtp_1
X_1244_ _1344_/CLK _1244_/D vssd1 vssd1 vccd1 vccd1 _1244_/Q sky130_fd_sc_hd__dfxtp_1
X_1175_ _1339_/CLK _1175_/D vssd1 vssd1 vccd1 vccd1 _1175_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1251_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0959_ hold52/X hold36/X _0961_/S vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0726__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _0840_/D sky130_fd_sc_hd__clkbuf_1
Xinput54 input54/A vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
Xinput43 input43/A vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _0839_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _0834_/B sky130_fd_sc_hd__clkbuf_1
X_0813_ _0814_/A _1043_/Q vssd1 vssd1 vccd1 vccd1 _0813_/X sky130_fd_sc_hd__and2b_1
XANTENNA__0662__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0675_ _0674_/X _0673_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0675_/X sky130_fd_sc_hd__mux2_1
X_0744_ hold674/X hold591/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1167_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0717__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1227_ _1266_/CLK _1227_/D vssd1 vssd1 vccd1 vccd1 _1227_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0865__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1158_ _1258_/CLK _1158_/D vssd1 vssd1 vccd1 vccd1 _1158_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0804__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1089_ _1321_/CLK _1089_/D vssd1 vssd1 vccd1 vccd1 _1089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0653__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ hold378/X hold335/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1012_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0624__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold635 _0826_/X vssd1 vssd1 vccd1 vccd1 _1209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _1154_/Q vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold602 _0904_/Y vssd1 vssd1 vccd1 vccd1 _0905_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold624 _0707_/X vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_0727_ _0726_/X _0725_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold679 _1188_/Q vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_0658_ hold378/X hold680/X hold425/X hold355/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0658_/X sky130_fd_sc_hd__mux4_1
X_0589_ hold137/X hold374/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0589_/X sky130_fd_sc_hd__mux2_1
Xhold668 _0759_/X vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _1177_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold646 _0735_/X vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0619__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold465 _1137_/Q vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _0804_/X vssd1 vssd1 vccd1 vccd1 _1202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _0562_/X vssd1 vssd1 vccd1 vccd1 _1060_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _0930_/X vssd1 vssd1 vccd1 vccd1 _1262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _1294_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold410 _0996_/X vssd1 vssd1 vccd1 vccd1 _1326_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _1293_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _1317_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold498 _0791_/X vssd1 vssd1 vccd1 vccd1 _1189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0992_ hold36/X hold56/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0873__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold273 _1057_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold262 _0610_/X vssd1 vssd1 vccd1 vccd1 _1107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _0573_/X vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _1252_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold295 _0602_/X vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0906__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 _1122_/Q vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1359_/CLK _1260_/D vssd1 vssd1 vccd1 vccd1 _1260_/Q sky130_fd_sc_hd__dfxtp_1
X_1191_ _1359_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
Xinput8 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ hold99/X hold91/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0975_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0632__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0807__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0760_ hold668/X hold605/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1171_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1295__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0691_ _0690_/X _0689_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0691_/X sky130_fd_sc_hd__mux2_1
X_1312_ _1343_/CLK _1312_/D vssd1 vssd1 vccd1 vccd1 _1312_/Q sky130_fd_sc_hd__dfxtp_1
X_1243_ _1251_/CLK _1243_/D vssd1 vssd1 vccd1 vccd1 _1243_/Q sky130_fd_sc_hd__dfxtp_1
X_1174_ _1337_/CLK _1174_/D vssd1 vssd1 vccd1 vccd1 _1174_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0627__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0958_ hold521/X hold497/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0889_ _0907_/A _0889_/B vssd1 vssd1 vccd1 vccd1 _1232_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout124_A _0775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0888__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0743_ _0742_/X _0741_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput55 hold64/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__clkbuf_1
Xinput22 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput44 input44/A vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
Xinput11 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _0833_/C sky130_fd_sc_hd__clkbuf_1
Xinput33 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _0837_/D sky130_fd_sc_hd__clkbuf_1
X_0812_ _0821_/A _0812_/B vssd1 vssd1 vccd1 vccd1 _0825_/A sky130_fd_sc_hd__nand2_2
XANTENNA__0662__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0674_ hold174/X hold669/X hold190/X hold147/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0674_/X sky130_fd_sc_hd__mux4_1
X_1157_ _1358_/CLK _1157_/D vssd1 vssd1 vccd1 vccd1 _1157_/Q sky130_fd_sc_hd__dfxtp_1
X_1226_ _1265_/CLK _1226_/D vssd1 vssd1 vccd1 vccd1 _1226_/Q sky130_fd_sc_hd__dfxtp_1
X_1088_ _1351_/CLK _1088_/D vssd1 vssd1 vccd1 vccd1 _1088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0881__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0653__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1011_ hold85/X hold70/X _1024_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0640__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold669 _1314_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _1323_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_0726_ hold22/X hold629/X hold31/X hold15/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0726_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold614 _0866_/Y vssd1 vssd1 vccd1 vccd1 _0867_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold647 _0736_/X vssd1 vssd1 vccd1 vccd1 _1165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold603 _1166_/Q vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _0708_/X vssd1 vssd1 vccd1 vccd1 _1158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold658 _0655_/X vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_0588_ hold197/X hold474/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0588_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0657_ hold404/X hold396/X hold449/X hold390/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0657_/X sky130_fd_sc_hd__mux4_1
X_1209_ _1346_/CLK _1209_/D vssd1 vssd1 vccd1 vccd1 _1209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1206__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0550__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0635__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold455 _1073_/Q vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _0641_/X vssd1 vssd1 vccd1 vccd1 _1137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _1129_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _1261_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold488 _1143_/Q vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _1275_/Q vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _0971_/X vssd1 vssd1 vccd1 vccd1 _1302_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _0963_/X vssd1 vssd1 vccd1 vccd1 _1294_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _0962_/X vssd1 vssd1 vccd1 vccd1 _1293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _0987_/X vssd1 vssd1 vccd1 vccd1 _1317_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0709_ hold429/X hold347/X hold384/X hold382/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0709_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0991_ hold497/X hold529/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0860__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0774__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold274 _0559_/X vssd1 vssd1 vccd1 vccd1 _1057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold230 _1103_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _1316_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _1184_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _0920_/X vssd1 vssd1 vccd1 vccd1 _1252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _1265_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _0626_/X vssd1 vssd1 vccd1 vccd1 _1122_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0765__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1190_ _1359_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 _1190_/Q sky130_fd_sc_hd__dfxtp_1
Xinput9 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0974_ hold151/X hold114/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0913__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0738__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0690_ hold648/X hold38/X hold27/X hold20/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0690_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1311_ _1343_/CLK _1311_/D vssd1 vssd1 vccd1 vccd1 _1311_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0729__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1242_ _1272_/CLK _1242_/D vssd1 vssd1 vccd1 vccd1 _1242_/Q sky130_fd_sc_hd__dfxtp_1
X_1173_ _1337_/CLK _1173_/D vssd1 vssd1 vccd1 vccd1 _1173_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0643__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ hold513/X hold470/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0957_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0888_ _1232_/Q _0906_/A2 _0908_/B1 hold585/X vssd1 vssd1 vccd1 vccd1 _0888_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__0879__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout117_A _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0553__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0728__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0673_ hold304/X hold374/X hold359/X hold288/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0673_/X sky130_fd_sc_hd__mux4_1
X_0742_ hold126/X hold673/X hold101/X hold97/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0742_/X sky130_fd_sc_hd__mux4_1
Xinput67 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _0910_/B sky130_fd_sc_hd__buf_1
Xinput34 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _0910_/D sky130_fd_sc_hd__buf_2
Xinput56 input56/A vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput12 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _0833_/B sky130_fd_sc_hd__clkbuf_1
Xinput45 hold12/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__clkbuf_1
Xinput23 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
X_0811_ _0810_/B _1042_/Q vssd1 vssd1 vccd1 vccd1 _0812_/B sky130_fd_sc_hd__nand2b_1
X_1156_ _1353_/CLK _1156_/D vssd1 vssd1 vccd1 vccd1 _1156_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0638__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1225_ _1254_/CLK _1225_/D vssd1 vssd1 vccd1 vccd1 _1225_/Q sky130_fd_sc_hd__dfxtp_1
X_1087_ _1251_/CLK _1087_/D vssd1 vssd1 vccd1 vccd1 _1087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ hold162/X hold134/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0921__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold615 hold725/X vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__buf_1
Xhold648 _1350_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _1183_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold659 _0656_/X vssd1 vssd1 vccd1 vccd1 _1145_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0656_ hold658/X hold565/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0656_/X sky130_fd_sc_hd__mux2_1
Xhold604 _0890_/Y vssd1 vssd1 vccd1 vccd1 _0891_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _0711_/X vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0725_ hold337/X hold294/X hold330/X hold413/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0725_/X sky130_fd_sc_hd__mux4_1
X_0587_ hold200/X hold226/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1208_ _1346_/CLK _1208_/D vssd1 vssd1 vccd1 vccd1 _1208_/Q sky130_fd_sc_hd__dfxtp_1
X_1139_ _1339_/CLK _1139_/D vssd1 vssd1 vccd1 vccd1 _1139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0916__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0651__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _0575_/X vssd1 vssd1 vccd1 vccd1 _1073_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _0647_/X vssd1 vssd1 vccd1 vccd1 _1143_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _0633_/X vssd1 vssd1 vccd1 vccd1 _1129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _0929_/X vssd1 vssd1 vccd1 vccd1 _1261_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _1185_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _1345_/Q vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _1192_/Q vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
X_0639_ hold238/X hold73/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0639_/X sky130_fd_sc_hd__mux2_1
Xhold445 _1292_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0708_ hold624/X hold593/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0708_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0887__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1323__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0561__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0736__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0990_ hold470/X hold525/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0990_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0774__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0646__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1346__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 _1248_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold231 _0606_/X vssd1 vssd1 vccd1 vccd1 _1103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 _1078_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _0786_/X vssd1 vssd1 vccd1 vccd1 _1184_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold264 _0986_/X vssd1 vssd1 vccd1 vccd1 _1316_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _1284_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0906__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 _0933_/X vssd1 vssd1 vccd1 vccd1 _1265_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0556__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0765__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0973_ hold124/X hold65/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1000__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0738__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0674__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1310_ _1344_/CLK _1310_/D vssd1 vssd1 vccd1 vccd1 _1310_/Q sky130_fd_sc_hd__dfxtp_1
X_1241_ _1337_/CLK _1241_/D vssd1 vssd1 vccd1 vccd1 _1241_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0729__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1191__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1172_ _1272_/CLK _1172_/D vssd1 vssd1 vccd1 vccd1 _1172_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0924__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0956_ hold319/X hold88/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0956_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0665__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0887_ _0907_/A _0887_/B vssd1 vssd1 vccd1 vccd1 _1231_/D sky130_fd_sc_hd__nor2_1
Xoutput100 _1219_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
XANTENNA__0895__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1064__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0744__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _0838_/A sky130_fd_sc_hd__clkbuf_1
X_0810_ _1042_/Q _0810_/B vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__nand2b_1
X_0672_ _0671_/X hold561/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1149_/D sky130_fd_sc_hd__mux2_1
X_0741_ hold238/X hold230/X hold250/X hold306/X _0757_/S0 _0757_/S1 vssd1 vssd1 vccd1
+ vccd1 _0741_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 input68/A vssd1 vssd1 vccd1 vccd1 _0530_/B sky130_fd_sc_hd__clkbuf_2
Xinput24 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _0838_/C sky130_fd_sc_hd__clkbuf_1
Xinput46 hold69/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__clkbuf_1
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_1224_ _1254_/CLK _1224_/D vssd1 vssd1 vccd1 vccd1 _1224_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0919__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1086_ _1351_/CLK _1086_/D vssd1 vssd1 vccd1 vccd1 _1086_/Q sky130_fd_sc_hd__dfxtp_1
X_1155_ _1359_/CLK _1155_/D vssd1 vssd1 vccd1 vccd1 _1155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0939_ hold357/X hold107/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0939_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0564__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0739__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0586_ hold276/X hold282/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0586_/X sky130_fd_sc_hd__mux2_1
X_0724_ hold678/X hold595/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1162_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold616 _0872_/Y vssd1 vssd1 vccd1 vccd1 _0873_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _0712_/X vssd1 vssd1 vccd1 vccd1 _1159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 _0679_/X vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _0691_/X vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_0655_ _0654_/X _0653_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0655_/X sky130_fd_sc_hd__mux2_1
Xhold605 _1171_/Q vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
X_1207_ _1339_/CLK _1207_/D vssd1 vssd1 vccd1 vccd1 _1207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ _1334_/CLK _1138_/D vssd1 vssd1 vccd1 vccd1 _1138_/Q sky130_fd_sc_hd__dfxtp_1
X_1069_ _1266_/CLK _1069_/D vssd1 vssd1 vccd1 vccd1 _1069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0559__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1337_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0932__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold435 _1358_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _0787_/X vssd1 vssd1 vccd1 vccd1 _1185_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold402 input52/X vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__buf_2
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold413 _1263_/Q vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ _0706_/X _0705_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0707_/X sky130_fd_sc_hd__mux2_1
Xhold479 _1015_/X vssd1 vssd1 vccd1 vccd1 _1345_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _0794_/X vssd1 vssd1 vccd1 vccd1 _1192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _0961_/X vssd1 vssd1 vccd1 vccd1 _1292_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0638_ hold141/X hold45/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0638_/X sky130_fd_sc_hd__mux2_1
Xhold457 _1062_/Q vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
X_0569_ hold330/X hold13/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0569_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1003__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0752__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0860__A2 _0843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1298__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0927__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold254 _1117_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _1052_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _0916_/X vssd1 vssd1 vccd1 vccd1 _1248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _0580_/X vssd1 vssd1 vccd1 vccd1 _1078_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _1075_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _0953_/X vssd1 vssd1 vccd1 vccd1 _1284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 input60/X vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__buf_2
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold210 _1254_/Q vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold298 _1348_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0572__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0747__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ hold145/X hold107/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0972_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0567__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0674__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1171_ _1363_/CLK _1171_/D vssd1 vssd1 vccd1 vccd1 _1171_/Q sky130_fd_sc_hd__dfxtp_1
X_1240_ _1272_/CLK _1240_/D vssd1 vssd1 vccd1 vccd1 _1240_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0665__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0955_ hold27/X hold18/X _0961_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
X_0886_ _1231_/Q _0906_/A2 _0908_/B1 hold581/X vssd1 vssd1 vccd1 vccd1 _0886_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__0940__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput101 _1220_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1011__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1209__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1359__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0760__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _0835_/B sky130_fd_sc_hd__clkbuf_1
Xinput36 hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__clkbuf_1
Xinput14 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _0832_/A sky130_fd_sc_hd__clkbuf_1
X_0740_ hold640/X hold603/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__mux2_1
X_0671_ hold691/X _0669_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput47 input47/A vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__clkbuf_1
X_1154_ _1254_/CLK _1154_/D vssd1 vssd1 vccd1 vccd1 _1154_/Q sky130_fd_sc_hd__dfxtp_1
X_1223_ _1254_/CLK _1223_/D vssd1 vssd1 vccd1 vccd1 _1223_/Q sky130_fd_sc_hd__dfxtp_1
X_1085_ _1321_/CLK _1085_/D vssd1 vssd1 vccd1 vccd1 _1085_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0935__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0938_ hold507/X hold399/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0938_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout122_A _0521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0869_ _0977_/C _0869_/B vssd1 vssd1 vccd1 vccd1 _1222_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1006__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0580__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__0755__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0890__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0723_ _0722_/X _0721_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold606 _0900_/Y vssd1 vssd1 vccd1 vccd1 _0901_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold617 _1160_/Q vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
X_0585_ hold335/X hold396/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0585_/X sky130_fd_sc_hd__mux2_1
X_0654_ hold85/X hold95/X hold79/X hold657/X _0810_/B _0814_/A vssd1 vssd1 vccd1 vccd1
+ _0654_/X sky130_fd_sc_hd__mux4_1
Xhold639 _1198_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _0680_/X vssd1 vssd1 vccd1 vccd1 _1151_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1137_ _1334_/CLK _1137_/D vssd1 vssd1 vccd1 vccd1 _1137_/Q sky130_fd_sc_hd__dfxtp_1
X_1206_ _1363_/CLK _1206_/D vssd1 vssd1 vccd1 vccd1 _1206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1068_ _1332_/CLK _1068_/D vssd1 vssd1 vccd1 vccd1 _1068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0575__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0872__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0977__C _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0710__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 _1111_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold403 _0522_/X vssd1 vssd1 vccd1 vccd1 _1035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _1028_/X vssd1 vssd1 vccd1 vccd1 _1358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _1278_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0706_ hold75/X hold56/X hold52/X hold623/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0706_/X sky130_fd_sc_hd__mux4_1
Xhold458 _0564_/X vssd1 vssd1 vccd1 vccd1 _1062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold414 _0931_/X vssd1 vssd1 vccd1 vccd1 _1263_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0568_ hold437/X hold409/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0637_ hold149/X hold6/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0637_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0854__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0701__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0943__S _0943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold233 _0554_/X vssd1 vssd1 vccd1 vccd1 _1052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0621_/X vssd1 vssd1 vccd1 vccd1 _1117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _1053_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _0981_/X vssd1 vssd1 vccd1 vccd1 _1311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _0577_/X vssd1 vssd1 vccd1 vccd1 _1075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _1250_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _1018_/X vssd1 vssd1 vccd1 vccd1 _1348_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _1037_/Q vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 input61/X vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__buf_2
XFILLER_0_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _0922_/X vssd1 vssd1 vccd1 vccd1 _1254_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1014__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0763__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0971_ hold687/X hold399/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0938__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1009__S _1009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0583__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1333_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1170_ _1339_/CLK _1170_/D vssd1 vssd1 vccd1 vccd1 _1170_/Q sky130_fd_sc_hd__dfxtp_1
X_0954_ hold523/X hold259/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0954_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0885_ _0907_/A _0885_/B vssd1 vssd1 vccd1 vccd1 _1230_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0668__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1299_ _1363_/CLK _1299_/D vssd1 vssd1 vccd1 vccd1 _1299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0578__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0670_ hold478/X hold206/X hold228/X hold690/X _0757_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0670_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1303__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _0833_/D sky130_fd_sc_hd__clkbuf_1
Xinput48 hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__clkbuf_1
Xinput37 hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _0835_/A sky130_fd_sc_hd__clkbuf_1
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
X_1084_ _1343_/CLK _1084_/D vssd1 vssd1 vccd1 vccd1 _1084_/Q sky130_fd_sc_hd__dfxtp_1
X_1153_ _1351_/CLK _1153_/D vssd1 vssd1 vccd1 vccd1 _1153_/Q sky130_fd_sc_hd__dfxtp_1
X_1222_ _1254_/CLK _1222_/D vssd1 vssd1 vccd1 vccd1 _1222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0951__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0937_ hold484/X hold402/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0799_ hold6/X hold645/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__mux2_1
X_0868_ _1222_/Q _0847_/D _0878_/B1 hold609/X vssd1 vssd1 vccd1 vccd1 _0868_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA_fanout115_A _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1022__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0771__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0722_ hold435/X hold677/X hold443/X hold451/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0722_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold629 _1327_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold618 _0878_/Y vssd1 vssd1 vccd1 vccd1 _0879_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0653_ hold93/X hold184/X hold81/X hold224/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0653_/X sky130_fd_sc_hd__mux4_1
Xhold607 _1152_/Q vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
X_0584_ hold70/X hold184/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0584_/X sky130_fd_sc_hd__mux2_1
X_1136_ _1333_/CLK _1136_/D vssd1 vssd1 vccd1 vccd1 _1136_/Q sky130_fd_sc_hd__dfxtp_1
X_1205_ _1337_/CLK _1205_/D vssd1 vssd1 vccd1 vccd1 _1205_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0946__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1067_ _1265_/CLK _1067_/D vssd1 vssd1 vccd1 vccd1 _1067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1017__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0591__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0710__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold448 _0614_/X vssd1 vssd1 vccd1 vccd1 _1111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _1079_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _1066_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold415 _1357_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 _1114_/Q vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
X_0636_ hold349/X hold156/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0636_/X sky130_fd_sc_hd__mux2_1
Xhold426 _0947_/X vssd1 vssd1 vccd1 vccd1 _1278_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0705_ hold417/X hold463/X hold457/X hold441/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0705_/X sky130_fd_sc_hd__mux4_1
X_0567_ hold392/X hold362/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1171__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0676__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119_ _1254_/CLK _1119_/D vssd1 vssd1 vccd1 vccd1 _1119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0701__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0586__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 _0982_/X vssd1 vssd1 vccd1 vccd1 _1312_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold223 _0555_/X vssd1 vssd1 vccd1 vccd1 _1053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _1249_/Q vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
X_0619_ hold323/X hold276/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0619_/X sky130_fd_sc_hd__mux2_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold267 _1139_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _1142_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _0918_/X vssd1 vssd1 vccd1 vccd1 _1250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _0524_/X vssd1 vssd1 vccd1 vccd1 _1037_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _1203_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _1266_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0686__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1030__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0970_ hold539/X hold402/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0677__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0954__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1025__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0953_ hold286/X hold104/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0953_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0884_ _1230_/Q _0906_/A2 _0908_/B1 hold571/X vssd1 vssd1 vccd1 vccd1 _0884_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0949__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1298_ _1363_/CLK hold55/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__0684__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0594__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _0838_/B sky130_fd_sc_hd__clkbuf_1
Xinput49 hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__clkbuf_1
Xinput16 input16/A vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_1221_ _1254_/CLK _1221_/D vssd1 vssd1 vccd1 vccd1 _1221_/Q sky130_fd_sc_hd__dfxtp_1
X_1083_ _1343_/CLK _1083_/D vssd1 vssd1 vccd1 vccd1 _1083_/Q sky130_fd_sc_hd__dfxtp_1
X_1152_ _1258_/CLK _1152_/D vssd1 vssd1 vccd1 vccd1 _1152_/Q sky130_fd_sc_hd__dfxtp_1
X_0936_ hold531/X hold313/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0936_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1128__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0798_ hold156/X hold675/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0798_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout108_A _0944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0867_ _0977_/C _0867_/B vssd1 vssd1 vccd1 vccd1 _1221_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0679__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0589__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0890__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0721_ hold547/X hold545/X hold437/X hold431/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0721_/X sky130_fd_sc_hd__mux4_1
X_0583_ hold134/X hold271/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0583_/X sky130_fd_sc_hd__mux2_1
X_0652_ _0651_/X hold665/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0652_/X sky130_fd_sc_hd__mux2_1
Xhold608 _0862_/Y vssd1 vssd1 vccd1 vccd1 _0863_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold619 _1159_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1204_ _1337_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
X_1066_ _1358_/CLK _1066_/D vssd1 vssd1 vccd1 vccd1 _1066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0962__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1135_ _1332_/CLK _1135_/D vssd1 vssd1 vccd1 vccd1 _1135_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0919_ hold164/X hold48/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0919_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1033__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0872__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0901__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0782__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold438 _0568_/X vssd1 vssd1 vccd1 vccd1 _1066_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold416 _1027_/X vssd1 vssd1 vccd1 vccd1 _1357_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _0618_/X vssd1 vssd1 vccd1 vccd1 _1114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _1050_/Q vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_0704_ hold693/X hold615/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1157_/D sky130_fd_sc_hd__mux2_1
Xhold427 _1324_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0566_ hold180/X hold129/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0635_ hold337/X hold13/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0635_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0957__S _0961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1118_ _1344_/CLK _1118_/D vssd1 vssd1 vccd1 vccd1 _1118_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0854__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0692__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1049_ _1346_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1028__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0845__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold213 _0646_/X vssd1 vssd1 vccd1 vccd1 _1142_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold235 _0805_/X vssd1 vssd1 vccd1 vccd1 _1203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 _1360_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold224 _1245_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold257 _0917_/X vssd1 vssd1 vccd1 vccd1 _1249_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0618_ hold404/X hold335/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0618_/X sky130_fd_sc_hd__mux2_1
Xhold268 _0643_/X vssd1 vssd1 vccd1 vccd1 _1139_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0687__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 _0934_/X vssd1 vssd1 vccd1 vccd1 _1266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _1102_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_0549_ _1044_/Q _1043_/Q _0944_/C vssd1 vssd1 vccd1 vccd1 _0581_/S sky130_fd_sc_hd__and3_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0686__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0597__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0677__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0970__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout138_A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0790__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ hold62/X hold48/X _0961_/S vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0883_ _0907_/A _0883_/B vssd1 vssd1 vccd1 vccd1 _1229_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0965__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1297_ _1359_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput28 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _0837_/A sky130_fd_sc_hd__clkbuf_1
Xinput17 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _0832_/B sky130_fd_sc_hd__clkbuf_1
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
XANTENNA__0785__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1220_ _1254_/CLK _1220_/D vssd1 vssd1 vccd1 vccd1 _1220_/Q sky130_fd_sc_hd__dfxtp_1
X_1151_ _1254_/CLK _1151_/D vssd1 vssd1 vccd1 vccd1 _1151_/Q sky130_fd_sc_hd__dfxtp_1
X_1082_ _1344_/CLK _1082_/D vssd1 vssd1 vccd1 vccd1 _1082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0935_ hold306/X hold73/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0935_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0866_ _1221_/Q _0847_/D _0878_/B1 hold613/X vssd1 vssd1 vccd1 vccd1 _0866_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__0814__A _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0797_ hold13/X hold15/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
X_1349_ _1353_/CLK _1349_/D vssd1 vssd1 vccd1 vccd1 _1349_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0695__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0884__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0722__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0720_ hold683/X hold575/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1161_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0651_ _0650_/X _0649_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0651_/X sky130_fd_sc_hd__mux2_1
X_0582_ _1043_/Q _0911_/A _0977_/D _1044_/Q vssd1 vssd1 vccd1 vccd1 _0613_/S sky130_fd_sc_hd__or4b_4
Xhold609 _1155_/Q vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
X_1203_ _1332_/CLK _1203_/D vssd1 vssd1 vccd1 vccd1 _1203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0866__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1134_ _1337_/CLK _1134_/D vssd1 vssd1 vccd1 vccd1 _1134_/Q sky130_fd_sc_hd__dfxtp_1
X_1065_ _1358_/CLK _1065_/D vssd1 vssd1 vccd1 vccd1 _1065_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0713__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0544__A _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0918_ hold288/X hold137/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0918_/X sky130_fd_sc_hd__mux2_1
X_0849_ _0911_/A _0849_/B vssd1 vssd1 vccd1 vccd1 _1212_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout120_A _0581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0848__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold406 _1247_/Q vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0703_ _0702_/X _0701_/X _0775_/S vssd1 vssd1 vccd1 vccd1 _0703_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold417 _1126_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _1105_/Q vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_0634_ hold547/X hold409/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold428 _0994_/X vssd1 vssd1 vccd1 vccd1 _1324_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0565_ hold384/X hold25/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0565_/X sky130_fd_sc_hd__mux2_1
X_1117_ _1343_/CLK _1117_/D vssd1 vssd1 vccd1 vccd1 _1117_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0973__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1048_ _1344_/CLK _1048_/D vssd1 vssd1 vccd1 vccd1 _1048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0793__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold236 _1116_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold214 _1280_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 _1030_/X vssd1 vssd1 vccd1 vccd1 _1360_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _0913_/X vssd1 vssd1 vccd1 vccd1 _1245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _1070_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _0605_/X vssd1 vssd1 vccd1 vccd1 _1102_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0968__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0548_ _0518_/Y _0546_/C _0547_/Y vssd1 vssd1 vccd1 vccd1 _0548_/X sky130_fd_sc_hd__o21a_1
X_0617_ hold93/X hold70/X _0630_/S vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0907__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1306__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0788__S _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1329__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0951_ hold190/X hold137/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0951_/X sky130_fd_sc_hd__mux2_1
X_0882_ _1229_/Q _0906_/A2 _0908_/B1 hold595/X vssd1 vssd1 vccd1 vccd1 _0882_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1296_ _1363_/CLK _1296_/D vssd1 vssd1 vccd1 vccd1 _1296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0981__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _0834_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _0838_/D sky130_fd_sc_hd__clkbuf_1
X_1150_ _1346_/CLK _1150_/D vssd1 vssd1 vccd1 vccd1 _1150_/Q sky130_fd_sc_hd__dfxtp_1
X_1081_ _1251_/CLK _1081_/D vssd1 vssd1 vccd1 vccd1 _1081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0865_ _0977_/C _0865_/B vssd1 vssd1 vccd1 vccd1 _1220_/D sky130_fd_sc_hd__nor2_1
X_0934_ hold278/X hold45/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0934_/X sky130_fd_sc_hd__mux2_1
X_0796_ hold409/X hold451/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0796_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0976__S _0976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1279_ _1343_/CLK _1279_/D vssd1 vssd1 vccd1 vccd1 _1279_/Q sky130_fd_sc_hd__dfxtp_1
X_1348_ _1351_/CLK _1348_/D vssd1 vssd1 vccd1 vccd1 _1348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0722__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0581_ hold459/X hold326/X _0581_/S vssd1 vssd1 vccd1 vccd1 _0581_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0796__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0650_ hold162/X _1308_/Q hold143/X hold176/X _0810_/B _0814_/A vssd1 vssd1 vccd1
+ vccd1 _0650_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1197__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1202_ _1334_/CLK _1202_/D vssd1 vssd1 vccd1 vccd1 _1202_/Q sky130_fd_sc_hd__dfxtp_1
X_1064_ _1359_/CLK _1064_/D vssd1 vssd1 vccd1 vccd1 _1064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1133_ _1266_/CLK _1133_/D vssd1 vssd1 vccd1 vccd1 _1133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0713__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0917_ hold256/X hold197/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0917_/X sky130_fd_sc_hd__mux2_1
X_0779_ hold70/X hold657/X _0792_/S vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout113_A _0792_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0848_ _1212_/Q _0847_/D _0878_/B1 hold565/X vssd1 vssd1 vccd1 vccd1 _0848_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold407 _0915_/X vssd1 vssd1 vccd1 vccd1 _1247_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0633_ hold411/X hold362/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0633_/X sky130_fd_sc_hd__mux2_1
X_0702_ hold533/X hold529/X hold521/X hold692/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0702_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold429 _1127_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _0630_/X vssd1 vssd1 vccd1 vccd1 _1126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0564_ hold457/X hold36/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ _1343_/CLK _1116_/D vssd1 vssd1 vccd1 vccd1 _1116_/Q sky130_fd_sc_hd__dfxtp_1
X_1047_ _1251_/CLK _1047_/D vssd1 vssd1 vccd1 vccd1 _1047_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0698__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1362__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0689__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold226 _1084_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _0620_/X vssd1 vssd1 vccd1 vccd1 _1116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _0949_/X vssd1 vssd1 vccd1 vccd1 _1280_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0616_ hold292/X hold134/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0616_/X sky130_fd_sc_hd__mux2_1
Xhold259 input66/X vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__clkbuf_2
Xhold248 _1272_/Q vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _1141_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0984__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0547_ _0518_/Y _0546_/C _0911_/A vssd1 vssd1 vccd1 vccd1 _0547_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0817__B _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0979__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0902__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold590 _0894_/Y vssd1 vssd1 vccd1 vccd1 _0895_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0950_ hold228/X hold197/X _0961_/S vssd1 vssd1 vccd1 vccd1 _0950_/X sky130_fd_sc_hd__mux2_1
X_0881_ _0907_/A _0881_/B vssd1 vssd1 vccd1 vccd1 _1228_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0799__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1295_ _1359_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _0832_/D sky130_fd_sc_hd__clkbuf_1
X_1080_ _1344_/CLK _1080_/D vssd1 vssd1 vccd1 vccd1 _1080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0795_ hold362/X hold682/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0795_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0864_ _1220_/Q _0847_/D _0878_/B1 hold587/X vssd1 vssd1 vccd1 vccd1 _0864_/Y sky130_fd_sc_hd__a22oi_1
X_0933_ hold296/X hold6/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1347_ _1359_/CLK hold59/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1278_ _1344_/CLK _1278_/D vssd1 vssd1 vccd1 vccd1 _1278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0884__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0992__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _0706_/S0 vssd1 vssd1 vccd1 vccd1 _0810_/B sky130_fd_sc_hd__buf_6
X_1201_ _1333_/CLK _1201_/D vssd1 vssd1 vccd1 vccd1 _1201_/Q sky130_fd_sc_hd__dfxtp_1
X_0580_ hold220/X hold91/X _0580_/S vssd1 vssd1 vccd1 vccd1 _0580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1132_ _1332_/CLK _1132_/D vssd1 vssd1 vccd1 vccd1 _1132_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0866__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1063_ _1258_/CLK _1063_/D vssd1 vssd1 vccd1 vccd1 _1063_/Q sky130_fd_sc_hd__dfxtp_1
X_0916_ hold242/X hold200/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0987__S _0994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0778_ hold134/X hold176/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0778_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout106_A _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0847_ hold2/X _0847_/B _0847_/C _0847_/D vssd1 vssd1 vccd1 vccd1 _0847_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__1291__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0848__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1164__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0701_ hold543/X hold527/X hold515/X hold537/X _0734_/S0 _0734_/S1 vssd1 vssd1 vccd1
+ vccd1 _0701_/X sky130_fd_sc_hd__mux4_1
X_0563_ hold515/X hold497/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0563_/X sky130_fd_sc_hd__mux2_1
Xhold419 _1036_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0632_ hold192/X hold129/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0632_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input44/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0600__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1115_ _1343_/CLK _1115_/D vssd1 vssd1 vccd1 vccd1 _1115_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0698__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1046_ _1346_/CLK _1046_/D vssd1 vssd1 vccd1 vccd1 _1046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0689__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold227 _0587_/X vssd1 vssd1 vccd1 vccd1 _1084_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold238 _1135_/Q vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0541__D _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 _1058_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _0940_/X vssd1 vssd1 vccd1 vccd1 _1272_/D sky130_fd_sc_hd__dlygate4sd3_1
X_0546_ _0911_/A _0546_/B _0546_/C vssd1 vssd1 vccd1 vccd1 _1046_/D sky130_fd_sc_hd__and3b_1
X_0615_ _1043_/Q _0944_/C _1044_/Q vssd1 vssd1 vccd1 vccd1 _0647_/S sky130_fd_sc_hd__and3b_4
Xhold205 _0645_/X vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ hold22/X hold13/X _1033_/S vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0770__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0995__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _1042_/Q _0530_/B _0910_/D vssd1 vssd1 vccd1 vccd1 _0533_/B sky130_fd_sc_hd__and3_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0761__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold580 _0908_/Y vssd1 vssd1 vccd1 vccd1 _0909_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold591 _1167_/Q vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ _1228_/Q _0906_/A2 _0908_/B1 hold575/X vssd1 vssd1 vccd1 vccd1 _0880_/Y sky130_fd_sc_hd__a22oi_1
X_1363_ _1363_/CLK _1363_/D vssd1 vssd1 vccd1 vccd1 _1363_/Q sky130_fd_sc_hd__dfxtp_1
X_1294_ _1358_/CLK _1294_/D vssd1 vssd1 vccd1 vccd1 _1294_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0896__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout136_A _0843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0734__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0878__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0725__S0 _0734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0932_ hold380/X hold156/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0932_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0603__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0794_ hold129/X hold467/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0794_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0863_ _0977_/C _0863_/B vssd1 vssd1 vccd1 vccd1 _1219_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1346_ _1346_/CLK _1346_/D vssd1 vssd1 vccd1 vccd1 _1346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1277_ _1346_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout131 _0757_/S0 vssd1 vssd1 vccd1 vccd1 _0706_/S0 sky130_fd_sc_hd__buf_8
Xfanout120 _0581_/S vssd1 vssd1 vccd1 vccd1 _0564_/S sky130_fd_sc_hd__buf_8
X_1200_ _1332_/CLK _1200_/D vssd1 vssd1 vccd1 vccd1 _1200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1062_ _1258_/CLK _1062_/D vssd1 vssd1 vccd1 vccd1 _1062_/Q sky130_fd_sc_hd__dfxtp_1
X_1131_ _1265_/CLK _1131_/D vssd1 vssd1 vccd1 vccd1 _1131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0915_ hold406/X hold276/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0846_ _0847_/D hold3/X _0845_/Y vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o21a_1
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0777_ _1044_/Q _0911_/A _0977_/D _1043_/Q vssd1 vssd1 vccd1 vccd1 _0809_/S sky130_fd_sc_hd__or4b_4
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _1363_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ _0699_/X hold597/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1156_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1309__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0562_ hold486/X hold470/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 input44/X vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0631_ hold429/X hold25/X _0646_/S vssd1 vssd1 vccd1 vccd1 _0631_/X sky130_fd_sc_hd__mux2_1
X_1114_ _1344_/CLK _1114_/D vssd1 vssd1 vccd1 vccd1 _1114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1045_ _1251_/CLK _1045_/D vssd1 vssd1 vccd1 vccd1 _1045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0998__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0829_ _0829_/A _0829_/B vssd1 vssd1 vccd1 vccd1 _0829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold206 _1313_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold217 _0560_/X vssd1 vssd1 vccd1 vccd1 _1058_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0614_ hold326/X hold447/X _0614_/S vssd1 vssd1 vccd1 vccd1 _0614_/X sky130_fd_sc_hd__mux2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold228 _1281_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _0639_/X vssd1 vssd1 vccd1 vccd1 _1135_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0611__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0545_ _0814_/A _0545_/B vssd1 vssd1 vccd1 vccd1 _0546_/C sky130_fd_sc_hd__nand2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ hold435/X hold409/X _1033_/S vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0521__S _0521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1254_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0606__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0770__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0528_ hold386/X hold326/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0528_/X sky130_fd_sc_hd__mux2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1177__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0902__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0761__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold570 _0858_/Y vssd1 vssd1 vccd1 vccd1 _0859_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _0892_/Y vssd1 vssd1 vccd1 vccd1 _0893_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold581 _1164_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1293_ _1358_/CLK _1293_/D vssd1 vssd1 vccd1 vccd1 _1293_/Q sky130_fd_sc_hd__dfxtp_1
X_1362_ _1363_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
Xoutput90 _1239_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0734__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0670__S0 _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0725__S1 _0734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0862_ _1219_/Q _0847_/D _0878_/B1 hold607/X vssd1 vssd1 vccd1 vccd1 _0862_/Y sky130_fd_sc_hd__a22oi_1
X_0931_ hold413/X hold13/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0931_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0661__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0793_ hold25/X hold29/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1345_ _1353_/CLK _1345_/D vssd1 vssd1 vccd1 vccd1 _1345_/Q sky130_fd_sc_hd__dfxtp_1
X_1276_ _1346_/CLK _1276_/D vssd1 vssd1 vccd1 vccd1 _1276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0855__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout121 _1024_/S vssd1 vssd1 vccd1 vccd1 _1033_/S sky130_fd_sc_hd__buf_6
Xfanout110 wire112/X vssd1 vssd1 vccd1 vccd1 _0878_/B1 sky130_fd_sc_hd__buf_4
Xfanout132 _0757_/S0 vssd1 vssd1 vccd1 vccd1 _0774_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__0704__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1130_ _1333_/CLK _1130_/D vssd1 vssd1 vccd1 vccd1 _1130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1061_ _1321_/CLK _1061_/D vssd1 vssd1 vccd1 vccd1 _1061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0614__S _0614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0914_ hold390/X hold335/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__mux2_1
X_0845_ _0517_/Y _0847_/D _0911_/A vssd1 vssd1 vccd1 vccd1 _0845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0776_ hold695/X hold579/X _0776_/S vssd1 vssd1 vccd1 vccd1 _1175_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1328_ _1363_/CLK _1328_/D vssd1 vssd1 vccd1 vccd1 _1328_/Q sky130_fd_sc_hd__dfxtp_1
X_1259_ _1265_/CLK _1259_/D vssd1 vssd1 vccd1 vccd1 _1259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0524__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0561_ hold343/X hold88/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0561_/X sky130_fd_sc_hd__mux2_1
X_0630_ hold417/X hold36/X _0630_/S vssd1 vssd1 vccd1 vccd1 _0630_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0609__S _0612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1044_ _1251_/CLK _1044_/D vssd1 vssd1 vccd1 vccd1 _1044_/Q sky130_fd_sc_hd__dfxtp_2
X_1113_ _1346_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0759_ _0758_/X _0757_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0828_ _0825_/A _0819_/C _0827_/A _0827_/B _0825_/B vssd1 vssd1 vccd1 vccd1 _0829_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout111_A wire112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 _0983_/X vssd1 vssd1 vccd1 vccd1 _1313_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold229 _0950_/X vssd1 vssd1 vccd1 vccd1 _1281_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0613_ hold91/X hold186/X _0613_/S vssd1 vssd1 vccd1 vccd1 _0613_/X sky130_fd_sc_hd__mux2_1
Xhold218 _1274_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0544_ _0814_/A _0545_/B vssd1 vssd1 vccd1 vccd1 _0546_/B sky130_fd_sc_hd__or2_1
X_1027_ hold415/X hold362/X _1033_/S vssd1 vssd1 vccd1 vccd1 _1027_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0863__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0802__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0712__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold90 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0622__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ hold651/X hold91/X _1033_/S vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold582 _0886_/Y vssd1 vssd1 vccd1 vccd1 _0887_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _0854_/Y vssd1 vssd1 vccd1 vccd1 _0855_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _1163_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _1158_/Q vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0707__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1292_ _1353_/CLK _1292_/D vssd1 vssd1 vccd1 vccd1 _1292_/Q sky130_fd_sc_hd__dfxtp_1
X_1361_ _1363_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
Xoutput91 _1240_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_12
Xoutput80 _1230_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__0896__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1343_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__0617__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1144__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0527__S _1033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0670__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 _1246_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0878__A2 _0906_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0930_ hold431/X hold409/X _0942_/S vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1167__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0792_ hold36/X hold623/X _0792_/S vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0861_ _0977_/C _0861_/B vssd1 vssd1 vccd1 vccd1 _1218_/D sky130_fd_sc_hd__nor2_1
XANTENNA__0661__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1275_ _1334_/CLK _1275_/D vssd1 vssd1 vccd1 vccd1 _1275_/Q sky130_fd_sc_hd__dfxtp_1
X_1344_ _1344_/CLK _1344_/D vssd1 vssd1 vccd1 vccd1 _1344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0871__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout122 _0521_/S vssd1 vssd1 vccd1 vccd1 _1024_/S sky130_fd_sc_hd__buf_8
Xfanout111 wire112/X vssd1 vssd1 vccd1 vccd1 _0908_/B1 sky130_fd_sc_hd__buf_4
Xfanout133 _0757_/S0 vssd1 vssd1 vccd1 vccd1 _0734_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0720__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1060_ _1321_/CLK _1060_/D vssd1 vssd1 vccd1 vccd1 _1060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0775_ _0774_/X _0773_/X _0775_/S vssd1 vssd1 vccd1 vccd1 _0775_/X sky130_fd_sc_hd__mux2_1
X_0844_ hold2/X _1144_/Q _0910_/C vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__o21a_1
XFILLER_0_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0913_ hold224/X hold70/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0913_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0630__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1189_ _1321_/CLK _1189_/D vssd1 vssd1 vccd1 vccd1 _1189_/Q sky130_fd_sc_hd__dfxtp_1
X_1327_ _1359_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _1327_/Q sky130_fd_sc_hd__dfxtp_1
X_1258_ _1258_/CLK _1258_/D vssd1 vssd1 vccd1 vccd1 _1258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0805__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0715__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1355__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0560_ hold216/X hold18/X _0564_/S vssd1 vssd1 vccd1 vccd1 _0560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1112_ _1344_/CLK _1112_/D vssd1 vssd1 vccd1 vccd1 _1112_/Q sky130_fd_sc_hd__dfxtp_1
X_1043_ _1251_/CLK _1043_/D vssd1 vssd1 vccd1 vccd1 _1043_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_44_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0625__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ hold244/X hold667/X hold145/X hold234/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0758_/X sky130_fd_sc_hd__mux4_1
X_0827_ _0827_/A _0827_/B vssd1 vssd1 vccd1 vccd1 _0829_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout104_A _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0689_ hold240/X hold364/X hold216/X hold210/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0689_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold208 _1180_/Q vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _0942_/X vssd1 vssd1 vccd1 vccd1 _1274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0612_ hold114/X hold170/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0612_/X sky130_fd_sc_hd__mux2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0543_ _0810_/B _0648_/B _0542_/Y vssd1 vssd1 vccd1 vccd1 _1045_/D sky130_fd_sc_hd__o21a_1
XANTENNA__0773__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1026_ hold376/X hold129/X _1033_/S vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0850__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 _1168_/Q vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0526_ hold153/X hold114/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0526_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0746__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1009_ hold326/X hold694/X _1009_/S vssd1 vssd1 vccd1 vccd1 _1009_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold561 hold721/X vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__buf_1
Xhold583 hold717/X vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__buf_1
Xhold550 input30/X vssd1 vssd1 vccd1 vccd1 _0837_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _0884_/Y vssd1 vssd1 vccd1 vccd1 _0885_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _0874_/Y vssd1 vssd1 vccd1 vccd1 _0875_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0737__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0723__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1360_ _1363_/CLK _1360_/D vssd1 vssd1 vccd1 vccd1 _1360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput70 _1211_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
XANTENNA__1096__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1291_ _1359_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
Xoutput81 _1212_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput92 _1213_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_0_46_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0633__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0869__A _0977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0808__S _0808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold380 _1264_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold391 _0914_/X vssd1 vssd1 vccd1 vccd1 _1246_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0791_ hold497/X hold692/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0860_ _1218_/Q _0843_/Y _0878_/B1 hold611/X vssd1 vssd1 vccd1 vccd1 _0860_/Y sky130_fd_sc_hd__a22oi_1
X_1343_ _1343_/CLK _1343_/D vssd1 vssd1 vccd1 vccd1 _1343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0628__S _0630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1274_ _1339_/CLK _1274_/D vssd1 vssd1 vccd1 vccd1 _1274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0989_ hold88/X hold280/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0989_/X sky130_fd_sc_hd__mux2_1
Xfanout134 _1045_/Q vssd1 vssd1 vccd1 vccd1 _0757_/S0 sky130_fd_sc_hd__clkbuf_8
Xfanout123 _0775_/S vssd1 vssd1 vccd1 vccd1 _0817_/B sky130_fd_sc_hd__buf_6
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ hold366/X hold134/X _0926_/S vssd1 vssd1 vccd1 vccd1 _0912_/X sky130_fd_sc_hd__mux2_1
X_0774_ hold386/X hold694/X hold388/X hold345/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0774_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0843_ _0530_/B _0910_/D _0910_/B vssd1 vssd1 vccd1 vccd1 _0843_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1326_ _1358_/CLK _1326_/D vssd1 vssd1 vccd1 vccd1 _1326_/Q sky130_fd_sc_hd__dfxtp_1
X_1257_ _1321_/CLK _1257_/D vssd1 vssd1 vccd1 vccd1 _1257_/Q sky130_fd_sc_hd__dfxtp_1
X_1188_ _1353_/CLK _1188_/D vssd1 vssd1 vccd1 vccd1 _1188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0731__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1111_ _1334_/CLK _1111_/D vssd1 vssd1 vccd1 vccd1 _1111_/Q sky130_fd_sc_hd__dfxtp_1
X_1042_ _1251_/CLK _1042_/D vssd1 vssd1 vccd1 vccd1 _1042_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0641__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0757_ hold267/X hold261/X hold265/X hold357/X _0757_/S0 _0757_/S1 vssd1 vssd1 vccd1
+ vccd1 _0757_/X sky130_fd_sc_hd__mux4_1
X_0688_ _0687_/X hold587/X _0708_/S vssd1 vssd1 vccd1 vccd1 _1153_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0826_ _0539_/A _0819_/Y _0824_/X _0825_/Y vssd1 vssd1 vccd1 vccd1 _0826_/X sky130_fd_sc_hd__a22o_1
XANTENNA__0877__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1309_ _1346_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0551__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold209 _0782_/X vssd1 vssd1 vccd1 vccd1 _1180_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1322__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0611_ hold65/X hold642/X _0612_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
X_0542_ _0911_/A _0545_/B vssd1 vssd1 vccd1 vccd1 _0542_/Y sky130_fd_sc_hd__nor2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0773__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0847__D _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0636__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1025_ hold42/X hold25/X _1033_/S vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0809_ hold326/X hold345/X _0809_/S vssd1 vssd1 vccd1 vccd1 _0809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold721 _1149_/Q vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold710 _1047_/Q vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ hold120/X hold65/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0525_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0746__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1008_ hold91/X hold188/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1008_/X sky130_fd_sc_hd__mux2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 _0970_/X vssd1 vssd1 vccd1 vccd1 _1301_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0682__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold551 _0837_/X vssd1 vssd1 vccd1 vccd1 _0841_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _0856_/Y vssd1 vssd1 vccd1 vccd1 _0857_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold724/X vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__buf_1
Xhold595 _1162_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold584 _0898_/Y vssd1 vssd1 vccd1 vccd1 _0899_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0737__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0673__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 _1241_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
Xoutput82 _1231_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput71 _1221_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1290_ _1359_/CLK hold53/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0914__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1040__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1190__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0885__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_5_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold392 _1065_/Q vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _1325_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold381 _0932_/X vssd1 vssd1 vccd1 vccd1 _1264_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0790_ hold470/X hold679/X _0792_/S vssd1 vssd1 vccd1 vccd1 _0790_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1342_ _1344_/CLK _1342_/D vssd1 vssd1 vccd1 vccd1 _1342_/Q sky130_fd_sc_hd__dfxtp_1
X_1273_ _1337_/CLK _1273_/D vssd1 vssd1 vccd1 vccd1 _1273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout127_A _0757_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0988_ hold18/X hold38/X _0994_/S vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0644__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 _0792_/S vssd1 vssd1 vccd1 vccd1 _0808_/S sky130_fd_sc_hd__buf_8
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout102 _0926_/S vssd1 vssd1 vccd1 vccd1 _0942_/S sky130_fd_sc_hd__buf_8
Xfanout135 _0843_/Y vssd1 vssd1 vccd1 vccd1 _0847_/D sky130_fd_sc_hd__buf_4
Xfanout124 _0775_/S vssd1 vssd1 vccd1 vccd1 _0771_/S sky130_fd_sc_hd__buf_8
XANTENNA__0554__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0842_ _0847_/B _0847_/C vssd1 vssd1 vccd1 vccd1 _0842_/Y sky130_fd_sc_hd__nor2_1
X_0911_ _0911_/A _0911_/B vssd1 vssd1 vccd1 vccd1 _0943_/S sky130_fd_sc_hd__nor2_4
X_0773_ hold488/X hold447/X hold459/X hold499/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0773_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1256_ _1321_/CLK _1256_/D vssd1 vssd1 vccd1 vccd1 _1256_/Q sky130_fd_sc_hd__dfxtp_1
X_1325_ _1358_/CLK _1325_/D vssd1 vssd1 vccd1 vccd1 _1325_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0639__S _0646_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1187_ _1351_/CLK _1187_/D vssd1 vssd1 vccd1 vccd1 _1187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1110_ _1339_/CLK _1110_/D vssd1 vssd1 vccd1 vccd1 _1110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1041_ _1339_/CLK _1041_/D vssd1 vssd1 vccd1 vccd1 _1041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0825_ _0825_/A _0825_/B _0825_/C _0825_/D vssd1 vssd1 vccd1 vccd1 _0825_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0922__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0756_ hold689/X hold583/X _0772_/S vssd1 vssd1 vccd1 vccd1 _1170_/D sky130_fd_sc_hd__mux2_1
X_0687_ _0686_/X _0685_/X _0817_/B vssd1 vssd1 vccd1 vccd1 _0687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1308_ _1346_/CLK _1308_/D vssd1 vssd1 vccd1 vccd1 _1308_/Q sky130_fd_sc_hd__dfxtp_1
X_1239_ _1272_/CLK _1239_/D vssd1 vssd1 vccd1 vccd1 _1239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0893__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0908__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0610_ hold107/X hold261/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0610_/X sky130_fd_sc_hd__mux2_1
X_0541_ _0530_/B _0910_/D _0541_/C _0810_/B vssd1 vssd1 vccd1 vccd1 _0545_/B sky130_fd_sc_hd__and4b_1
XANTENNA__0917__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ hold75/X hold36/X _1024_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0652__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0850__A2 _0847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold700 _1035_/Q vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold722 _1175_/Q vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
X_0808_ hold91/X hold122/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0808_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1297__CLK _1359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 _0548_/X vssd1 vssd1 vccd1 vccd1 _1047_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0739_ _0738_/X _0737_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0562__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ hold244/X hold107/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0524_/X sky130_fd_sc_hd__mux2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0647__S _0647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1007_ hold114/X hold654/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1007_/X sky130_fd_sc_hd__mux2_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold541 _1121_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold530 _0991_/X vssd1 vssd1 vccd1 vccd1 _1321_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0682__S1 _0706_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 hold723/X vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__buf_1
Xhold552 _0841_/X vssd1 vssd1 vccd1 vccd1 _0847_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _0896_/Y vssd1 vssd1 vccd1 vccd1 _0897_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _0882_/Y vssd1 vssd1 vccd1 vccd1 _0883_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold585 _1165_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__0557__S _0564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0673__S1 _0814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 _1232_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput72 _1222_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput94 _1242_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0930__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1335__CLK _1363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1001__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 _0567_/X vssd1 vssd1 vccd1 vccd1 _1065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _0995_/X vssd1 vssd1 vccd1 vccd1 _1325_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _0556_/X vssd1 vssd1 vccd1 vccd1 _1054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _1259_/Q vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1208__CLK _1346_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1341_ _1346_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_1272_ _1272_/CLK _1272_/D vssd1 vssd1 vccd1 vccd1 _1272_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0925__S _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0987_ hold259/X hold476/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0987_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0660__S _0708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout114 _0809_/S vssd1 vssd1 vccd1 vccd1 _0792_/S sky130_fd_sc_hd__buf_8
XFILLER_0_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout136 _0843_/Y vssd1 vssd1 vccd1 vccd1 _0906_/A2 sky130_fd_sc_hd__buf_4
Xfanout103 _0943_/S vssd1 vssd1 vccd1 vccd1 _0926_/S sky130_fd_sc_hd__buf_8
Xfanout125 _0757_/S1 vssd1 vssd1 vccd1 vccd1 _0814_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0570__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold190 _1282_/Q vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0841_ _0841_/A _0841_/B _0841_/C _0841_/D vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__or4_1
X_0910_ _0911_/A _0910_/B _0910_/C _0910_/D vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__and4b_1
X_0772_ hold652/X hold577/X _0772_/S vssd1 vssd1 vccd1 vccd1 _0772_/X sky130_fd_sc_hd__mux2_1
X_1324_ _1353_/CLK _1324_/D vssd1 vssd1 vccd1 vccd1 _1324_/Q sky130_fd_sc_hd__dfxtp_1
X_1255_ _1351_/CLK _1255_/D vssd1 vssd1 vccd1 vccd1 _1255_/Q sky130_fd_sc_hd__dfxtp_1
X_1186_ _1359_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0655__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0880__B1 _0908_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0565__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ _1363_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 _1040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0862__B1 _0878_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0755_ hold688/X _0753_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0755_/X sky130_fd_sc_hd__mux2_1
X_0824_ _0825_/A _0825_/B _0825_/D _0825_/C vssd1 vssd1 vccd1 vccd1 _0824_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0686_ hold535/X hold476/X hold523/X hold423/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0686_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1307_ _1339_/CLK _1307_/D vssd1 vssd1 vccd1 vccd1 _1307_/Q sky130_fd_sc_hd__dfxtp_1
X_1169_ _1339_/CLK _1169_/D vssd1 vssd1 vccd1 vccd1 _1169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1238_ _1272_/CLK _1238_/D vssd1 vssd1 vccd1 vccd1 _1238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0758__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0540_ _0530_/B _0910_/D _0541_/C vssd1 vssd1 vccd1 vccd1 _0648_/B sky130_fd_sc_hd__and3b_1
X_1023_ hold533/X hold497/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1023_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _1358_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0933__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 _0751_/X vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold723 _1147_/Q vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
X_0738_ hold77/X hold50/X hold54/X hold639/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0738_/X sky130_fd_sc_hd__mux4_1
X_0807_ hold114/X hold116/X _0808_/S vssd1 vssd1 vccd1 vccd1 _0807_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold712 _1046_/Q vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout102_A _0926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0669_ hold254/X hold474/X hold222/X hold256/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0669_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0749__S0 _0774_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1004__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0523_ hold419/X hold399/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0523_/X sky130_fd_sc_hd__mux2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0663__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1006_ hold65/X hold83/X _1008_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0899__A _0907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 _0625_/X vssd1 vssd1 vccd1 vccd1 _1121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _1268_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold520 _0803_/X vssd1 vssd1 vccd1 vccd1 _1201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _1161_/Q vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold564 _0852_/Y vssd1 vssd1 vccd1 vccd1 _0853_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _0842_/Y vssd1 vssd1 vccd1 vccd1 _0910_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _0888_/Y vssd1 vssd1 vccd1 vccd1 _0889_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold716/X vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__buf_1
XANTENNA__0573__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0748__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 _1233_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput73 _1223_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput95 _1214_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0568__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold394 _1097_/Q vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _1344_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 _0636_/X vssd1 vssd1 vccd1 vccd1 _1132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _0927_/X vssd1 vssd1 vccd1 vccd1 _1259_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1346_/CLK _1340_/D vssd1 vssd1 vccd1 vccd1 _1340_/Q sky130_fd_sc_hd__dfxtp_1
X_1271_ _1332_/CLK _1271_/D vssd1 vssd1 vccd1 vccd1 _1271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0986_ hold104/X hold263/X _0994_/S vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0941__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _0977_/C vssd1 vssd1 vccd1 vccd1 _0911_/A sky130_fd_sc_hd__buf_4
Xfanout104 _0708_/S vssd1 vssd1 vccd1 vccd1 _0772_/S sky130_fd_sc_hd__buf_8
Xfanout126 _0757_/S1 vssd1 vssd1 vccd1 vccd1 _0706_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout115 _0630_/S vssd1 vssd1 vccd1 vccd1 _0646_/S sky130_fd_sc_hd__buf_8
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1012__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold180 _1064_/Q vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold191 _0951_/X vssd1 vssd1 vccd1 vccd1 _1282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0771_ _0770_/X _0769_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0771_/X sky130_fd_sc_hd__mux2_1
X_0840_ input5/X input8/X input7/X _0840_/D vssd1 vssd1 vccd1 vccd1 _0841_/D sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1323_ _1359_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 _1323_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0936__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1185_ _1351_/CLK _1185_/D vssd1 vssd1 vccd1 vccd1 _1185_/Q sky130_fd_sc_hd__dfxtp_1
X_1254_ _1254_/CLK _1254_/D vssd1 vssd1 vccd1 vccd1 _1254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0671__S _0817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout132_A _0757_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0969_ hold321/X hold313/X _0976_/S vssd1 vssd1 vccd1 vccd1 _0969_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1007__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0581__S _0581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0756__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0685_ hold541/X hold480/X hold273/X hold684/X _0706_/S0 _0706_/S1 vssd1 vssd1 vccd1
+ vccd1 _0685_/X sky130_fd_sc_hd__mux4_1
X_0754_ hold419/X hold494/X hold687/X hold453/X _0757_/S0 _0757_/S1 vssd1 vssd1 vccd1
+ vccd1 _0754_/X sky130_fd_sc_hd__mux4_1
X_0823_ _0827_/A _0827_/B vssd1 vssd1 vccd1 vccd1 _0825_/D sky130_fd_sc_hd__or2_1
X_1306_ _1363_/CLK _1306_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
X_1168_ _1332_/CLK _1168_/D vssd1 vssd1 vccd1 vccd1 _1168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1237_ _1272_/CLK _1237_/D vssd1 vssd1 vccd1 vccd1 _1237_/Q sky130_fd_sc_hd__dfxtp_1
X_1099_ _1265_/CLK _1099_/D vssd1 vssd1 vccd1 vccd1 _1099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0908__A2 _0843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0576__S _0580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0758__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ hold492/X hold470/X _1024_/S vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0694__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0668_ _0667_/X hold696/X _0708_/S vssd1 vssd1 vccd1 vccd1 _0668_/X sky130_fd_sc_hd__mux2_1
Xhold724 _1169_/Q vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold713 _1120_/Q vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
X_0806_ hold65/X hold67/X _0808_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold702 _1043_/Q vssd1 vssd1 vccd1 vccd1 _0533_/A sky130_fd_sc_hd__dlygate4sd3_1
X_0737_ hold141/X hold246/X hold269/X hold278/X _0774_/S0 _0774_/S1 vssd1 vssd1 vccd1
+ vccd1 _0737_/X sky130_fd_sc_hd__mux4_1
XANTENNA__0749__S1 _0774_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0599_ hold129/X hold671/X _0612_/S vssd1 vssd1 vccd1 vccd1 _0599_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0685__S0 _0706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1020__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0522_ hold700/X hold402/X _1033_/S vssd1 vssd1 vccd1 vccd1 _0522_/X sky130_fd_sc_hd__mux2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ hold107/X hold667/X _1008_/S vssd1 vssd1 vccd1 vccd1 _1005_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold510 _0595_/X vssd1 vssd1 vccd1 vccd1 _1092_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold543 _1125_/Q vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _0936_/X vssd1 vssd1 vccd1 vccd1 _1268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _1289_/Q vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 hold719/X vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold554 _0910_/X vssd1 vssd1 vccd1 vccd1 _1243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 _0870_/Y vssd1 vssd1 vccd1 vccd1 _0871_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _0880_/Y vssd1 vssd1 vccd1 vccd1 _0881_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _1145_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1015__S _1024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0658__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput85 _1234_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput74 _1224_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput96 _1215_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0764__S _0772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0649__S0 _0810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0939__S _0942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

