magic
tech sky130A
magscale 1 2
timestamp 1725878007
<< viali >>
rect 51641 27421 51675 27455
rect 52285 27285 52319 27319
rect 31493 27013 31527 27047
rect 18613 26877 18647 26911
rect 28365 26877 28399 26911
rect 28733 26877 28767 26911
rect 29285 26877 29319 26911
rect 30757 26877 30791 26911
rect 45201 26877 45235 26911
rect 46489 26877 46523 26911
rect 46673 26877 46707 26911
rect 48145 26877 48179 26911
rect 49249 26877 49283 26911
rect 50813 26877 50847 26911
rect 51089 26877 51123 26911
rect 52285 26877 52319 26911
rect 54677 26877 54711 26911
rect 45937 26809 45971 26843
rect 48697 26809 48731 26843
rect 51733 26809 51767 26843
rect 18521 26741 18555 26775
rect 19257 26741 19291 26775
rect 27813 26741 27847 26775
rect 30205 26741 30239 26775
rect 31217 26741 31251 26775
rect 45845 26741 45879 26775
rect 47317 26741 47351 26775
rect 47593 26741 47627 26775
rect 48605 26741 48639 26775
rect 50261 26741 50295 26775
rect 51641 26741 51675 26775
rect 54125 26741 54159 26775
rect 17325 26537 17359 26571
rect 47869 26537 47903 26571
rect 51549 26537 51583 26571
rect 31217 26469 31251 26503
rect 48697 26469 48731 26503
rect 53573 26469 53607 26503
rect 19257 26401 19291 26435
rect 31861 26401 31895 26435
rect 48145 26401 48179 26435
rect 49341 26401 49375 26435
rect 15393 26333 15427 26367
rect 18449 26333 18483 26367
rect 18705 26333 18739 26367
rect 19809 26333 19843 26367
rect 27905 26333 27939 26367
rect 29837 26333 29871 26367
rect 30104 26333 30138 26367
rect 45017 26333 45051 26367
rect 46489 26333 46523 26367
rect 46756 26333 46790 26367
rect 48329 26333 48363 26367
rect 50169 26333 50203 26367
rect 52193 26333 52227 26367
rect 54217 26333 54251 26367
rect 54401 26333 54435 26367
rect 15660 26265 15694 26299
rect 17141 26265 17175 26299
rect 28172 26265 28206 26299
rect 44741 26265 44775 26299
rect 45284 26265 45318 26299
rect 48789 26265 48823 26299
rect 50436 26265 50470 26299
rect 52460 26265 52494 26299
rect 53665 26265 53699 26299
rect 16773 26197 16807 26231
rect 18981 26197 19015 26231
rect 29285 26197 29319 26231
rect 31309 26197 31343 26231
rect 32229 26197 32263 26231
rect 46397 26197 46431 26231
rect 48237 26197 48271 26231
rect 51825 26197 51859 26231
rect 55045 26197 55079 26231
rect 19441 25993 19475 26027
rect 31493 25993 31527 26027
rect 44189 25993 44223 26027
rect 46029 25993 46063 26027
rect 46397 25993 46431 26027
rect 46489 25993 46523 26027
rect 46857 25993 46891 26027
rect 46949 25993 46983 26027
rect 48973 25993 49007 26027
rect 51181 25993 51215 26027
rect 52009 25993 52043 26027
rect 54125 25993 54159 26027
rect 54217 25993 54251 26027
rect 14933 25925 14967 25959
rect 15270 25925 15304 25959
rect 19073 25925 19107 25959
rect 27804 25925 27838 25959
rect 45324 25925 45358 25959
rect 50068 25925 50102 25959
rect 53012 25925 53046 25959
rect 15025 25857 15059 25891
rect 18337 25857 18371 25891
rect 18981 25857 19015 25891
rect 19809 25857 19843 25891
rect 27537 25857 27571 25891
rect 29929 25857 29963 25891
rect 30067 25857 30101 25891
rect 31125 25857 31159 25891
rect 31585 25857 31619 25891
rect 45569 25857 45603 25891
rect 45937 25857 45971 25891
rect 47593 25857 47627 25891
rect 47860 25857 47894 25891
rect 49801 25857 49835 25891
rect 51549 25857 51583 25891
rect 51641 25857 51675 25891
rect 52377 25857 52411 25891
rect 54585 25857 54619 25891
rect 7021 25789 7055 25823
rect 7757 25789 7791 25823
rect 8493 25789 8527 25823
rect 10977 25789 11011 25823
rect 13829 25789 13863 25823
rect 14381 25789 14415 25823
rect 17325 25789 17359 25823
rect 17463 25789 17497 25823
rect 17601 25789 17635 25823
rect 18521 25789 18555 25823
rect 19165 25789 19199 25823
rect 19901 25789 19935 25823
rect 20085 25789 20119 25823
rect 30205 25789 30239 25823
rect 30941 25789 30975 25823
rect 31309 25789 31343 25823
rect 32689 25789 32723 25823
rect 45753 25789 45787 25823
rect 47041 25789 47075 25823
rect 51365 25789 51399 25823
rect 52745 25789 52779 25823
rect 54677 25789 54711 25823
rect 54769 25789 54803 25823
rect 55229 25789 55263 25823
rect 11805 25721 11839 25755
rect 17877 25721 17911 25755
rect 28917 25721 28951 25755
rect 30481 25721 30515 25755
rect 31953 25721 31987 25755
rect 6469 25653 6503 25687
rect 7205 25653 7239 25687
rect 7941 25653 7975 25687
rect 8861 25653 8895 25687
rect 10425 25653 10459 25687
rect 12173 25653 12207 25687
rect 13277 25653 13311 25687
rect 16405 25653 16439 25687
rect 16681 25653 16715 25687
rect 18613 25653 18647 25687
rect 20453 25653 20487 25687
rect 29285 25653 29319 25687
rect 32137 25653 32171 25687
rect 7757 25449 7791 25483
rect 7941 25449 7975 25483
rect 10609 25449 10643 25483
rect 15209 25449 15243 25483
rect 19257 25449 19291 25483
rect 27813 25449 27847 25483
rect 31677 25449 31711 25483
rect 48237 25449 48271 25483
rect 49893 25449 49927 25483
rect 50353 25449 50387 25483
rect 54033 25449 54067 25483
rect 10517 25381 10551 25415
rect 13737 25381 13771 25415
rect 18981 25381 19015 25415
rect 27721 25381 27755 25415
rect 28641 25381 28675 25415
rect 47317 25381 47351 25415
rect 8493 25313 8527 25347
rect 11253 25313 11287 25347
rect 14105 25313 14139 25347
rect 15761 25313 15795 25347
rect 16497 25313 16531 25347
rect 16589 25313 16623 25347
rect 16865 25313 16899 25347
rect 19809 25313 19843 25347
rect 28365 25313 28399 25347
rect 29193 25313 29227 25347
rect 31585 25313 31619 25347
rect 44833 25313 44867 25347
rect 45661 25313 45695 25347
rect 47041 25313 47075 25347
rect 47777 25313 47811 25347
rect 50905 25313 50939 25347
rect 52147 25313 52181 25347
rect 52285 25313 52319 25347
rect 52561 25313 52595 25347
rect 53021 25313 53055 25347
rect 53389 25313 53423 25347
rect 54677 25313 54711 25347
rect 5549 25245 5583 25279
rect 6377 25245 6411 25279
rect 6633 25245 6667 25279
rect 9505 25245 9539 25279
rect 11437 25245 11471 25279
rect 12357 25245 12391 25279
rect 12624 25245 12658 25279
rect 15669 25245 15703 25279
rect 16405 25245 16439 25279
rect 17509 25245 17543 25279
rect 17601 25245 17635 25279
rect 26249 25245 26283 25279
rect 31329 25245 31363 25279
rect 32229 25245 32263 25279
rect 45385 25245 45419 25279
rect 46765 25245 46799 25279
rect 46903 25245 46937 25279
rect 47961 25245 47995 25279
rect 50721 25245 50755 25279
rect 52009 25245 52043 25279
rect 53205 25245 53239 25279
rect 8309 25177 8343 25211
rect 8953 25177 8987 25211
rect 10977 25177 11011 25211
rect 12081 25177 12115 25211
rect 15025 25177 15059 25211
rect 15577 25177 15611 25211
rect 17868 25177 17902 25211
rect 28181 25177 28215 25211
rect 29009 25177 29043 25211
rect 45477 25177 45511 25211
rect 53573 25177 53607 25211
rect 54125 25177 54159 25211
rect 4905 25109 4939 25143
rect 8401 25109 8435 25143
rect 11069 25109 11103 25143
rect 14749 25109 14783 25143
rect 16037 25109 16071 25143
rect 25145 25109 25179 25143
rect 25605 25109 25639 25143
rect 27261 25109 27295 25143
rect 28273 25109 28307 25143
rect 29101 25109 29135 25143
rect 30205 25109 30239 25143
rect 45017 25109 45051 25143
rect 46121 25109 46155 25143
rect 48697 25109 48731 25143
rect 50813 25109 50847 25143
rect 51365 25109 51399 25143
rect 53665 25109 53699 25143
rect 5457 24905 5491 24939
rect 6745 24905 6779 24939
rect 7113 24905 7147 24939
rect 7205 24905 7239 24939
rect 8953 24905 8987 24939
rect 11253 24905 11287 24939
rect 13829 24905 13863 24939
rect 14289 24905 14323 24939
rect 17325 24905 17359 24939
rect 18245 24905 18279 24939
rect 29837 24905 29871 24939
rect 30665 24905 30699 24939
rect 43269 24905 43303 24939
rect 45937 24905 45971 24939
rect 53205 24905 53239 24939
rect 4344 24837 4378 24871
rect 7840 24837 7874 24871
rect 10140 24837 10174 24871
rect 30573 24837 30607 24871
rect 5549 24769 5583 24803
rect 13737 24769 13771 24803
rect 14197 24769 14231 24803
rect 15025 24769 15059 24803
rect 15853 24769 15887 24803
rect 16405 24769 16439 24803
rect 16681 24769 16715 24803
rect 18797 24769 18831 24803
rect 24041 24769 24075 24803
rect 26269 24769 26303 24803
rect 26525 24769 26559 24803
rect 28457 24769 28491 24803
rect 29009 24769 29043 24803
rect 29285 24769 29319 24803
rect 42901 24769 42935 24803
rect 43913 24769 43947 24803
rect 45201 24769 45235 24803
rect 45845 24769 45879 24803
rect 46489 24769 46523 24803
rect 50353 24769 50387 24803
rect 50721 24769 50755 24803
rect 52561 24769 52595 24803
rect 4077 24701 4111 24735
rect 7389 24701 7423 24735
rect 7573 24701 7607 24735
rect 9229 24701 9263 24735
rect 9873 24701 9907 24735
rect 12541 24701 12575 24735
rect 12679 24701 12713 24735
rect 12817 24701 12851 24735
rect 13553 24701 13587 24735
rect 14381 24701 14415 24735
rect 20085 24701 20119 24735
rect 24225 24701 24259 24735
rect 26985 24701 27019 24735
rect 27537 24701 27571 24735
rect 30849 24701 30883 24735
rect 31217 24701 31251 24735
rect 42625 24701 42659 24735
rect 42809 24701 42843 24735
rect 44097 24701 44131 24735
rect 44649 24701 44683 24735
rect 13093 24633 13127 24667
rect 15393 24633 15427 24667
rect 24777 24633 24811 24667
rect 6193 24565 6227 24599
rect 11713 24565 11747 24599
rect 11897 24565 11931 24599
rect 25145 24565 25179 24599
rect 30205 24565 30239 24599
rect 42257 24565 42291 24599
rect 43361 24565 43395 24599
rect 46949 24565 46983 24599
rect 47777 24565 47811 24599
rect 51273 24565 51307 24599
rect 5457 24361 5491 24395
rect 14105 24361 14139 24395
rect 26525 24361 26559 24395
rect 41613 24361 41647 24395
rect 43821 24361 43855 24395
rect 13921 24293 13955 24327
rect 3985 24225 4019 24259
rect 5917 24225 5951 24259
rect 6101 24225 6135 24259
rect 7205 24225 7239 24259
rect 7481 24225 7515 24259
rect 7941 24225 7975 24259
rect 11989 24225 12023 24259
rect 14657 24225 14691 24259
rect 24501 24225 24535 24259
rect 5825 24157 5859 24191
rect 6929 24157 6963 24191
rect 7067 24157 7101 24191
rect 8125 24157 8159 24191
rect 9965 24157 9999 24191
rect 12541 24157 12575 24191
rect 15393 24157 15427 24191
rect 20085 24157 20119 24191
rect 20177 24157 20211 24191
rect 20913 24157 20947 24191
rect 22661 24157 22695 24191
rect 23949 24157 23983 24191
rect 25053 24157 25087 24191
rect 25237 24157 25271 24191
rect 27077 24157 27111 24191
rect 33517 24157 33551 24191
rect 33701 24157 33735 24191
rect 36001 24157 36035 24191
rect 37565 24157 37599 24191
rect 37749 24157 37783 24191
rect 40417 24157 40451 24191
rect 41153 24157 41187 24191
rect 42349 24157 42383 24191
rect 42441 24157 42475 24191
rect 42708 24157 42742 24191
rect 44005 24157 44039 24191
rect 46489 24157 46523 24191
rect 46765 24157 46799 24191
rect 48145 24157 48179 24191
rect 50997 24157 51031 24191
rect 51917 24157 51951 24191
rect 52653 24157 52687 24191
rect 53297 24157 53331 24191
rect 54401 24157 54435 24191
rect 55321 24157 55355 24191
rect 57161 24157 57195 24191
rect 57897 24157 57931 24191
rect 4252 24089 4286 24123
rect 10232 24089 10266 24123
rect 11805 24089 11839 24123
rect 12808 24089 12842 24123
rect 14841 24089 14875 24123
rect 23213 24089 23247 24123
rect 47317 24089 47351 24123
rect 5365 24021 5399 24055
rect 6285 24021 6319 24055
rect 8401 24021 8435 24055
rect 11345 24021 11379 24055
rect 11437 24021 11471 24055
rect 11897 24021 11931 24055
rect 19441 24021 19475 24055
rect 20821 24021 20855 24055
rect 21557 24021 21591 24055
rect 22109 24021 22143 24055
rect 23397 24021 23431 24055
rect 27721 24021 27755 24055
rect 32965 24021 32999 24055
rect 34345 24021 34379 24055
rect 35449 24021 35483 24055
rect 37013 24021 37047 24055
rect 38393 24021 38427 24055
rect 39681 24021 39715 24055
rect 39865 24021 39899 24055
rect 40601 24021 40635 24055
rect 41705 24021 41739 24055
rect 44649 24021 44683 24055
rect 45937 24021 45971 24055
rect 47501 24021 47535 24055
rect 50445 24021 50479 24055
rect 51273 24021 51307 24055
rect 52009 24021 52043 24055
rect 52745 24021 52779 24055
rect 53665 24021 53699 24055
rect 53849 24021 53883 24055
rect 54769 24021 54803 24055
rect 55965 24021 55999 24055
rect 56609 24021 56643 24055
rect 57345 24021 57379 24055
rect 5181 23817 5215 23851
rect 10701 23817 10735 23851
rect 13737 23817 13771 23851
rect 14105 23817 14139 23851
rect 18613 23817 18647 23851
rect 20177 23817 20211 23851
rect 20269 23817 20303 23851
rect 23581 23817 23615 23851
rect 26801 23817 26835 23851
rect 31585 23817 31619 23851
rect 33517 23817 33551 23851
rect 36645 23817 36679 23851
rect 37289 23817 37323 23851
rect 37657 23817 37691 23851
rect 40693 23817 40727 23851
rect 46029 23817 46063 23851
rect 48329 23817 48363 23851
rect 50445 23817 50479 23851
rect 52285 23817 52319 23851
rect 53849 23817 53883 23851
rect 55413 23817 55447 23851
rect 11529 23749 11563 23783
rect 14381 23749 14415 23783
rect 19064 23749 19098 23783
rect 21557 23749 21591 23783
rect 22201 23749 22235 23783
rect 31217 23749 31251 23783
rect 34520 23749 34554 23783
rect 38752 23749 38786 23783
rect 42441 23749 42475 23783
rect 44557 23749 44591 23783
rect 47869 23749 47903 23783
rect 49065 23749 49099 23783
rect 51917 23749 51951 23783
rect 54217 23749 54251 23783
rect 56600 23749 56634 23783
rect 5089 23681 5123 23715
rect 5549 23681 5583 23715
rect 11345 23681 11379 23715
rect 13645 23681 13679 23715
rect 20637 23681 20671 23715
rect 23949 23681 23983 23715
rect 24041 23681 24075 23715
rect 24777 23681 24811 23715
rect 25688 23681 25722 23715
rect 26985 23681 27019 23715
rect 32137 23681 32171 23715
rect 32404 23681 32438 23715
rect 38301 23681 38335 23715
rect 38485 23681 38519 23715
rect 40233 23681 40267 23715
rect 40325 23681 40359 23715
rect 40785 23681 40819 23715
rect 44649 23681 44683 23715
rect 46397 23681 46431 23715
rect 46489 23681 46523 23715
rect 47961 23681 47995 23715
rect 50813 23681 50847 23715
rect 50905 23681 50939 23715
rect 52929 23681 52963 23715
rect 54309 23681 54343 23715
rect 54953 23681 54987 23715
rect 55045 23681 55079 23715
rect 56149 23681 56183 23715
rect 5365 23613 5399 23647
rect 13461 23613 13495 23647
rect 15393 23613 15427 23647
rect 16405 23613 16439 23647
rect 17417 23613 17451 23647
rect 18797 23613 18831 23647
rect 20729 23613 20763 23647
rect 20821 23613 20855 23647
rect 21925 23613 21959 23647
rect 22109 23613 22143 23647
rect 22661 23613 22695 23647
rect 24133 23613 24167 23647
rect 24869 23613 24903 23647
rect 24961 23613 24995 23647
rect 25421 23613 25455 23647
rect 27629 23613 27663 23647
rect 29745 23613 29779 23647
rect 34253 23613 34287 23647
rect 36277 23613 36311 23647
rect 37749 23613 37783 23647
rect 37933 23613 37967 23647
rect 40049 23613 40083 23647
rect 41429 23613 41463 23647
rect 42073 23613 42107 23647
rect 44465 23613 44499 23647
rect 45661 23613 45695 23647
rect 46673 23613 46707 23647
rect 47041 23613 47075 23647
rect 47685 23613 47719 23647
rect 48513 23613 48547 23647
rect 50997 23613 51031 23647
rect 51641 23613 51675 23647
rect 51825 23613 51859 23647
rect 54401 23613 54435 23647
rect 54769 23613 54803 23647
rect 56333 23613 56367 23647
rect 58449 23613 58483 23647
rect 6193 23545 6227 23579
rect 22569 23545 22603 23579
rect 35633 23545 35667 23579
rect 39865 23545 39899 23579
rect 45017 23545 45051 23579
rect 49893 23545 49927 23579
rect 57713 23545 57747 23579
rect 4721 23477 4755 23511
rect 6561 23477 6595 23511
rect 8217 23477 8251 23511
rect 13001 23477 13035 23511
rect 14841 23477 14875 23511
rect 15853 23477 15887 23511
rect 16865 23477 16899 23511
rect 23305 23477 23339 23511
rect 24409 23477 24443 23511
rect 28457 23477 28491 23511
rect 30389 23477 30423 23511
rect 33885 23477 33919 23511
rect 35725 23477 35759 23511
rect 37105 23477 37139 23511
rect 41521 23477 41555 23511
rect 43913 23477 43947 23511
rect 45109 23477 45143 23511
rect 50261 23477 50295 23511
rect 53573 23477 53607 23511
rect 55505 23477 55539 23511
rect 57897 23477 57931 23511
rect 4537 23273 4571 23307
rect 5549 23273 5583 23307
rect 12265 23273 12299 23307
rect 15945 23273 15979 23307
rect 24225 23273 24259 23307
rect 25145 23273 25179 23307
rect 27077 23273 27111 23307
rect 33425 23273 33459 23307
rect 37749 23273 37783 23307
rect 39865 23273 39899 23307
rect 45293 23273 45327 23307
rect 46857 23273 46891 23307
rect 48513 23273 48547 23307
rect 51549 23273 51583 23307
rect 54861 23273 54895 23307
rect 57253 23273 57287 23307
rect 28641 23205 28675 23239
rect 39037 23205 39071 23239
rect 51641 23205 51675 23239
rect 58265 23205 58299 23239
rect 5089 23137 5123 23171
rect 11621 23137 11655 23171
rect 17325 23137 17359 23171
rect 19901 23137 19935 23171
rect 20085 23137 20119 23171
rect 20729 23137 20763 23171
rect 21189 23137 21223 23171
rect 21582 23137 21616 23171
rect 22845 23137 22879 23171
rect 24961 23137 24995 23171
rect 26065 23137 26099 23171
rect 26341 23137 26375 23171
rect 26801 23137 26835 23171
rect 27629 23137 27663 23171
rect 28549 23137 28583 23171
rect 29193 23137 29227 23171
rect 30665 23137 30699 23171
rect 30757 23137 30791 23171
rect 34069 23137 34103 23171
rect 38485 23137 38519 23171
rect 38644 23137 38678 23171
rect 39497 23137 39531 23171
rect 40417 23137 40451 23171
rect 42717 23137 42751 23171
rect 42901 23137 42935 23171
rect 43361 23137 43395 23171
rect 43913 23137 43947 23171
rect 56103 23137 56137 23171
rect 56241 23137 56275 23171
rect 56517 23137 56551 23171
rect 57805 23137 57839 23171
rect 13553 23069 13587 23103
rect 14473 23069 14507 23103
rect 17969 23069 18003 23103
rect 18521 23069 18555 23103
rect 20545 23069 20579 23103
rect 21465 23069 21499 23103
rect 21741 23069 21775 23103
rect 22661 23069 22695 23103
rect 23112 23069 23146 23103
rect 25789 23069 25823 23103
rect 25927 23069 25961 23103
rect 26985 23069 27019 23103
rect 27445 23069 27479 23103
rect 31585 23069 31619 23103
rect 31953 23069 31987 23103
rect 33793 23069 33827 23103
rect 34713 23069 34747 23103
rect 36369 23069 36403 23103
rect 38761 23069 38795 23103
rect 39681 23069 39715 23103
rect 41245 23069 41279 23103
rect 43637 23069 43671 23103
rect 43754 23069 43788 23103
rect 45477 23069 45511 23103
rect 47133 23069 47167 23103
rect 47400 23069 47434 23103
rect 50169 23069 50203 23103
rect 53021 23069 53055 23103
rect 53481 23069 53515 23103
rect 55965 23069 55999 23103
rect 56977 23069 57011 23103
rect 57161 23069 57195 23103
rect 57713 23069 57747 23103
rect 12909 23001 12943 23035
rect 14740 23001 14774 23035
rect 17058 23001 17092 23035
rect 19809 23001 19843 23035
rect 29101 23001 29135 23035
rect 32220 23001 32254 23035
rect 34980 23001 35014 23035
rect 36636 23001 36670 23035
rect 40233 23001 40267 23035
rect 40325 23001 40359 23035
rect 41512 23001 41546 23035
rect 45744 23001 45778 23035
rect 50436 23001 50470 23035
rect 52754 23001 52788 23035
rect 53748 23001 53782 23035
rect 9137 22933 9171 22967
rect 13001 22933 13035 22967
rect 15853 22933 15887 22967
rect 17417 22933 17451 22967
rect 19073 22933 19107 22967
rect 19441 22933 19475 22967
rect 22385 22933 22419 22967
rect 24409 22933 24443 22967
rect 27537 22933 27571 22967
rect 27905 22933 27939 22967
rect 29009 22933 29043 22967
rect 30021 22933 30055 22967
rect 30205 22933 30239 22967
rect 30573 22933 30607 22967
rect 31033 22933 31067 22967
rect 33333 22933 33367 22967
rect 33885 22933 33919 22967
rect 36093 22933 36127 22967
rect 37841 22933 37875 22967
rect 40969 22933 41003 22967
rect 42625 22933 42659 22967
rect 44557 22933 44591 22967
rect 55321 22933 55355 22967
rect 57621 22933 57655 22967
rect 8309 22729 8343 22763
rect 13185 22729 13219 22763
rect 14933 22729 14967 22763
rect 16037 22729 16071 22763
rect 16129 22729 16163 22763
rect 16497 22729 16531 22763
rect 17693 22729 17727 22763
rect 20177 22729 20211 22763
rect 21833 22729 21867 22763
rect 25973 22729 26007 22763
rect 27261 22729 27295 22763
rect 29193 22729 29227 22763
rect 29285 22729 29319 22763
rect 31217 22729 31251 22763
rect 32873 22729 32907 22763
rect 35725 22729 35759 22763
rect 36185 22729 36219 22763
rect 40233 22729 40267 22763
rect 42441 22729 42475 22763
rect 42901 22729 42935 22763
rect 43269 22729 43303 22763
rect 50445 22729 50479 22763
rect 50721 22729 50755 22763
rect 53113 22729 53147 22763
rect 53205 22729 53239 22763
rect 55781 22729 55815 22763
rect 57621 22729 57655 22763
rect 11713 22661 11747 22695
rect 15393 22661 15427 22695
rect 19064 22661 19098 22695
rect 26065 22661 26099 22695
rect 28058 22661 28092 22695
rect 42809 22661 42843 22695
rect 44404 22661 44438 22695
rect 45385 22661 45419 22695
rect 45845 22661 45879 22695
rect 56508 22661 56542 22695
rect 8401 22593 8435 22627
rect 13553 22593 13587 22627
rect 13645 22593 13679 22627
rect 14013 22593 14047 22627
rect 15301 22593 15335 22627
rect 17601 22593 17635 22627
rect 18061 22593 18095 22627
rect 18797 22593 18831 22627
rect 21189 22593 21223 22627
rect 21281 22593 21315 22627
rect 22957 22593 22991 22627
rect 23213 22593 23247 22627
rect 23673 22593 23707 22627
rect 23940 22593 23974 22627
rect 27813 22593 27847 22627
rect 31585 22593 31619 22627
rect 31677 22593 31711 22627
rect 32781 22593 32815 22627
rect 34345 22593 34379 22627
rect 35081 22593 35115 22627
rect 37556 22593 37590 22627
rect 38853 22593 38887 22627
rect 39120 22593 39154 22627
rect 40877 22593 40911 22627
rect 41144 22593 41178 22627
rect 44649 22593 44683 22627
rect 45937 22593 45971 22627
rect 46204 22593 46238 22627
rect 48375 22593 48409 22627
rect 49433 22593 49467 22627
rect 51365 22593 51399 22627
rect 51641 22593 51675 22627
rect 52561 22593 52595 22627
rect 53665 22593 53699 22627
rect 53932 22593 53966 22627
rect 56241 22593 56275 22627
rect 58449 22593 58483 22627
rect 5917 22525 5951 22559
rect 8217 22525 8251 22559
rect 9413 22525 9447 22559
rect 11345 22525 11379 22559
rect 11897 22525 11931 22559
rect 13737 22525 13771 22559
rect 14565 22525 14599 22559
rect 15485 22525 15519 22559
rect 15853 22525 15887 22559
rect 17785 22525 17819 22559
rect 18613 22525 18647 22559
rect 20821 22525 20855 22559
rect 21005 22525 21039 22559
rect 25789 22525 25823 22559
rect 29929 22525 29963 22559
rect 30088 22525 30122 22559
rect 30205 22525 30239 22559
rect 30941 22525 30975 22559
rect 31125 22525 31159 22559
rect 31769 22525 31803 22559
rect 33057 22525 33091 22559
rect 34069 22525 34103 22559
rect 34207 22525 34241 22559
rect 34621 22525 34655 22559
rect 35265 22525 35299 22559
rect 35817 22525 35851 22559
rect 35909 22525 35943 22559
rect 36737 22525 36771 22559
rect 37289 22525 37323 22559
rect 43085 22525 43119 22559
rect 48237 22525 48271 22559
rect 48513 22525 48547 22559
rect 49249 22525 49283 22559
rect 51503 22525 51537 22559
rect 52377 22525 52411 22559
rect 53297 22525 53331 22559
rect 55137 22525 55171 22559
rect 5273 22457 5307 22491
rect 8769 22457 8803 22491
rect 17141 22457 17175 22491
rect 21649 22457 21683 22491
rect 25513 22457 25547 22491
rect 26433 22457 26467 22491
rect 30481 22457 30515 22491
rect 35357 22457 35391 22491
rect 48789 22457 48823 22491
rect 51917 22457 51951 22491
rect 55045 22457 55079 22491
rect 5365 22389 5399 22423
rect 6653 22389 6687 22423
rect 8861 22389 8895 22423
rect 10701 22389 10735 22423
rect 12541 22389 12575 22423
rect 17233 22389 17267 22423
rect 25053 22389 25087 22423
rect 32413 22389 32447 22423
rect 33425 22389 33459 22423
rect 38669 22389 38703 22423
rect 42257 22389 42291 22423
rect 45017 22389 45051 22423
rect 47317 22389 47351 22423
rect 47593 22389 47627 22423
rect 49801 22389 49835 22423
rect 52745 22389 52779 22423
rect 57897 22389 57931 22423
rect 5641 22185 5675 22219
rect 8953 22185 8987 22219
rect 11621 22185 11655 22219
rect 13921 22185 13955 22219
rect 18061 22185 18095 22219
rect 20177 22185 20211 22219
rect 11713 22117 11747 22151
rect 31217 22117 31251 22151
rect 32137 22117 32171 22151
rect 32321 22117 32355 22151
rect 33793 22117 33827 22151
rect 35541 22117 35575 22151
rect 38025 22117 38059 22151
rect 38761 22117 38795 22151
rect 41521 22117 41555 22151
rect 43729 22117 43763 22151
rect 55597 22117 55631 22151
rect 5457 22049 5491 22083
rect 6193 22049 6227 22083
rect 9597 22049 9631 22083
rect 12265 22049 12299 22083
rect 14289 22049 14323 22083
rect 14749 22049 14783 22083
rect 16221 22049 16255 22083
rect 16865 22049 16899 22083
rect 17141 22049 17175 22083
rect 17417 22049 17451 22083
rect 22293 22049 22327 22083
rect 22937 22049 22971 22083
rect 27813 22049 27847 22083
rect 29837 22049 29871 22083
rect 31493 22049 31527 22083
rect 32873 22049 32907 22083
rect 33241 22049 33275 22083
rect 34805 22049 34839 22083
rect 34989 22049 35023 22083
rect 36093 22049 36127 22083
rect 37013 22049 37047 22083
rect 37289 22049 37323 22083
rect 39313 22049 39347 22083
rect 41429 22049 41463 22083
rect 42809 22049 42843 22083
rect 43085 22049 43119 22083
rect 46397 22049 46431 22083
rect 47041 22049 47075 22083
rect 47869 22049 47903 22083
rect 48053 22049 48087 22083
rect 51733 22049 51767 22083
rect 52653 22049 52687 22083
rect 57161 22049 57195 22083
rect 6469 21981 6503 22015
rect 8513 21981 8547 22015
rect 8769 21981 8803 22015
rect 10241 21981 10275 22015
rect 12541 21981 12575 22015
rect 12808 21981 12842 22015
rect 15577 21981 15611 22015
rect 16405 21981 16439 22015
rect 17258 21981 17292 22015
rect 20821 21981 20855 22015
rect 30104 21981 30138 22015
rect 37565 21981 37599 22015
rect 38577 21981 38611 22015
rect 42165 21981 42199 22015
rect 42625 21981 42659 22015
rect 46949 21981 46983 22015
rect 48145 21981 48179 22015
rect 50169 21981 50203 22015
rect 52377 21981 52411 22015
rect 56977 21981 57011 22015
rect 57069 21981 57103 22015
rect 57989 21981 58023 22015
rect 5181 21913 5215 21947
rect 9321 21913 9355 21947
rect 10508 21913 10542 21947
rect 22048 21913 22082 21947
rect 22385 21913 22419 21947
rect 28080 21913 28114 21947
rect 34529 21913 34563 21947
rect 47685 21913 47719 21947
rect 50436 21913 50470 21947
rect 4813 21845 4847 21879
rect 5273 21845 5307 21879
rect 6009 21845 6043 21879
rect 6101 21845 6135 21879
rect 7113 21845 7147 21879
rect 7389 21845 7423 21879
rect 9413 21845 9447 21879
rect 10057 21845 10091 21879
rect 12081 21845 12115 21879
rect 12173 21845 12207 21879
rect 16129 21845 16163 21879
rect 18429 21845 18463 21879
rect 20085 21845 20119 21879
rect 20913 21845 20947 21879
rect 24961 21845 24995 21879
rect 25329 21845 25363 21879
rect 29193 21845 29227 21879
rect 34069 21845 34103 21879
rect 35081 21845 35115 21879
rect 35449 21845 35483 21879
rect 37473 21845 37507 21879
rect 37933 21845 37967 21879
rect 42257 21845 42291 21879
rect 42717 21845 42751 21879
rect 46489 21845 46523 21879
rect 46857 21845 46891 21879
rect 48513 21845 48547 21879
rect 49985 21845 50019 21879
rect 51549 21845 51583 21879
rect 55045 21845 55079 21879
rect 56425 21845 56459 21879
rect 56609 21845 56643 21879
rect 57437 21845 57471 21879
rect 4721 21641 4755 21675
rect 6193 21641 6227 21675
rect 8953 21641 8987 21675
rect 11069 21641 11103 21675
rect 12081 21641 12115 21675
rect 14381 21641 14415 21675
rect 28825 21641 28859 21675
rect 29929 21641 29963 21675
rect 31401 21641 31435 21675
rect 32413 21641 32447 21675
rect 35265 21641 35299 21675
rect 43269 21641 43303 21675
rect 46397 21641 46431 21675
rect 48237 21641 48271 21675
rect 50997 21641 51031 21675
rect 54769 21641 54803 21675
rect 56701 21641 56735 21675
rect 57161 21641 57195 21675
rect 5080 21573 5114 21607
rect 6377 21573 6411 21607
rect 14473 21573 14507 21607
rect 28917 21573 28951 21607
rect 50537 21573 50571 21607
rect 54401 21573 54435 21607
rect 7180 21505 7214 21539
rect 7297 21505 7331 21539
rect 8217 21505 8251 21539
rect 8309 21505 8343 21539
rect 9137 21505 9171 21539
rect 10977 21505 11011 21539
rect 12725 21505 12759 21539
rect 13001 21505 13035 21539
rect 13921 21505 13955 21539
rect 29285 21505 29319 21539
rect 30389 21505 30423 21539
rect 42625 21505 42659 21539
rect 46949 21505 46983 21539
rect 47593 21505 47627 21539
rect 48973 21505 49007 21539
rect 52377 21505 52411 21539
rect 56793 21505 56827 21539
rect 4169 21437 4203 21471
rect 4813 21437 4847 21471
rect 7021 21437 7055 21471
rect 8033 21437 8067 21471
rect 9965 21437 9999 21471
rect 11161 21437 11195 21471
rect 12863 21437 12897 21471
rect 13737 21437 13771 21471
rect 14565 21437 14599 21471
rect 16129 21437 16163 21471
rect 19073 21437 19107 21471
rect 29009 21437 29043 21471
rect 37105 21437 37139 21471
rect 49157 21437 49191 21471
rect 50261 21437 50295 21471
rect 50445 21437 50479 21471
rect 51549 21437 51583 21471
rect 56241 21437 56275 21471
rect 56517 21437 56551 21471
rect 58449 21437 58483 21471
rect 7573 21369 7607 21403
rect 10609 21369 10643 21403
rect 13277 21369 13311 21403
rect 50905 21369 50939 21403
rect 9781 21301 9815 21335
rect 10517 21301 10551 21335
rect 11989 21301 12023 21335
rect 14013 21301 14047 21335
rect 15577 21301 15611 21335
rect 19625 21301 19659 21335
rect 25329 21301 25363 21335
rect 28365 21301 28399 21335
rect 28457 21301 28491 21335
rect 31033 21301 31067 21335
rect 35633 21301 35667 21335
rect 37565 21301 37599 21335
rect 42165 21301 42199 21335
rect 48421 21301 48455 21335
rect 49801 21301 49835 21335
rect 51733 21301 51767 21335
rect 57437 21301 57471 21335
rect 57897 21301 57931 21335
rect 4537 21097 4571 21131
rect 10241 21097 10275 21131
rect 12541 21097 12575 21131
rect 15761 21097 15795 21131
rect 17233 21097 17267 21131
rect 28273 21097 28307 21131
rect 34897 21097 34931 21131
rect 42165 21097 42199 21131
rect 50353 21097 50387 21131
rect 51641 21097 51675 21131
rect 57621 21097 57655 21131
rect 9137 21029 9171 21063
rect 11805 21029 11839 21063
rect 42993 21029 43027 21063
rect 45201 21029 45235 21063
rect 10425 20961 10459 20995
rect 11897 20961 11931 20995
rect 16405 20961 16439 20995
rect 28825 20961 28859 20995
rect 42441 20961 42475 20995
rect 43637 20961 43671 20995
rect 58173 20961 58207 20995
rect 5917 20893 5951 20927
rect 6377 20893 6411 20927
rect 7849 20893 7883 20927
rect 10681 20893 10715 20927
rect 13461 20893 13495 20927
rect 16129 20893 16163 20927
rect 16589 20893 16623 20927
rect 19349 20893 19383 20927
rect 22937 20893 22971 20927
rect 23673 20893 23707 20927
rect 25237 20893 25271 20927
rect 25329 20893 25363 20927
rect 26065 20893 26099 20927
rect 27537 20893 27571 20927
rect 29745 20893 29779 20927
rect 34161 20893 34195 20927
rect 35173 20893 35207 20927
rect 37565 20893 37599 20927
rect 37749 20893 37783 20927
rect 38945 20893 38979 20927
rect 40785 20893 40819 20927
rect 44373 20893 44407 20927
rect 52193 20893 52227 20927
rect 53941 20893 53975 20927
rect 54309 20893 54343 20927
rect 56149 20893 56183 20927
rect 56416 20893 56450 20927
rect 5650 20825 5684 20859
rect 6644 20825 6678 20859
rect 9597 20825 9631 20859
rect 15669 20825 15703 20859
rect 37013 20825 37047 20859
rect 40141 20825 40175 20859
rect 42533 20825 42567 20859
rect 43821 20825 43855 20859
rect 7757 20757 7791 20791
rect 8493 20757 8527 20791
rect 12817 20757 12851 20791
rect 13921 20757 13955 20791
rect 16221 20757 16255 20791
rect 19993 20757 20027 20791
rect 21833 20757 21867 20791
rect 22293 20757 22327 20791
rect 23029 20757 23063 20791
rect 24593 20757 24627 20791
rect 25973 20757 26007 20791
rect 26709 20757 26743 20791
rect 26985 20757 27019 20791
rect 30389 20757 30423 20791
rect 32045 20757 32079 20791
rect 33609 20757 33643 20791
rect 36645 20757 36679 20791
rect 38393 20757 38427 20791
rect 38761 20757 38795 20791
rect 39589 20757 39623 20791
rect 40233 20757 40267 20791
rect 42625 20757 42659 20791
rect 43085 20757 43119 20791
rect 44741 20757 44775 20791
rect 45569 20757 45603 20791
rect 53389 20757 53423 20791
rect 54861 20757 54895 20791
rect 56057 20757 56091 20791
rect 57529 20757 57563 20791
rect 57989 20757 58023 20791
rect 58081 20757 58115 20791
rect 5457 20553 5491 20587
rect 7757 20553 7791 20587
rect 13645 20553 13679 20587
rect 16497 20553 16531 20587
rect 17601 20553 17635 20587
rect 18521 20553 18555 20587
rect 22293 20553 22327 20587
rect 25329 20553 25363 20587
rect 25881 20553 25915 20587
rect 27261 20553 27295 20587
rect 29653 20553 29687 20587
rect 30021 20553 30055 20587
rect 30573 20553 30607 20587
rect 38853 20553 38887 20587
rect 42901 20553 42935 20587
rect 44741 20553 44775 20587
rect 48145 20553 48179 20587
rect 51181 20553 51215 20587
rect 53573 20553 53607 20587
rect 54033 20553 54067 20587
rect 54769 20553 54803 20587
rect 57069 20553 57103 20587
rect 7297 20485 7331 20519
rect 13277 20485 13311 20519
rect 19634 20485 19668 20519
rect 24216 20485 24250 20519
rect 37565 20485 37599 20519
rect 39212 20485 39246 20519
rect 44833 20485 44867 20519
rect 48237 20485 48271 20519
rect 58541 20485 58575 20519
rect 4813 20417 4847 20451
rect 8677 20417 8711 20451
rect 9680 20417 9714 20451
rect 14657 20417 14691 20451
rect 15117 20417 15151 20451
rect 15373 20417 15407 20451
rect 19901 20417 19935 20451
rect 22201 20417 22235 20451
rect 25789 20417 25823 20451
rect 27353 20417 27387 20451
rect 32505 20417 32539 20451
rect 33609 20417 33643 20451
rect 33793 20417 33827 20451
rect 34060 20417 34094 20451
rect 35265 20417 35299 20451
rect 37657 20417 37691 20451
rect 38485 20417 38519 20451
rect 42809 20417 42843 20451
rect 43913 20417 43947 20451
rect 52305 20417 52339 20451
rect 52561 20417 52595 20451
rect 53941 20417 53975 20451
rect 55413 20417 55447 20451
rect 56609 20417 56643 20451
rect 57897 20417 57931 20451
rect 2237 20349 2271 20383
rect 7113 20349 7147 20383
rect 7205 20349 7239 20383
rect 8309 20349 8343 20383
rect 9413 20349 9447 20383
rect 12817 20349 12851 20383
rect 13093 20349 13127 20383
rect 13185 20349 13219 20383
rect 13737 20349 13771 20383
rect 14381 20349 14415 20383
rect 16957 20349 16991 20383
rect 18245 20349 18279 20383
rect 19993 20349 20027 20383
rect 21005 20349 21039 20383
rect 22109 20349 22143 20383
rect 23765 20349 23799 20383
rect 23949 20349 23983 20383
rect 25973 20349 26007 20383
rect 26801 20349 26835 20383
rect 27077 20349 27111 20383
rect 27813 20349 27847 20383
rect 30113 20349 30147 20383
rect 30205 20349 30239 20383
rect 31125 20349 31159 20383
rect 31953 20349 31987 20383
rect 32597 20349 32631 20383
rect 32689 20349 32723 20383
rect 32965 20349 32999 20383
rect 35817 20349 35851 20383
rect 36553 20349 36587 20383
rect 37473 20349 37507 20383
rect 38209 20349 38243 20383
rect 38393 20349 38427 20383
rect 38945 20349 38979 20383
rect 40417 20349 40451 20383
rect 42257 20349 42291 20383
rect 42993 20349 43027 20383
rect 43269 20349 43303 20383
rect 44557 20349 44591 20383
rect 45293 20349 45327 20383
rect 46029 20349 46063 20383
rect 48329 20349 48363 20383
rect 49157 20349 49191 20383
rect 53297 20349 53331 20383
rect 54125 20349 54159 20383
rect 54585 20349 54619 20383
rect 55572 20349 55606 20383
rect 55689 20349 55723 20383
rect 55965 20349 55999 20383
rect 56425 20349 56459 20383
rect 57161 20349 57195 20383
rect 57253 20349 57287 20383
rect 7665 20281 7699 20315
rect 22661 20281 22695 20315
rect 25421 20281 25455 20315
rect 32137 20281 32171 20315
rect 35173 20281 35207 20315
rect 40325 20281 40359 20315
rect 42441 20281 42475 20315
rect 45201 20281 45235 20315
rect 48605 20281 48639 20315
rect 52745 20281 52779 20315
rect 2881 20213 2915 20247
rect 10793 20213 10827 20247
rect 11713 20213 11747 20247
rect 17693 20213 17727 20247
rect 20637 20213 20671 20247
rect 21649 20213 21683 20247
rect 23213 20213 23247 20247
rect 27721 20213 27755 20247
rect 28457 20213 28491 20247
rect 29469 20213 29503 20247
rect 31309 20213 31343 20247
rect 36001 20213 36035 20247
rect 37105 20213 37139 20247
rect 38025 20213 38059 20247
rect 41061 20213 41095 20247
rect 41429 20213 41463 20247
rect 41613 20213 41647 20247
rect 44373 20213 44407 20247
rect 45937 20213 45971 20247
rect 46673 20213 46707 20247
rect 47317 20213 47351 20247
rect 47777 20213 47811 20247
rect 56701 20213 56735 20247
rect 9597 20009 9631 20043
rect 16497 20009 16531 20043
rect 19073 20009 19107 20043
rect 20545 20009 20579 20043
rect 23857 20009 23891 20043
rect 24685 20009 24719 20043
rect 25605 20009 25639 20043
rect 27537 20009 27571 20043
rect 30941 20009 30975 20043
rect 32505 20009 32539 20043
rect 35449 20009 35483 20043
rect 37473 20009 37507 20043
rect 42809 20009 42843 20043
rect 45017 20009 45051 20043
rect 48605 20009 48639 20043
rect 48697 20009 48731 20043
rect 49801 20009 49835 20043
rect 52377 20009 52411 20043
rect 55045 20009 55079 20043
rect 57161 20009 57195 20043
rect 13921 19941 13955 19975
rect 21741 19941 21775 19975
rect 26801 19941 26835 19975
rect 33885 19941 33919 19975
rect 40693 19941 40727 19975
rect 42993 19941 43027 19975
rect 51549 19941 51583 19975
rect 57069 19941 57103 19975
rect 10241 19873 10275 19907
rect 14657 19873 14691 19907
rect 15485 19873 15519 19907
rect 17877 19873 17911 19907
rect 18521 19873 18555 19907
rect 19717 19873 19751 19907
rect 19809 19873 19843 19907
rect 21348 19873 21382 19907
rect 21465 19873 21499 19907
rect 22201 19873 22235 19907
rect 22385 19873 22419 19907
rect 25421 19873 25455 19907
rect 26387 19873 26421 19907
rect 26525 19873 26559 19907
rect 27261 19873 27295 19907
rect 33333 19873 33367 19907
rect 33492 19873 33526 19907
rect 34345 19873 34379 19907
rect 34805 19873 34839 19907
rect 35725 19873 35759 19907
rect 38393 19873 38427 19907
rect 38669 19873 38703 19907
rect 38945 19873 38979 19907
rect 39405 19873 39439 19907
rect 40325 19873 40359 19907
rect 40417 19873 40451 19907
rect 41429 19873 41463 19907
rect 43637 19873 43671 19907
rect 43796 19873 43830 19907
rect 43913 19873 43947 19907
rect 44189 19873 44223 19907
rect 46397 19873 46431 19907
rect 47225 19873 47259 19907
rect 49341 19873 49375 19907
rect 50169 19873 50203 19907
rect 51825 19873 51859 19907
rect 52837 19873 52871 19907
rect 54401 19873 54435 19907
rect 55505 19873 55539 19907
rect 57805 19873 57839 19907
rect 58173 19873 58207 19907
rect 2145 19805 2179 19839
rect 2881 19805 2915 19839
rect 3433 19805 3467 19839
rect 3801 19805 3835 19839
rect 6929 19805 6963 19839
rect 7573 19805 7607 19839
rect 9965 19805 9999 19839
rect 12541 19805 12575 19839
rect 14473 19805 14507 19839
rect 14933 19805 14967 19839
rect 17610 19805 17644 19839
rect 21189 19805 21223 19839
rect 22477 19805 22511 19839
rect 22744 19805 22778 19839
rect 26249 19805 26283 19839
rect 27445 19805 27479 19839
rect 28917 19805 28951 19839
rect 29561 19805 29595 19839
rect 29828 19805 29862 19839
rect 31125 19805 31159 19839
rect 31392 19805 31426 19839
rect 33609 19805 33643 19839
rect 34529 19805 34563 19839
rect 35081 19805 35115 19839
rect 36093 19805 36127 19839
rect 38531 19805 38565 19839
rect 39589 19805 39623 19839
rect 41245 19805 41279 19839
rect 41696 19805 41730 19839
rect 44649 19805 44683 19839
rect 44833 19805 44867 19839
rect 47041 19805 47075 19839
rect 49065 19805 49099 19839
rect 52009 19805 52043 19839
rect 55689 19805 55723 19839
rect 57529 19805 57563 19839
rect 6285 19737 6319 19771
rect 12808 19737 12842 19771
rect 14565 19737 14599 19771
rect 18613 19737 18647 19771
rect 24133 19737 24167 19771
rect 28650 19737 28684 19771
rect 36360 19737 36394 19771
rect 40233 19737 40267 19771
rect 46152 19737 46186 19771
rect 46489 19737 46523 19771
rect 47492 19737 47526 19771
rect 50414 19737 50448 19771
rect 53104 19737 53138 19771
rect 54677 19737 54711 19771
rect 55956 19737 55990 19771
rect 2789 19669 2823 19703
rect 4445 19669 4479 19703
rect 7021 19669 7055 19703
rect 7941 19669 7975 19703
rect 10057 19669 10091 19703
rect 10609 19669 10643 19703
rect 10977 19669 11011 19703
rect 14105 19669 14139 19703
rect 18153 19669 18187 19703
rect 18705 19669 18739 19703
rect 19257 19669 19291 19703
rect 19625 19669 19659 19703
rect 20361 19669 20395 19703
rect 24777 19669 24811 19703
rect 25145 19669 25179 19703
rect 25237 19669 25271 19703
rect 32689 19669 32723 19703
rect 34989 19669 35023 19703
rect 37749 19669 37783 19703
rect 39865 19669 39899 19703
rect 49157 19669 49191 19703
rect 51917 19669 51951 19703
rect 54217 19669 54251 19703
rect 54585 19669 54619 19703
rect 57621 19669 57655 19703
rect 1961 19465 1995 19499
rect 3433 19465 3467 19499
rect 3801 19465 3835 19499
rect 6745 19465 6779 19499
rect 7113 19465 7147 19499
rect 13921 19465 13955 19499
rect 16497 19465 16531 19499
rect 17325 19465 17359 19499
rect 17693 19465 17727 19499
rect 19993 19465 20027 19499
rect 20913 19465 20947 19499
rect 21373 19465 21407 19499
rect 23213 19465 23247 19499
rect 25513 19465 25547 19499
rect 26341 19465 26375 19499
rect 26801 19465 26835 19499
rect 28641 19465 28675 19499
rect 30113 19465 30147 19499
rect 30481 19465 30515 19499
rect 35449 19465 35483 19499
rect 35541 19465 35575 19499
rect 37289 19465 37323 19499
rect 37657 19465 37691 19499
rect 40141 19465 40175 19499
rect 43821 19465 43855 19499
rect 45385 19465 45419 19499
rect 48973 19465 49007 19499
rect 50169 19465 50203 19499
rect 50537 19465 50571 19499
rect 51549 19465 51583 19499
rect 54309 19465 54343 19499
rect 54401 19465 54435 19499
rect 55781 19465 55815 19499
rect 57897 19465 57931 19499
rect 3074 19397 3108 19431
rect 3893 19397 3927 19431
rect 12716 19397 12750 19431
rect 29776 19397 29810 19431
rect 40601 19397 40635 19431
rect 56508 19397 56542 19431
rect 3341 19329 3375 19363
rect 4261 19329 4295 19363
rect 6653 19329 6687 19363
rect 9781 19329 9815 19363
rect 12449 19329 12483 19363
rect 14473 19329 14507 19363
rect 15117 19329 15151 19363
rect 15384 19329 15418 19363
rect 17233 19329 17267 19363
rect 18613 19329 18647 19363
rect 18880 19329 18914 19363
rect 21281 19329 21315 19363
rect 21833 19329 21867 19363
rect 22089 19329 22123 19363
rect 24133 19329 24167 19363
rect 24400 19329 24434 19363
rect 26433 19329 26467 19363
rect 26985 19329 27019 19363
rect 27252 19329 27286 19363
rect 30021 19329 30055 19363
rect 30573 19329 30607 19363
rect 31953 19329 31987 19363
rect 32137 19329 32171 19363
rect 32393 19329 32427 19363
rect 34733 19329 34767 19363
rect 34989 19329 35023 19363
rect 35909 19329 35943 19363
rect 37749 19329 37783 19363
rect 38761 19329 38795 19363
rect 39028 19329 39062 19363
rect 40693 19329 40727 19363
rect 42708 19329 42742 19363
rect 44281 19329 44315 19363
rect 45293 19329 45327 19363
rect 45845 19329 45879 19363
rect 46112 19329 46146 19363
rect 47582 19329 47616 19363
rect 47860 19329 47894 19363
rect 50629 19329 50663 19363
rect 52929 19329 52963 19363
rect 53196 19329 53230 19363
rect 55045 19329 55079 19363
rect 56241 19329 56275 19363
rect 58449 19329 58483 19363
rect 3985 19261 4019 19295
rect 4813 19261 4847 19295
rect 6469 19261 6503 19295
rect 7849 19261 7883 19295
rect 9597 19261 9631 19295
rect 9689 19261 9723 19295
rect 10793 19261 10827 19295
rect 17049 19261 17083 19295
rect 21465 19261 21499 19295
rect 26249 19261 26283 19295
rect 30665 19261 30699 19295
rect 31401 19261 31435 19295
rect 35633 19261 35667 19295
rect 36461 19261 36495 19295
rect 37841 19261 37875 19295
rect 40785 19261 40819 19295
rect 42441 19261 42475 19295
rect 44005 19261 44039 19295
rect 44189 19261 44223 19295
rect 45109 19261 45143 19295
rect 50721 19261 50755 19295
rect 55137 19261 55171 19295
rect 8493 19193 8527 19227
rect 10149 19193 10183 19227
rect 33517 19193 33551 19227
rect 37105 19193 37139 19227
rect 40233 19193 40267 19227
rect 45753 19193 45787 19227
rect 5273 19125 5307 19159
rect 5825 19125 5859 19159
rect 7205 19125 7239 19159
rect 8217 19125 8251 19159
rect 10241 19125 10275 19159
rect 13829 19125 13863 19159
rect 18245 19125 18279 19159
rect 20361 19125 20395 19159
rect 20821 19125 20855 19159
rect 23949 19125 23983 19159
rect 25973 19125 26007 19159
rect 28365 19125 28399 19159
rect 33609 19125 33643 19159
rect 35081 19125 35115 19159
rect 38301 19125 38335 19159
rect 44649 19125 44683 19159
rect 47225 19125 47259 19159
rect 49985 19125 50019 19159
rect 57621 19125 57655 19159
rect 2145 18921 2179 18955
rect 7113 18921 7147 18955
rect 7941 18921 7975 18955
rect 10517 18921 10551 18955
rect 16037 18921 16071 18955
rect 17049 18921 17083 18955
rect 19257 18921 19291 18955
rect 24593 18921 24627 18955
rect 27077 18921 27111 18955
rect 30021 18921 30055 18955
rect 32045 18921 32079 18955
rect 34253 18921 34287 18955
rect 39129 18921 39163 18955
rect 40141 18921 40175 18955
rect 45017 18921 45051 18955
rect 46029 18921 46063 18955
rect 54125 18921 54159 18955
rect 57345 18921 57379 18955
rect 3617 18853 3651 18887
rect 10425 18853 10459 18887
rect 37657 18853 37691 18887
rect 44005 18853 44039 18887
rect 1593 18785 1627 18819
rect 3801 18785 3835 18819
rect 4445 18785 4479 18819
rect 4838 18785 4872 18819
rect 4997 18785 5031 18819
rect 5733 18785 5767 18819
rect 7389 18785 7423 18819
rect 11069 18785 11103 18819
rect 15945 18785 15979 18819
rect 16589 18785 16623 18819
rect 19809 18785 19843 18819
rect 22293 18785 22327 18819
rect 22385 18785 22419 18819
rect 25145 18785 25179 18819
rect 27997 18785 28031 18819
rect 28825 18785 28859 18819
rect 31953 18785 31987 18819
rect 32689 18785 32723 18819
rect 33425 18785 33459 18819
rect 33701 18785 33735 18819
rect 33793 18785 33827 18819
rect 35265 18785 35299 18819
rect 36277 18785 36311 18819
rect 38301 18785 38335 18819
rect 38485 18785 38519 18819
rect 44649 18785 44683 18819
rect 45569 18785 45603 18819
rect 46581 18785 46615 18819
rect 57989 18785 58023 18819
rect 1777 18717 1811 18751
rect 2237 18717 2271 18751
rect 3985 18717 4019 18751
rect 4721 18717 4755 18751
rect 6000 18717 6034 18751
rect 7573 18717 7607 18751
rect 8033 18717 8067 18751
rect 9045 18717 9079 18751
rect 9312 18717 9346 18751
rect 16405 18717 16439 18751
rect 22201 18717 22235 18751
rect 27813 18717 27847 18751
rect 28273 18717 28307 18751
rect 32505 18717 32539 18751
rect 42625 18717 42659 18751
rect 46397 18717 46431 18751
rect 51825 18717 51859 18751
rect 52469 18717 52503 18751
rect 52837 18717 52871 18751
rect 57161 18717 57195 18751
rect 1685 18649 1719 18683
rect 2504 18649 2538 18683
rect 7481 18649 7515 18683
rect 8677 18649 8711 18683
rect 25605 18649 25639 18683
rect 32413 18649 32447 18683
rect 33885 18649 33919 18683
rect 36544 18649 36578 18683
rect 37749 18649 37783 18683
rect 42892 18649 42926 18683
rect 44097 18649 44131 18683
rect 5641 18581 5675 18615
rect 16497 18581 16531 18615
rect 21649 18581 21683 18615
rect 21833 18581 21867 18615
rect 27445 18581 27479 18615
rect 27905 18581 27939 18615
rect 34713 18581 34747 18615
rect 35633 18581 35667 18615
rect 46489 18581 46523 18615
rect 51181 18581 51215 18615
rect 51917 18581 51951 18615
rect 56609 18581 56643 18615
rect 3341 18377 3375 18411
rect 3985 18377 4019 18411
rect 4077 18377 4111 18411
rect 7849 18377 7883 18411
rect 8125 18377 8159 18411
rect 8309 18377 8343 18411
rect 10609 18377 10643 18411
rect 10701 18377 10735 18411
rect 20269 18377 20303 18411
rect 27353 18377 27387 18411
rect 33793 18377 33827 18411
rect 34897 18377 34931 18411
rect 51825 18377 51859 18411
rect 52929 18377 52963 18411
rect 56609 18377 56643 18411
rect 2228 18309 2262 18343
rect 6736 18309 6770 18343
rect 50712 18309 50746 18343
rect 1961 18241 1995 18275
rect 9229 18241 9263 18275
rect 10149 18241 10183 18275
rect 27905 18241 27939 18275
rect 34345 18241 34379 18275
rect 39405 18241 39439 18275
rect 50445 18241 50479 18275
rect 56977 18241 57011 18275
rect 57897 18241 57931 18275
rect 4169 18173 4203 18207
rect 6469 18173 6503 18207
rect 8953 18173 8987 18207
rect 9112 18173 9146 18207
rect 9505 18173 9539 18207
rect 9965 18173 9999 18207
rect 10885 18173 10919 18207
rect 13001 18173 13035 18207
rect 13277 18173 13311 18207
rect 15577 18173 15611 18207
rect 15853 18173 15887 18207
rect 19165 18173 19199 18207
rect 44649 18173 44683 18207
rect 48421 18173 48455 18207
rect 48789 18173 48823 18207
rect 52561 18173 52595 18207
rect 54125 18173 54159 18207
rect 57069 18173 57103 18207
rect 57161 18173 57195 18207
rect 58449 18173 58483 18207
rect 11345 18105 11379 18139
rect 27169 18105 27203 18139
rect 45845 18105 45879 18139
rect 56517 18105 56551 18139
rect 1869 18037 1903 18071
rect 3617 18037 3651 18071
rect 4721 18037 4755 18071
rect 6009 18037 6043 18071
rect 10241 18037 10275 18071
rect 12449 18037 12483 18071
rect 13829 18037 13863 18071
rect 15025 18037 15059 18071
rect 16497 18037 16531 18071
rect 19809 18037 19843 18071
rect 25513 18037 25547 18071
rect 37565 18037 37599 18071
rect 38761 18037 38795 18071
rect 43729 18037 43763 18071
rect 44097 18037 44131 18071
rect 45017 18037 45051 18071
rect 45385 18037 45419 18071
rect 47869 18037 47903 18071
rect 49341 18037 49375 18071
rect 51917 18037 51951 18071
rect 53573 18037 53607 18071
rect 3801 17833 3835 17867
rect 10701 17833 10735 17867
rect 12541 17833 12575 17867
rect 25237 17833 25271 17867
rect 47869 17833 47903 17867
rect 51641 17833 51675 17867
rect 53665 17833 53699 17867
rect 57713 17833 57747 17867
rect 12449 17765 12483 17799
rect 14473 17765 14507 17799
rect 43821 17765 43855 17799
rect 48697 17765 48731 17799
rect 51549 17765 51583 17799
rect 4353 17697 4387 17731
rect 5549 17697 5583 17731
rect 9229 17697 9263 17731
rect 13185 17697 13219 17731
rect 15853 17697 15887 17731
rect 37933 17697 37967 17731
rect 43913 17697 43947 17731
rect 47777 17697 47811 17731
rect 48513 17697 48547 17731
rect 49249 17697 49283 17731
rect 49709 17697 49743 17731
rect 52285 17697 52319 17731
rect 53021 17697 53055 17731
rect 53573 17697 53607 17731
rect 54217 17697 54251 17731
rect 56333 17697 56367 17731
rect 7021 17629 7055 17663
rect 8769 17629 8803 17663
rect 11253 17629 11287 17663
rect 12909 17629 12943 17663
rect 16773 17629 16807 17663
rect 18245 17629 18279 17663
rect 18981 17629 19015 17663
rect 20269 17629 20303 17663
rect 21005 17629 21039 17663
rect 21649 17629 21683 17663
rect 25881 17629 25915 17663
rect 26617 17629 26651 17663
rect 30573 17629 30607 17663
rect 30849 17629 30883 17663
rect 33057 17629 33091 17663
rect 33793 17629 33827 17663
rect 36369 17629 36403 17663
rect 36645 17629 36679 17663
rect 37657 17629 37691 17663
rect 40417 17629 40451 17663
rect 41153 17629 41187 17663
rect 41337 17629 41371 17663
rect 41889 17629 41923 17663
rect 42441 17629 42475 17663
rect 45017 17629 45051 17663
rect 49065 17629 49099 17663
rect 50169 17629 50203 17663
rect 50436 17629 50470 17663
rect 54493 17629 54527 17663
rect 56600 17629 56634 17663
rect 5816 17561 5850 17595
rect 9496 17561 9530 17595
rect 15608 17561 15642 17595
rect 16221 17561 16255 17595
rect 23397 17561 23431 17595
rect 37197 17561 37231 17595
rect 42708 17561 42742 17595
rect 48237 17561 48271 17595
rect 54033 17561 54067 17595
rect 55137 17561 55171 17595
rect 6929 17493 6963 17527
rect 10609 17493 10643 17527
rect 13001 17493 13035 17527
rect 17693 17493 17727 17527
rect 18429 17493 18463 17527
rect 19625 17493 19659 17527
rect 20361 17493 20395 17527
rect 21097 17493 21131 17527
rect 25329 17493 25363 17527
rect 26065 17493 26099 17527
rect 30021 17493 30055 17527
rect 31401 17493 31435 17527
rect 33701 17493 33735 17527
rect 34437 17493 34471 17527
rect 35817 17493 35851 17527
rect 37289 17493 37323 17527
rect 37749 17493 37783 17527
rect 39681 17493 39715 17527
rect 39865 17493 39899 17527
rect 40601 17493 40635 17527
rect 44557 17493 44591 17527
rect 45661 17493 45695 17527
rect 48329 17493 48363 17527
rect 49157 17493 49191 17527
rect 52009 17493 52043 17527
rect 52101 17493 52135 17527
rect 52469 17493 52503 17527
rect 54125 17493 54159 17527
rect 4997 17289 5031 17323
rect 7113 17289 7147 17323
rect 8677 17289 8711 17323
rect 14473 17289 14507 17323
rect 16681 17289 16715 17323
rect 18061 17289 18095 17323
rect 18521 17289 18555 17323
rect 20361 17289 20395 17323
rect 20821 17289 20855 17323
rect 21189 17289 21223 17323
rect 23949 17289 23983 17323
rect 25421 17289 25455 17323
rect 27353 17289 27387 17323
rect 30941 17289 30975 17323
rect 33517 17289 33551 17323
rect 34345 17289 34379 17323
rect 35909 17289 35943 17323
rect 36921 17289 36955 17323
rect 39681 17289 39715 17323
rect 40141 17289 40175 17323
rect 40969 17289 41003 17323
rect 42257 17289 42291 17323
rect 44373 17289 44407 17323
rect 44833 17289 44867 17323
rect 45937 17289 45971 17323
rect 48973 17289 49007 17323
rect 51825 17289 51859 17323
rect 52193 17289 52227 17323
rect 54493 17289 54527 17323
rect 8217 17221 8251 17255
rect 9413 17221 9447 17255
rect 9873 17221 9907 17255
rect 14924 17221 14958 17255
rect 33057 17221 33091 17255
rect 42441 17221 42475 17255
rect 47860 17221 47894 17255
rect 49341 17221 49375 17255
rect 54953 17221 54987 17255
rect 7573 17153 7607 17187
rect 10885 17153 10919 17187
rect 11989 17153 12023 17187
rect 12256 17153 12290 17187
rect 13829 17153 13863 17187
rect 13921 17153 13955 17187
rect 14657 17153 14691 17187
rect 17049 17153 17083 17187
rect 18429 17153 18463 17187
rect 18981 17153 19015 17187
rect 19248 17153 19282 17187
rect 21833 17153 21867 17187
rect 22089 17153 22123 17187
rect 24041 17153 24075 17187
rect 25053 17153 25087 17187
rect 25789 17153 25823 17187
rect 25881 17153 25915 17187
rect 29561 17153 29595 17187
rect 29817 17153 29851 17187
rect 33149 17153 33183 17187
rect 36277 17153 36311 17187
rect 37289 17153 37323 17187
rect 37545 17153 37579 17187
rect 39773 17153 39807 17187
rect 40601 17153 40635 17187
rect 44741 17153 44775 17187
rect 45477 17153 45511 17187
rect 45569 17153 45603 17187
rect 46765 17153 46799 17187
rect 47593 17153 47627 17187
rect 50169 17153 50203 17187
rect 50445 17153 50479 17187
rect 51181 17153 51215 17187
rect 51365 17153 51399 17187
rect 53113 17153 53147 17187
rect 53380 17153 53414 17187
rect 56011 17153 56045 17187
rect 56885 17153 56919 17187
rect 3985 17085 4019 17119
rect 7205 17085 7239 17119
rect 7389 17085 7423 17119
rect 8861 17085 8895 17119
rect 9965 17085 9999 17119
rect 10149 17085 10183 17119
rect 14105 17085 14139 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 18613 17085 18647 17119
rect 20545 17085 20579 17119
rect 20729 17085 20763 17119
rect 24133 17085 24167 17119
rect 24409 17085 24443 17119
rect 26065 17085 26099 17119
rect 27445 17085 27479 17119
rect 27537 17085 27571 17119
rect 28825 17085 28859 17119
rect 31585 17085 31619 17119
rect 32965 17085 32999 17119
rect 34161 17085 34195 17119
rect 34253 17085 34287 17119
rect 36369 17085 36403 17119
rect 36461 17085 36495 17119
rect 39497 17085 39531 17119
rect 40325 17085 40359 17119
rect 40509 17085 40543 17119
rect 41613 17085 41647 17119
rect 44925 17085 44959 17119
rect 45385 17085 45419 17119
rect 46673 17085 46707 17119
rect 47317 17085 47351 17119
rect 50307 17085 50341 17119
rect 50721 17085 50755 17119
rect 51641 17085 51675 17119
rect 51733 17085 51767 17119
rect 55873 17085 55907 17119
rect 56149 17085 56183 17119
rect 56425 17085 56459 17119
rect 57069 17085 57103 17119
rect 4721 17017 4755 17051
rect 9505 17017 9539 17051
rect 13369 17017 13403 17051
rect 23213 17017 23247 17051
rect 26801 17017 26835 17051
rect 3433 16949 3467 16983
rect 6745 16949 6779 16983
rect 10333 16949 10367 16983
rect 13461 16949 13495 16983
rect 16037 16949 16071 16983
rect 16497 16949 16531 16983
rect 17969 16949 18003 16983
rect 21557 16949 21591 16983
rect 23581 16949 23615 16983
rect 26985 16949 27019 16983
rect 29469 16949 29503 16983
rect 31033 16949 31067 16983
rect 33885 16949 33919 16983
rect 34713 16949 34747 16983
rect 35725 16949 35759 16983
rect 38669 16949 38703 16983
rect 39221 16949 39255 16983
rect 41061 16949 41095 16983
rect 43729 16949 43763 16983
rect 46029 16949 46063 16983
rect 49525 16949 49559 16983
rect 52561 16949 52595 16983
rect 55229 16949 55263 16983
rect 6285 16745 6319 16779
rect 7573 16745 7607 16779
rect 10425 16745 10459 16779
rect 18797 16745 18831 16779
rect 19257 16745 19291 16779
rect 22477 16745 22511 16779
rect 26249 16745 26283 16779
rect 29929 16745 29963 16779
rect 32781 16745 32815 16779
rect 34529 16745 34563 16779
rect 36829 16745 36863 16779
rect 37841 16745 37875 16779
rect 51365 16745 51399 16779
rect 55137 16745 55171 16779
rect 3801 16677 3835 16711
rect 39037 16677 39071 16711
rect 44833 16677 44867 16711
rect 49801 16677 49835 16711
rect 3617 16609 3651 16643
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 6837 16609 6871 16643
rect 9781 16609 9815 16643
rect 9965 16609 9999 16643
rect 10701 16609 10735 16643
rect 11069 16609 11103 16643
rect 11897 16609 11931 16643
rect 13921 16609 13955 16643
rect 14749 16609 14783 16643
rect 14908 16609 14942 16643
rect 15301 16609 15335 16643
rect 15945 16609 15979 16643
rect 16589 16609 16623 16643
rect 17417 16609 17451 16643
rect 20039 16609 20073 16643
rect 20177 16609 20211 16643
rect 20453 16609 20487 16643
rect 20913 16609 20947 16643
rect 21097 16609 21131 16643
rect 24869 16609 24903 16643
rect 26617 16609 26651 16643
rect 28457 16609 28491 16643
rect 29193 16609 29227 16643
rect 30113 16609 30147 16643
rect 30297 16609 30331 16643
rect 30849 16609 30883 16643
rect 31033 16609 31067 16643
rect 31493 16609 31527 16643
rect 31769 16609 31803 16643
rect 31886 16609 31920 16643
rect 32689 16609 32723 16643
rect 34161 16609 34195 16643
rect 37013 16609 37047 16643
rect 37197 16609 37231 16643
rect 39497 16609 39531 16643
rect 39681 16609 39715 16643
rect 41245 16609 41279 16643
rect 41705 16609 41739 16643
rect 43453 16609 43487 16643
rect 45017 16609 45051 16643
rect 47317 16609 47351 16643
rect 49341 16609 49375 16643
rect 51457 16609 51491 16643
rect 53389 16609 53423 16643
rect 56149 16609 56183 16643
rect 58173 16609 58207 16643
rect 4629 16541 4663 16575
rect 9689 16541 9723 16575
rect 15025 16541 15059 16575
rect 15761 16541 15795 16575
rect 17684 16541 17718 16575
rect 19901 16541 19935 16575
rect 23949 16541 23983 16575
rect 26884 16541 26918 16575
rect 29009 16541 29043 16575
rect 30389 16541 30423 16575
rect 32045 16541 32079 16575
rect 33905 16541 33939 16575
rect 35449 16541 35483 16575
rect 37289 16541 37323 16575
rect 38485 16541 38519 16575
rect 38623 16541 38657 16575
rect 38761 16541 38795 16575
rect 40989 16541 41023 16575
rect 43720 16541 43754 16575
rect 45284 16541 45318 16575
rect 55873 16541 55907 16575
rect 4169 16473 4203 16507
rect 5273 16473 5307 16507
rect 12164 16473 12198 16507
rect 16037 16473 16071 16507
rect 21189 16473 21223 16507
rect 25136 16473 25170 16507
rect 29101 16473 29135 16507
rect 35716 16473 35750 16507
rect 41950 16473 41984 16507
rect 47584 16473 47618 16507
rect 48789 16473 48823 16507
rect 53656 16473 53690 16507
rect 55321 16473 55355 16507
rect 56416 16473 56450 16507
rect 57621 16473 57655 16507
rect 2973 16405 3007 16439
rect 9321 16405 9355 16439
rect 11713 16405 11747 16439
rect 13277 16405 13311 16439
rect 14105 16405 14139 16439
rect 23397 16405 23431 16439
rect 24685 16405 24719 16439
rect 27997 16405 28031 16439
rect 28641 16405 28675 16439
rect 30757 16405 30791 16439
rect 37657 16405 37691 16439
rect 39865 16405 39899 16439
rect 43085 16405 43119 16439
rect 46397 16405 46431 16439
rect 48697 16405 48731 16439
rect 52101 16405 52135 16439
rect 54769 16405 54803 16439
rect 57529 16405 57563 16439
rect 3709 16201 3743 16235
rect 4077 16201 4111 16235
rect 12817 16201 12851 16235
rect 14289 16201 14323 16235
rect 15117 16201 15151 16235
rect 15485 16201 15519 16235
rect 19073 16201 19107 16235
rect 19533 16201 19567 16235
rect 21281 16201 21315 16235
rect 21833 16201 21867 16235
rect 22201 16201 22235 16235
rect 24225 16201 24259 16235
rect 27261 16201 27295 16235
rect 28549 16201 28583 16235
rect 31401 16201 31435 16235
rect 32781 16201 32815 16235
rect 38669 16201 38703 16235
rect 40509 16201 40543 16235
rect 41613 16201 41647 16235
rect 49617 16201 49651 16235
rect 52285 16201 52319 16235
rect 54309 16201 54343 16235
rect 55413 16201 55447 16235
rect 57161 16201 57195 16235
rect 2320 16133 2354 16167
rect 7512 16133 7546 16167
rect 7849 16133 7883 16167
rect 9220 16133 9254 16167
rect 15577 16133 15611 16167
rect 19441 16133 19475 16167
rect 20168 16133 20202 16167
rect 23112 16133 23146 16167
rect 27353 16133 27387 16167
rect 27813 16133 27847 16167
rect 34560 16133 34594 16167
rect 39396 16133 39430 16167
rect 4169 16065 4203 16099
rect 4537 16065 4571 16099
rect 7757 16065 7791 16099
rect 8953 16065 8987 16099
rect 13461 16065 13495 16099
rect 13645 16065 13679 16099
rect 17049 16065 17083 16099
rect 17316 16065 17350 16099
rect 19901 16065 19935 16099
rect 21649 16065 21683 16099
rect 25421 16065 25455 16099
rect 26157 16065 26191 16099
rect 26341 16065 26375 16099
rect 26709 16065 26743 16099
rect 29662 16065 29696 16099
rect 29929 16065 29963 16099
rect 30021 16065 30055 16099
rect 30288 16065 30322 16099
rect 34805 16065 34839 16099
rect 35725 16065 35759 16099
rect 35992 16065 36026 16099
rect 37289 16065 37323 16099
rect 37841 16065 37875 16099
rect 39129 16065 39163 16099
rect 42809 16065 42843 16099
rect 44327 16065 44361 16099
rect 45385 16065 45419 16099
rect 48145 16065 48179 16099
rect 48973 16065 49007 16099
rect 49709 16065 49743 16099
rect 52009 16065 52043 16099
rect 54861 16065 54895 16099
rect 56793 16065 56827 16099
rect 58449 16065 58483 16099
rect 2053 15997 2087 16031
rect 4353 15997 4387 16031
rect 5089 15997 5123 16031
rect 6193 15997 6227 16031
rect 8401 15997 8435 16031
rect 14933 15997 14967 16031
rect 15669 15997 15703 16031
rect 19625 15997 19659 16031
rect 22293 15997 22327 16031
rect 22477 15997 22511 16031
rect 22845 15997 22879 16031
rect 25145 15997 25179 16031
rect 25283 15997 25317 16031
rect 27077 15997 27111 16031
rect 28365 15997 28399 16031
rect 38025 15997 38059 16031
rect 42257 15997 42291 16031
rect 42901 15997 42935 16031
rect 43085 15997 43119 16031
rect 44189 15997 44223 16031
rect 44465 15997 44499 16031
rect 45201 15997 45235 16031
rect 50997 15997 51031 16031
rect 54033 15997 54067 16031
rect 54217 15997 54251 16031
rect 56517 15997 56551 16031
rect 56701 15997 56735 16031
rect 57897 15997 57931 16031
rect 3433 15929 3467 15963
rect 6377 15929 6411 15963
rect 25697 15929 25731 15963
rect 37105 15929 37139 15963
rect 42441 15929 42475 15963
rect 44741 15929 44775 15963
rect 53757 15929 53791 15963
rect 54677 15929 54711 15963
rect 5549 15861 5583 15895
rect 10333 15861 10367 15895
rect 14657 15861 14691 15895
rect 18429 15861 18463 15895
rect 18981 15861 19015 15895
rect 24501 15861 24535 15895
rect 27721 15861 27755 15895
rect 33149 15861 33183 15895
rect 33425 15861 33459 15895
rect 43545 15861 43579 15895
rect 47593 15861 47627 15895
rect 50353 15861 50387 15895
rect 50445 15861 50479 15895
rect 51365 15861 51399 15895
rect 56241 15861 56275 15895
rect 6929 15657 6963 15691
rect 8493 15657 8527 15691
rect 4537 15589 4571 15623
rect 10149 15589 10183 15623
rect 24133 15589 24167 15623
rect 27445 15589 27479 15623
rect 30113 15589 30147 15623
rect 30941 15589 30975 15623
rect 31953 15589 31987 15623
rect 42349 15589 42383 15623
rect 43177 15589 43211 15623
rect 43269 15589 43303 15623
rect 44281 15589 44315 15623
rect 48605 15589 48639 15623
rect 52377 15589 52411 15623
rect 57253 15589 57287 15623
rect 3893 15521 3927 15555
rect 4077 15521 4111 15555
rect 4930 15521 4964 15555
rect 5089 15521 5123 15555
rect 6377 15521 6411 15555
rect 7665 15521 7699 15555
rect 16773 15521 16807 15555
rect 18429 15521 18463 15555
rect 22753 15521 22787 15555
rect 24409 15521 24443 15555
rect 26065 15521 26099 15555
rect 28089 15521 28123 15555
rect 28733 15521 28767 15555
rect 30665 15521 30699 15555
rect 31493 15521 31527 15555
rect 41981 15521 42015 15555
rect 42625 15521 42659 15555
rect 43821 15521 43855 15555
rect 44557 15521 44591 15555
rect 47777 15521 47811 15555
rect 48053 15521 48087 15555
rect 49249 15521 49283 15555
rect 50997 15521 51031 15555
rect 51733 15521 51767 15555
rect 53021 15521 53055 15555
rect 56333 15521 56367 15555
rect 56609 15521 56643 15555
rect 57897 15521 57931 15555
rect 2053 15453 2087 15487
rect 4813 15453 4847 15487
rect 6469 15453 6503 15487
rect 6561 15453 6595 15487
rect 7389 15453 7423 15487
rect 9689 15453 9723 15487
rect 12541 15453 12575 15487
rect 12909 15453 12943 15487
rect 15761 15453 15795 15487
rect 18153 15453 18187 15487
rect 30481 15453 30515 15487
rect 37565 15453 37599 15487
rect 42809 15453 42843 15487
rect 48237 15453 48271 15487
rect 51089 15453 51123 15487
rect 52009 15453 52043 15487
rect 54125 15453 54159 15487
rect 54861 15453 54895 15487
rect 55321 15453 55355 15487
rect 2298 15385 2332 15419
rect 5733 15385 5767 15419
rect 18245 15385 18279 15419
rect 23020 15385 23054 15419
rect 26332 15385 26366 15419
rect 27537 15385 27571 15419
rect 30573 15385 30607 15419
rect 48145 15385 48179 15419
rect 49709 15385 49743 15419
rect 3433 15317 3467 15351
rect 6101 15317 6135 15351
rect 7021 15317 7055 15351
rect 7481 15317 7515 15351
rect 8125 15317 8159 15351
rect 9137 15317 9171 15351
rect 11989 15317 12023 15351
rect 13461 15317 13495 15351
rect 15117 15317 15151 15351
rect 17417 15317 17451 15351
rect 17785 15317 17819 15351
rect 18981 15317 19015 15351
rect 19533 15317 19567 15351
rect 25053 15317 25087 15351
rect 29377 15317 29411 15351
rect 37933 15317 37967 15351
rect 42717 15317 42751 15351
rect 48697 15317 48731 15351
rect 50629 15317 50663 15351
rect 51181 15317 51215 15351
rect 51549 15317 51583 15351
rect 51917 15317 51951 15351
rect 52469 15317 52503 15351
rect 53573 15317 53607 15351
rect 54309 15317 54343 15351
rect 55965 15317 55999 15351
rect 56793 15317 56827 15351
rect 56885 15317 56919 15351
rect 57345 15317 57379 15351
rect 2145 15113 2179 15147
rect 4261 15113 4295 15147
rect 5365 15113 5399 15147
rect 6745 15113 6779 15147
rect 7941 15113 7975 15147
rect 9229 15113 9263 15147
rect 12173 15113 12207 15147
rect 14105 15113 14139 15147
rect 17601 15113 17635 15147
rect 18981 15113 19015 15147
rect 23765 15113 23799 15147
rect 29377 15113 29411 15147
rect 30113 15113 30147 15147
rect 43637 15113 43671 15147
rect 49709 15113 49743 15147
rect 50629 15113 50663 15147
rect 50721 15113 50755 15147
rect 53665 15113 53699 15147
rect 54493 15113 54527 15147
rect 3148 15045 3182 15079
rect 12081 15045 12115 15079
rect 12633 15045 12667 15079
rect 17509 15045 17543 15079
rect 23857 15045 23891 15079
rect 24501 15045 24535 15079
rect 36001 15045 36035 15079
rect 47860 15045 47894 15079
rect 51856 15045 51890 15079
rect 54953 15045 54987 15079
rect 56600 15045 56634 15079
rect 2881 14977 2915 15011
rect 4353 14977 4387 15011
rect 6193 14977 6227 15011
rect 7849 14977 7883 15011
rect 12541 14977 12575 15011
rect 14841 14977 14875 15011
rect 15209 14977 15243 15011
rect 15301 14977 15335 15011
rect 18153 14977 18187 15011
rect 18429 14977 18463 15011
rect 23213 14977 23247 15011
rect 28733 14977 28767 15011
rect 30205 14977 30239 15011
rect 43085 14977 43119 15011
rect 47593 14977 47627 15011
rect 50261 14977 50295 15011
rect 52101 14977 52135 15011
rect 54033 14977 54067 15011
rect 54125 14977 54159 15011
rect 54861 14977 54895 15011
rect 56333 14977 56367 15011
rect 57897 14977 57931 15011
rect 2789 14909 2823 14943
rect 7389 14909 7423 14943
rect 8493 14909 8527 14943
rect 9045 14909 9079 14943
rect 9137 14909 9171 14943
rect 9873 14909 9907 14943
rect 12817 14909 12851 14943
rect 13185 14909 13219 14943
rect 15117 14909 15151 14943
rect 15761 14909 15795 14943
rect 23949 14909 23983 14943
rect 37289 14909 37323 14943
rect 43729 14909 43763 14943
rect 49065 14909 49099 14943
rect 50077 14909 50111 14943
rect 50169 14909 50203 14943
rect 54217 14909 54251 14943
rect 55045 14909 55079 14943
rect 55321 14909 55355 14943
rect 9597 14841 9631 14875
rect 10793 14841 10827 14875
rect 15669 14841 15703 14875
rect 36277 14841 36311 14875
rect 48973 14841 49007 14875
rect 55965 14841 55999 14875
rect 4997 14773 5031 14807
rect 5549 14773 5583 14807
rect 10517 14773 10551 14807
rect 11253 14773 11287 14807
rect 13829 14773 13863 14807
rect 16405 14773 16439 14807
rect 23397 14773 23431 14807
rect 31493 14773 31527 14807
rect 32413 14773 32447 14807
rect 33057 14773 33091 14807
rect 33609 14773 33643 14807
rect 36829 14773 36863 14807
rect 37933 14773 37967 14807
rect 41797 14773 41831 14807
rect 44373 14773 44407 14807
rect 45017 14773 45051 14807
rect 45385 14773 45419 14807
rect 53573 14773 53607 14807
rect 57713 14773 57747 14807
rect 58541 14773 58575 14807
rect 3801 14569 3835 14603
rect 6837 14569 6871 14603
rect 8953 14569 8987 14603
rect 12909 14569 12943 14603
rect 14105 14569 14139 14603
rect 23213 14569 23247 14603
rect 24225 14569 24259 14603
rect 35265 14569 35299 14603
rect 38761 14569 38795 14603
rect 39129 14569 39163 14603
rect 44741 14569 44775 14603
rect 50169 14569 50203 14603
rect 54493 14569 54527 14603
rect 8125 14501 8159 14535
rect 17969 14501 18003 14535
rect 22937 14501 22971 14535
rect 29561 14501 29595 14535
rect 32965 14501 32999 14535
rect 37657 14501 37691 14535
rect 40049 14501 40083 14535
rect 41889 14501 41923 14535
rect 51365 14501 51399 14535
rect 4353 14433 4387 14467
rect 4813 14433 4847 14467
rect 7573 14433 7607 14467
rect 8585 14433 8619 14467
rect 11069 14433 11103 14467
rect 13553 14433 13587 14467
rect 15025 14433 15059 14467
rect 15301 14433 15335 14467
rect 15761 14433 15795 14467
rect 16405 14433 16439 14467
rect 19809 14433 19843 14467
rect 20085 14433 20119 14467
rect 23765 14433 23799 14467
rect 24961 14433 24995 14467
rect 26157 14433 26191 14467
rect 29377 14433 29411 14467
rect 30113 14433 30147 14467
rect 31953 14433 31987 14467
rect 32321 14433 32355 14467
rect 33057 14433 33091 14467
rect 34345 14433 34379 14467
rect 35909 14433 35943 14467
rect 37105 14433 37139 14467
rect 38301 14433 38335 14467
rect 41797 14433 41831 14467
rect 42441 14433 42475 14467
rect 43269 14433 43303 14467
rect 44189 14433 44223 14467
rect 45109 14433 45143 14467
rect 45293 14433 45327 14467
rect 49341 14433 49375 14467
rect 49525 14433 49559 14467
rect 50951 14433 50985 14467
rect 51089 14433 51123 14467
rect 51825 14433 51859 14467
rect 55965 14433 55999 14467
rect 56103 14433 56137 14467
rect 56241 14433 56275 14467
rect 56517 14433 56551 14467
rect 57161 14433 57195 14467
rect 57713 14433 57747 14467
rect 57805 14433 57839 14467
rect 58265 14433 58299 14467
rect 4169 14365 4203 14399
rect 5457 14365 5491 14399
rect 7732 14365 7766 14399
rect 7849 14365 7883 14399
rect 8769 14365 8803 14399
rect 10077 14365 10111 14399
rect 10333 14365 10367 14399
rect 11529 14365 11563 14399
rect 13461 14365 13495 14399
rect 14749 14365 14783 14399
rect 14887 14365 14921 14399
rect 15945 14365 15979 14399
rect 16957 14365 16991 14399
rect 18521 14365 18555 14399
rect 20269 14365 20303 14399
rect 20821 14365 20855 14399
rect 25973 14365 26007 14399
rect 26985 14365 27019 14399
rect 31217 14365 31251 14399
rect 32597 14365 32631 14399
rect 35817 14365 35851 14399
rect 36737 14365 36771 14399
rect 37289 14365 37323 14399
rect 40233 14365 40267 14399
rect 42257 14365 42291 14399
rect 43545 14365 43579 14399
rect 47409 14365 47443 14399
rect 49249 14365 49283 14399
rect 50813 14365 50847 14399
rect 52009 14365 52043 14399
rect 53113 14365 53147 14399
rect 53380 14365 53414 14399
rect 56977 14365 57011 14399
rect 4261 14297 4295 14331
rect 5702 14297 5736 14331
rect 10793 14297 10827 14331
rect 11796 14297 11830 14331
rect 13369 14297 13403 14331
rect 19073 14297 19107 14331
rect 25421 14297 25455 14331
rect 29929 14297 29963 14331
rect 31401 14297 31435 14331
rect 35725 14297 35759 14331
rect 42349 14297 42383 14331
rect 43177 14297 43211 14331
rect 47676 14297 47710 14331
rect 57621 14297 57655 14331
rect 6929 14229 6963 14263
rect 10425 14229 10459 14263
rect 10885 14229 10919 14263
rect 13001 14229 13035 14263
rect 20177 14229 20211 14263
rect 20637 14229 20671 14263
rect 21373 14229 21407 14263
rect 24409 14229 24443 14263
rect 25605 14229 25639 14263
rect 26065 14229 26099 14263
rect 26433 14229 26467 14263
rect 28733 14229 28767 14263
rect 30021 14229 30055 14263
rect 30665 14229 30699 14263
rect 32505 14229 32539 14263
rect 33701 14229 33735 14263
rect 33793 14229 33827 14263
rect 35357 14229 35391 14263
rect 36185 14229 36219 14263
rect 37197 14229 37231 14263
rect 37749 14229 37783 14263
rect 40877 14229 40911 14263
rect 41153 14229 41187 14263
rect 42717 14229 42751 14263
rect 43085 14229 43119 14263
rect 45385 14229 45419 14263
rect 45753 14229 45787 14263
rect 47317 14229 47351 14263
rect 48789 14229 48823 14263
rect 48881 14229 48915 14263
rect 49985 14229 50019 14263
rect 53021 14229 53055 14263
rect 54861 14229 54895 14263
rect 55321 14229 55355 14263
rect 57253 14229 57287 14263
rect 7297 14025 7331 14059
rect 8033 14025 8067 14059
rect 12909 14025 12943 14059
rect 14933 14025 14967 14059
rect 16497 14025 16531 14059
rect 18061 14025 18095 14059
rect 18429 14025 18463 14059
rect 20821 14025 20855 14059
rect 23121 14025 23155 14059
rect 23489 14025 23523 14059
rect 24593 14025 24627 14059
rect 26249 14025 26283 14059
rect 26617 14025 26651 14059
rect 29837 14025 29871 14059
rect 31953 14025 31987 14059
rect 36001 14025 36035 14059
rect 36093 14025 36127 14059
rect 39497 14025 39531 14059
rect 39957 14025 39991 14059
rect 40417 14025 40451 14059
rect 42257 14025 42291 14059
rect 46673 14025 46707 14059
rect 48329 14025 48363 14059
rect 49341 14025 49375 14059
rect 50813 14025 50847 14059
rect 51549 14025 51583 14059
rect 54493 14025 54527 14059
rect 56057 14025 56091 14059
rect 57529 14025 57563 14059
rect 7389 13957 7423 13991
rect 8309 13957 8343 13991
rect 9628 13957 9662 13991
rect 10057 13957 10091 13991
rect 11345 13957 11379 13991
rect 11796 13957 11830 13991
rect 18521 13957 18555 13991
rect 28724 13957 28758 13991
rect 33272 13957 33306 13991
rect 34888 13957 34922 13991
rect 36553 13957 36587 13991
rect 41133 13957 41167 13991
rect 44741 13957 44775 13991
rect 56394 13957 56428 13991
rect 57897 13957 57931 13991
rect 11529 13889 11563 13923
rect 13553 13889 13587 13923
rect 13820 13889 13854 13923
rect 15117 13889 15151 13923
rect 15373 13889 15407 13923
rect 17969 13889 18003 13923
rect 19441 13889 19475 13923
rect 19708 13889 19742 13923
rect 23029 13889 23063 13923
rect 25697 13889 25731 13923
rect 27169 13889 27203 13923
rect 30113 13889 30147 13923
rect 30297 13889 30331 13923
rect 31033 13889 31067 13923
rect 33517 13889 33551 13923
rect 34621 13889 34655 13923
rect 36461 13889 36495 13923
rect 37289 13889 37323 13923
rect 38209 13889 38243 13923
rect 38485 13889 38519 13923
rect 39129 13889 39163 13923
rect 39589 13889 39623 13923
rect 43821 13889 43855 13923
rect 43938 13889 43972 13923
rect 44097 13889 44131 13923
rect 45293 13889 45327 13923
rect 45560 13889 45594 13923
rect 47409 13889 47443 13923
rect 48881 13889 48915 13923
rect 49433 13889 49467 13923
rect 49700 13889 49734 13923
rect 50905 13889 50939 13923
rect 52193 13889 52227 13923
rect 53380 13889 53414 13923
rect 54953 13889 54987 13923
rect 58449 13889 58483 13923
rect 7573 13821 7607 13855
rect 9873 13821 9907 13855
rect 10609 13821 10643 13855
rect 13369 13821 13403 13855
rect 18705 13821 18739 13855
rect 21465 13821 21499 13855
rect 23581 13821 23615 13855
rect 23673 13821 23707 13855
rect 23949 13821 23983 13855
rect 25145 13821 25179 13855
rect 25973 13821 26007 13855
rect 26157 13821 26191 13855
rect 28457 13821 28491 13855
rect 31150 13821 31184 13855
rect 31309 13821 31343 13855
rect 34161 13821 34195 13855
rect 36645 13821 36679 13855
rect 37473 13821 37507 13855
rect 38347 13821 38381 13855
rect 39405 13821 39439 13855
rect 40509 13821 40543 13855
rect 40693 13821 40727 13855
rect 40877 13821 40911 13855
rect 42717 13821 42751 13855
rect 42901 13821 42935 13855
rect 43085 13821 43119 13855
rect 51641 13821 51675 13855
rect 53113 13821 53147 13855
rect 55505 13821 55539 13855
rect 56149 13821 56183 13855
rect 24961 13753 24995 13787
rect 30757 13753 30791 13787
rect 32137 13753 32171 13787
rect 37933 13753 37967 13787
rect 43545 13753 43579 13787
rect 6837 13685 6871 13719
rect 6929 13685 6963 13719
rect 8493 13685 8527 13719
rect 17325 13685 17359 13719
rect 19073 13685 19107 13719
rect 20913 13685 20947 13719
rect 22385 13685 22419 13719
rect 27813 13685 27847 13719
rect 28089 13685 28123 13719
rect 33609 13685 33643 13719
rect 40049 13685 40083 13719
rect 45017 13685 45051 13719
rect 46765 13685 46799 13719
rect 53021 13685 53055 13719
rect 10057 13481 10091 13515
rect 12449 13481 12483 13515
rect 18705 13481 18739 13515
rect 19257 13481 19291 13515
rect 21189 13481 21223 13515
rect 23857 13481 23891 13515
rect 26433 13481 26467 13515
rect 45845 13481 45879 13515
rect 46673 13481 46707 13515
rect 49709 13481 49743 13515
rect 55597 13481 55631 13515
rect 56057 13481 56091 13515
rect 7389 13413 7423 13447
rect 15669 13413 15703 13447
rect 31033 13413 31067 13447
rect 32505 13413 32539 13447
rect 33977 13413 34011 13447
rect 43085 13413 43119 13447
rect 56241 13413 56275 13447
rect 7481 13345 7515 13379
rect 9413 13345 9447 13379
rect 10701 13345 10735 13379
rect 13001 13345 13035 13379
rect 13921 13345 13955 13379
rect 14749 13345 14783 13379
rect 16221 13345 16255 13379
rect 16405 13345 16439 13379
rect 17325 13345 17359 13379
rect 20453 13345 20487 13379
rect 21833 13345 21867 13379
rect 24225 13345 24259 13379
rect 25145 13345 25179 13379
rect 25421 13345 25455 13379
rect 25697 13345 25731 13379
rect 26157 13345 26191 13379
rect 31953 13345 31987 13379
rect 34713 13345 34747 13379
rect 41705 13345 41739 13379
rect 45201 13345 45235 13379
rect 46397 13345 46431 13379
rect 49065 13345 49099 13379
rect 56793 13345 56827 13379
rect 57253 13345 57287 13379
rect 58449 13345 58483 13379
rect 3525 13277 3559 13311
rect 4261 13277 4295 13311
rect 6009 13277 6043 13311
rect 14565 13277 14599 13311
rect 16129 13277 16163 13311
rect 17581 13277 17615 13311
rect 19901 13277 19935 13311
rect 20060 13277 20094 13311
rect 20177 13277 20211 13311
rect 20913 13277 20947 13311
rect 21097 13277 21131 13311
rect 21649 13277 21683 13311
rect 22477 13277 22511 13311
rect 22733 13277 22767 13311
rect 25304 13277 25338 13311
rect 26341 13277 26375 13311
rect 27813 13277 27847 13311
rect 27997 13277 28031 13311
rect 29653 13277 29687 13311
rect 31401 13277 31435 13311
rect 32597 13277 32631 13311
rect 36369 13277 36403 13311
rect 37933 13277 37967 13311
rect 39589 13277 39623 13311
rect 39865 13277 39899 13311
rect 44557 13277 44591 13311
rect 46213 13277 46247 13311
rect 47225 13277 47259 13311
rect 47961 13277 47995 13311
rect 50721 13277 50755 13311
rect 56609 13277 56643 13311
rect 57897 13277 57931 13311
rect 6276 13209 6310 13243
rect 9229 13209 9263 13243
rect 14473 13209 14507 13243
rect 15209 13209 15243 13243
rect 27568 13209 27602 13243
rect 28264 13209 28298 13243
rect 29920 13209 29954 13243
rect 32045 13209 32079 13243
rect 32864 13209 32898 13243
rect 34980 13209 35014 13243
rect 36636 13209 36670 13243
rect 38200 13209 38234 13243
rect 41972 13209 42006 13243
rect 44312 13209 44346 13243
rect 2973 13141 3007 13175
rect 8125 13141 8159 13175
rect 10149 13141 10183 13175
rect 13461 13141 13495 13175
rect 14105 13141 14139 13175
rect 15761 13141 15795 13175
rect 17233 13141 17267 13175
rect 19073 13141 19107 13175
rect 21557 13141 21591 13175
rect 22201 13141 22235 13175
rect 24501 13141 24535 13175
rect 29377 13141 29411 13175
rect 32137 13141 32171 13175
rect 34345 13141 34379 13175
rect 36093 13141 36127 13175
rect 37749 13141 37783 13175
rect 39313 13141 39347 13175
rect 41337 13141 41371 13175
rect 43177 13141 43211 13175
rect 45293 13141 45327 13175
rect 45385 13141 45419 13175
rect 45753 13141 45787 13175
rect 46305 13141 46339 13175
rect 47409 13141 47443 13175
rect 50445 13141 50479 13175
rect 56701 13141 56735 13175
rect 6929 12937 6963 12971
rect 12265 12937 12299 12971
rect 13093 12937 13127 12971
rect 13461 12937 13495 12971
rect 13737 12937 13771 12971
rect 14013 12937 14047 12971
rect 18521 12937 18555 12971
rect 21465 12937 21499 12971
rect 24225 12937 24259 12971
rect 25329 12937 25363 12971
rect 26985 12937 27019 12971
rect 27997 12937 28031 12971
rect 30665 12937 30699 12971
rect 32321 12937 32355 12971
rect 32873 12937 32907 12971
rect 33241 12937 33275 12971
rect 33977 12937 34011 12971
rect 35173 12937 35207 12971
rect 36921 12937 36955 12971
rect 38485 12937 38519 12971
rect 41429 12937 41463 12971
rect 42165 12937 42199 12971
rect 42625 12937 42659 12971
rect 43269 12937 43303 12971
rect 43361 12937 43395 12971
rect 45385 12937 45419 12971
rect 47133 12937 47167 12971
rect 50077 12937 50111 12971
rect 55045 12937 55079 12971
rect 55505 12937 55539 12971
rect 2964 12869 2998 12903
rect 7021 12869 7055 12903
rect 15117 12869 15151 12903
rect 15577 12869 15611 12903
rect 19993 12869 20027 12903
rect 30573 12869 30607 12903
rect 33333 12869 33367 12903
rect 36645 12869 36679 12903
rect 37565 12869 37599 12903
rect 39212 12869 39246 12903
rect 40785 12869 40819 12903
rect 43913 12869 43947 12903
rect 46020 12869 46054 12903
rect 58265 12869 58299 12903
rect 12633 12801 12667 12835
rect 13921 12801 13955 12835
rect 14565 12801 14599 12835
rect 16129 12801 16163 12835
rect 16773 12801 16807 12835
rect 17040 12801 17074 12835
rect 20085 12801 20119 12835
rect 20352 12801 20386 12835
rect 22385 12801 22419 12835
rect 22652 12801 22686 12835
rect 24317 12801 24351 12835
rect 25688 12801 25722 12835
rect 27905 12801 27939 12835
rect 28181 12801 28215 12835
rect 29377 12801 29411 12835
rect 29469 12801 29503 12835
rect 31033 12801 31067 12835
rect 35725 12801 35759 12835
rect 36001 12801 36035 12835
rect 38117 12801 38151 12835
rect 38945 12801 38979 12835
rect 41797 12801 41831 12835
rect 45753 12801 45787 12835
rect 50261 12801 50295 12835
rect 50528 12801 50562 12835
rect 56977 12801 57011 12835
rect 58449 12801 58483 12835
rect 2697 12733 2731 12767
rect 4169 12733 4203 12767
rect 7205 12733 7239 12767
rect 7941 12733 7975 12767
rect 15209 12733 15243 12767
rect 15301 12733 15335 12767
rect 24409 12733 24443 12767
rect 24685 12733 24719 12767
rect 25421 12733 25455 12767
rect 27537 12733 27571 12767
rect 29653 12733 29687 12767
rect 30849 12733 30883 12767
rect 33517 12733 33551 12767
rect 40877 12733 40911 12767
rect 40969 12733 41003 12767
rect 43085 12733 43119 12767
rect 48329 12733 48363 12767
rect 54677 12733 54711 12767
rect 55965 12733 55999 12767
rect 57069 12733 57103 12767
rect 57161 12733 57195 12767
rect 57621 12733 57655 12767
rect 4077 12665 4111 12699
rect 5365 12665 5399 12699
rect 7665 12665 7699 12699
rect 23765 12665 23799 12699
rect 26801 12665 26835 12699
rect 31677 12665 31711 12699
rect 56609 12665 56643 12699
rect 4813 12597 4847 12631
rect 6561 12597 6595 12631
rect 10057 12597 10091 12631
rect 14749 12597 14783 12631
rect 18153 12597 18187 12631
rect 23857 12597 23891 12631
rect 28825 12597 28859 12631
rect 29009 12597 29043 12631
rect 30021 12597 30055 12631
rect 30205 12597 30239 12631
rect 32689 12597 32723 12631
rect 40325 12597 40359 12631
rect 40417 12597 40451 12631
rect 43729 12597 43763 12631
rect 47777 12597 47811 12631
rect 51641 12597 51675 12631
rect 54125 12597 54159 12631
rect 56517 12597 56551 12631
rect 6469 12393 6503 12427
rect 10609 12393 10643 12427
rect 15853 12393 15887 12427
rect 16681 12393 16715 12427
rect 17601 12393 17635 12427
rect 19809 12393 19843 12427
rect 21005 12393 21039 12427
rect 21557 12393 21591 12427
rect 23305 12393 23339 12427
rect 24869 12393 24903 12427
rect 26617 12393 26651 12427
rect 28641 12393 28675 12427
rect 29745 12393 29779 12427
rect 30113 12393 30147 12427
rect 40509 12393 40543 12427
rect 42349 12393 42383 12427
rect 43085 12393 43119 12427
rect 44741 12393 44775 12427
rect 45569 12393 45603 12427
rect 46029 12393 46063 12427
rect 50721 12393 50755 12427
rect 52009 12393 52043 12427
rect 53941 12393 53975 12427
rect 54125 12393 54159 12427
rect 5181 12325 5215 12359
rect 18337 12325 18371 12359
rect 21373 12325 21407 12359
rect 47041 12325 47075 12359
rect 48697 12325 48731 12359
rect 50629 12325 50663 12359
rect 57805 12325 57839 12359
rect 2973 12257 3007 12291
rect 5825 12257 5859 12291
rect 7021 12257 7055 12291
rect 8125 12257 8159 12291
rect 10333 12257 10367 12291
rect 18245 12257 18279 12291
rect 18889 12257 18923 12291
rect 20545 12257 20579 12291
rect 22109 12257 22143 12291
rect 23857 12257 23891 12291
rect 25513 12257 25547 12291
rect 25881 12257 25915 12291
rect 26065 12257 26099 12291
rect 29193 12257 29227 12291
rect 30665 12257 30699 12291
rect 39865 12257 39899 12291
rect 41153 12257 41187 12291
rect 42901 12257 42935 12291
rect 43637 12257 43671 12291
rect 44097 12257 44131 12291
rect 47317 12257 47351 12291
rect 49341 12257 49375 12291
rect 51273 12257 51307 12291
rect 54677 12257 54711 12291
rect 58449 12257 58483 12291
rect 3249 12189 3283 12223
rect 3525 12189 3559 12223
rect 3801 12189 3835 12223
rect 7481 12189 7515 12223
rect 10793 12189 10827 12223
rect 12725 12189 12759 12223
rect 14197 12189 14231 12223
rect 14464 12189 14498 12223
rect 17049 12189 17083 12223
rect 18705 12189 18739 12223
rect 20361 12189 20395 12223
rect 25329 12189 25363 12223
rect 27169 12189 27203 12223
rect 37473 12189 37507 12223
rect 40601 12189 40635 12223
rect 45201 12189 45235 12223
rect 46305 12189 46339 12223
rect 46857 12189 46891 12223
rect 47225 12189 47259 12223
rect 51089 12189 51123 12223
rect 52653 12189 52687 12223
rect 55321 12189 55355 12223
rect 56425 12189 56459 12223
rect 56692 12189 56726 12223
rect 2728 12121 2762 12155
rect 4068 12121 4102 12155
rect 10885 12121 10919 12155
rect 13553 12121 13587 12155
rect 15761 12121 15795 12155
rect 18797 12121 18831 12155
rect 20913 12121 20947 12155
rect 47584 12121 47618 12155
rect 52101 12121 52135 12155
rect 54493 12121 54527 12155
rect 55965 12121 55999 12155
rect 1593 12053 1627 12087
rect 3065 12053 3099 12087
rect 3433 12053 3467 12087
rect 5273 12053 5307 12087
rect 7573 12053 7607 12087
rect 8585 12053 8619 12087
rect 9781 12053 9815 12087
rect 12173 12053 12207 12087
rect 15577 12053 15611 12087
rect 16865 12053 16899 12087
rect 19901 12053 19935 12087
rect 20269 12053 20303 12087
rect 24961 12053 24995 12087
rect 25421 12053 25455 12087
rect 26157 12053 26191 12087
rect 26525 12053 26559 12087
rect 27629 12053 27663 12087
rect 31125 12053 31159 12087
rect 36001 12053 36035 12087
rect 37105 12053 37139 12087
rect 42165 12053 42199 12087
rect 48789 12053 48823 12087
rect 51181 12053 51215 12087
rect 53297 12053 53331 12087
rect 54585 12053 54619 12087
rect 57897 12053 57931 12087
rect 2973 11849 3007 11883
rect 3893 11849 3927 11883
rect 4261 11849 4295 11883
rect 19809 11849 19843 11883
rect 23765 11849 23799 11883
rect 28917 11849 28951 11883
rect 34989 11849 35023 11883
rect 38209 11849 38243 11883
rect 41429 11849 41463 11883
rect 43361 11849 43395 11883
rect 44097 11849 44131 11883
rect 46765 11849 46799 11883
rect 47593 11849 47627 11883
rect 49065 11849 49099 11883
rect 55137 11849 55171 11883
rect 24584 11781 24618 11815
rect 29837 11781 29871 11815
rect 35449 11781 35483 11815
rect 54024 11781 54058 11815
rect 2237 11713 2271 11747
rect 3525 11713 3559 11747
rect 4997 11713 5031 11747
rect 7490 11713 7524 11747
rect 7757 11713 7791 11747
rect 8677 11713 8711 11747
rect 11345 11713 11379 11747
rect 11785 11713 11819 11747
rect 13093 11713 13127 11747
rect 13645 11713 13679 11747
rect 15117 11713 15151 11747
rect 15393 11713 15427 11747
rect 18521 11713 18555 11747
rect 20361 11713 20395 11747
rect 21189 11713 21223 11747
rect 29193 11713 29227 11747
rect 35081 11713 35115 11747
rect 38117 11713 38151 11747
rect 46949 11713 46983 11747
rect 48717 11713 48751 11747
rect 48973 11713 49007 11747
rect 50445 11713 50479 11747
rect 51181 11713 51215 11747
rect 56195 11713 56229 11747
rect 57253 11713 57287 11747
rect 58541 11713 58575 11747
rect 4813 11645 4847 11679
rect 5089 11645 5123 11679
rect 7941 11645 7975 11679
rect 9045 11645 9079 11679
rect 9965 11645 9999 11679
rect 11529 11645 11563 11679
rect 17509 11645 17543 11679
rect 19165 11645 19199 11679
rect 24317 11645 24351 11679
rect 28457 11645 28491 11679
rect 30205 11645 30239 11679
rect 31585 11645 31619 11679
rect 33609 11645 33643 11679
rect 33793 11645 33827 11679
rect 34805 11645 34839 11679
rect 36185 11645 36219 11679
rect 36369 11645 36403 11679
rect 37841 11645 37875 11679
rect 40877 11645 40911 11679
rect 42993 11645 43027 11679
rect 45661 11645 45695 11679
rect 45937 11645 45971 11679
rect 49617 11645 49651 11679
rect 52469 11645 52503 11679
rect 53297 11645 53331 11679
rect 53757 11645 53791 11679
rect 56057 11645 56091 11679
rect 56333 11645 56367 11679
rect 57069 11645 57103 11679
rect 32413 11577 32447 11611
rect 32781 11577 32815 11611
rect 37289 11577 37323 11611
rect 47133 11577 47167 11611
rect 56609 11577 56643 11611
rect 2881 11509 2915 11543
rect 4997 11509 5031 11543
rect 5365 11509 5399 11543
rect 6377 11509 6411 11543
rect 8585 11509 8619 11543
rect 10609 11509 10643 11543
rect 10977 11509 11011 11543
rect 11161 11509 11195 11543
rect 12909 11509 12943 11543
rect 14105 11509 14139 11543
rect 14657 11509 14691 11543
rect 16957 11509 16991 11543
rect 18245 11509 18279 11543
rect 20545 11509 20579 11543
rect 25697 11509 25731 11543
rect 25973 11509 26007 11543
rect 28089 11509 28123 11543
rect 29009 11509 29043 11543
rect 30849 11509 30883 11543
rect 31033 11509 31067 11543
rect 33057 11509 33091 11543
rect 34437 11509 34471 11543
rect 35633 11509 35667 11543
rect 37013 11509 37047 11543
rect 40325 11509 40359 11543
rect 42441 11509 42475 11543
rect 43729 11509 43763 11543
rect 45109 11509 45143 11543
rect 46489 11509 46523 11543
rect 50261 11509 50295 11543
rect 50997 11509 51031 11543
rect 51917 11509 51951 11543
rect 52745 11509 52779 11543
rect 55413 11509 55447 11543
rect 58357 11509 58391 11543
rect 4353 11305 4387 11339
rect 8033 11305 8067 11339
rect 8953 11305 8987 11339
rect 13921 11305 13955 11339
rect 18429 11305 18463 11339
rect 24869 11305 24903 11339
rect 26801 11305 26835 11339
rect 29929 11305 29963 11339
rect 30113 11305 30147 11339
rect 37565 11305 37599 11339
rect 41245 11305 41279 11339
rect 44465 11305 44499 11339
rect 45201 11305 45235 11339
rect 46305 11305 46339 11339
rect 49157 11305 49191 11339
rect 50721 11305 50755 11339
rect 52377 11305 52411 11339
rect 52469 11305 52503 11339
rect 53481 11305 53515 11339
rect 2329 11237 2363 11271
rect 17417 11237 17451 11271
rect 28641 11237 28675 11271
rect 35265 11237 35299 11271
rect 37473 11237 37507 11271
rect 43453 11237 43487 11271
rect 47685 11237 47719 11271
rect 49249 11237 49283 11271
rect 57621 11237 57655 11271
rect 7297 11169 7331 11203
rect 7481 11169 7515 11203
rect 8585 11169 8619 11203
rect 11621 11169 11655 11203
rect 12081 11169 12115 11203
rect 16589 11169 16623 11203
rect 16773 11169 16807 11203
rect 17509 11169 17543 11203
rect 23581 11169 23615 11203
rect 28549 11169 28583 11203
rect 29193 11169 29227 11203
rect 30757 11169 30791 11203
rect 31677 11169 31711 11203
rect 33609 11169 33643 11203
rect 35817 11169 35851 11203
rect 38117 11169 38151 11203
rect 39865 11169 39899 11203
rect 42073 11169 42107 11203
rect 45845 11169 45879 11203
rect 47135 11169 47169 11203
rect 48329 11169 48363 11203
rect 48605 11169 48639 11203
rect 52929 11169 52963 11203
rect 53113 11169 53147 11203
rect 53757 11169 53791 11203
rect 56241 11169 56275 11203
rect 2513 11101 2547 11135
rect 2789 11101 2823 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 3157 11101 3191 11135
rect 3249 11101 3283 11135
rect 3821 11101 3855 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4169 11101 4203 11135
rect 4445 11101 4479 11135
rect 4629 11101 4663 11135
rect 7205 11101 7239 11135
rect 8401 11101 8435 11135
rect 10333 11101 10367 11135
rect 11069 11101 11103 11135
rect 11207 11101 11241 11135
rect 11345 11101 11379 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 13185 11101 13219 11135
rect 15209 11101 15243 11135
rect 20361 11101 20395 11135
rect 21189 11101 21223 11135
rect 21465 11101 21499 11135
rect 22201 11101 22235 11135
rect 25697 11101 25731 11135
rect 27813 11101 27847 11135
rect 30941 11101 30975 11135
rect 33793 11101 33827 11135
rect 36093 11101 36127 11135
rect 39037 11101 39071 11135
rect 41337 11101 41371 11135
rect 44097 11101 44131 11135
rect 45569 11101 45603 11135
rect 47271 11101 47305 11135
rect 47409 11101 47443 11135
rect 48145 11101 48179 11135
rect 48789 11101 48823 11135
rect 49801 11101 49835 11135
rect 50997 11101 51031 11135
rect 55873 11101 55907 11135
rect 58265 11101 58299 11135
rect 2697 11033 2731 11067
rect 7849 11033 7883 11067
rect 8493 11033 8527 11067
rect 10088 11033 10122 11067
rect 10425 11033 10459 11067
rect 16957 11033 16991 11067
rect 19809 11033 19843 11067
rect 22753 11033 22787 11067
rect 26709 11033 26743 11067
rect 27905 11033 27939 11067
rect 29101 11033 29135 11067
rect 30481 11033 30515 11067
rect 30573 11033 30607 11067
rect 33364 11033 33398 11067
rect 34345 11033 34379 11067
rect 34897 11033 34931 11067
rect 35633 11033 35667 11067
rect 36360 11033 36394 11067
rect 38393 11033 38427 11067
rect 40132 11033 40166 11067
rect 42340 11033 42374 11067
rect 46489 11033 46523 11067
rect 51264 11033 51298 11067
rect 54024 11033 54058 11067
rect 55321 11033 55355 11067
rect 56508 11033 56542 11067
rect 57713 11033 57747 11067
rect 3433 10965 3467 10999
rect 4445 10965 4479 10999
rect 6837 10965 6871 10999
rect 14381 10965 14415 10999
rect 14565 10965 14599 10999
rect 17049 10965 17083 10999
rect 18153 10965 18187 10999
rect 20637 10965 20671 10999
rect 22017 10965 22051 10999
rect 22937 10965 22971 10999
rect 23857 10965 23891 10999
rect 27169 10965 27203 10999
rect 29009 10965 29043 10999
rect 32229 10965 32263 10999
rect 35725 10965 35759 10999
rect 37933 10965 37967 10999
rect 38025 10965 38059 10999
rect 39313 10965 39347 10999
rect 41981 10965 42015 10999
rect 43545 10965 43579 10999
rect 45661 10965 45695 10999
rect 48697 10965 48731 10999
rect 52837 10965 52871 10999
rect 55137 10965 55171 10999
rect 2789 10761 2823 10795
rect 2881 10761 2915 10795
rect 3893 10761 3927 10795
rect 4169 10761 4203 10795
rect 4261 10761 4295 10795
rect 7389 10761 7423 10795
rect 7757 10761 7791 10795
rect 10241 10761 10275 10795
rect 14473 10761 14507 10795
rect 14657 10761 14691 10795
rect 16681 10761 16715 10795
rect 19533 10761 19567 10795
rect 19901 10761 19935 10795
rect 21649 10761 21683 10795
rect 26341 10761 26375 10795
rect 33609 10761 33643 10795
rect 34069 10761 34103 10795
rect 36185 10761 36219 10795
rect 36645 10761 36679 10795
rect 39221 10761 39255 10795
rect 40785 10761 40819 10795
rect 40877 10761 40911 10795
rect 41981 10761 42015 10795
rect 43913 10761 43947 10795
rect 46029 10761 46063 10795
rect 47869 10761 47903 10795
rect 47961 10761 47995 10795
rect 49709 10761 49743 10795
rect 55045 10761 55079 10795
rect 56977 10761 57011 10795
rect 57345 10761 57379 10795
rect 8300 10693 8334 10727
rect 10333 10693 10367 10727
rect 13645 10693 13679 10727
rect 15761 10693 15795 10727
rect 30389 10693 30423 10727
rect 30757 10693 30791 10727
rect 32404 10693 32438 10727
rect 34980 10693 35014 10727
rect 36553 10693 36587 10727
rect 39672 10693 39706 10727
rect 42708 10693 42742 10727
rect 44916 10693 44950 10727
rect 46581 10693 46615 10727
rect 48605 10693 48639 10727
rect 51448 10693 51482 10727
rect 54585 10693 54619 10727
rect 55781 10693 55815 10727
rect 57897 10693 57931 10727
rect 2605 10625 2639 10659
rect 2789 10625 2823 10659
rect 3065 10625 3099 10659
rect 3249 10625 3283 10659
rect 3525 10625 3559 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 6837 10625 6871 10659
rect 11796 10625 11830 10659
rect 13553 10625 13587 10659
rect 15025 10625 15059 10659
rect 15117 10625 15151 10659
rect 16497 10625 16531 10659
rect 17805 10625 17839 10659
rect 18061 10625 18095 10659
rect 20269 10625 20303 10659
rect 20536 10625 20570 10659
rect 22109 10625 22143 10659
rect 22376 10625 22410 10659
rect 24225 10625 24259 10659
rect 26249 10625 26283 10659
rect 27425 10625 27459 10659
rect 28641 10625 28675 10659
rect 30941 10625 30975 10659
rect 32137 10625 32171 10659
rect 33977 10625 34011 10659
rect 34713 10625 34747 10659
rect 37740 10625 37774 10659
rect 39405 10625 39439 10659
rect 41245 10625 41279 10659
rect 42441 10625 42475 10659
rect 44649 10625 44683 10659
rect 46489 10625 46523 10659
rect 49433 10625 49467 10659
rect 49893 10625 49927 10659
rect 51181 10625 51215 10659
rect 53113 10625 53147 10659
rect 53573 10625 53607 10659
rect 54677 10625 54711 10659
rect 56885 10625 56919 10659
rect 58449 10625 58483 10659
rect 3433 10557 3467 10591
rect 3617 10557 3651 10591
rect 8033 10557 8067 10591
rect 10149 10557 10183 10591
rect 11529 10557 11563 10591
rect 13737 10557 13771 10591
rect 15209 10557 15243 10591
rect 15853 10557 15887 10591
rect 18705 10557 18739 10591
rect 19257 10557 19291 10591
rect 19441 10557 19475 10591
rect 23765 10557 23799 10591
rect 25789 10557 25823 10591
rect 26433 10557 26467 10591
rect 27169 10557 27203 10591
rect 31309 10557 31343 10591
rect 34161 10557 34195 10591
rect 36737 10557 36771 10591
rect 37473 10557 37507 10591
rect 41337 10557 41371 10591
rect 41521 10557 41555 10591
rect 44465 10557 44499 10591
rect 46673 10557 46707 10591
rect 47133 10557 47167 10591
rect 47777 10557 47811 10591
rect 48973 10557 49007 10591
rect 50261 10557 50295 10591
rect 53205 10557 53239 10591
rect 53389 10557 53423 10591
rect 54125 10557 54159 10591
rect 54493 10557 54527 10591
rect 55229 10557 55263 10591
rect 56517 10557 56551 10591
rect 56793 10557 56827 10591
rect 9873 10489 9907 10523
rect 24041 10489 24075 10523
rect 25881 10489 25915 10523
rect 33517 10489 33551 10523
rect 36093 10489 36127 10523
rect 48329 10489 48363 10523
rect 52561 10489 52595 10523
rect 6561 10421 6595 10455
rect 9413 10421 9447 10455
rect 10701 10421 10735 10455
rect 11345 10421 11379 10455
rect 12909 10421 12943 10455
rect 13185 10421 13219 10455
rect 18153 10421 18187 10455
rect 23489 10421 23523 10455
rect 25145 10421 25179 10455
rect 28549 10421 28583 10455
rect 38853 10421 38887 10455
rect 43821 10421 43855 10455
rect 46121 10421 46155 10455
rect 50813 10421 50847 10455
rect 52745 10421 52779 10455
rect 3157 10217 3191 10251
rect 3433 10217 3467 10251
rect 4537 10217 4571 10251
rect 8769 10217 8803 10251
rect 10149 10217 10183 10251
rect 10425 10217 10459 10251
rect 12541 10217 12575 10251
rect 15485 10217 15519 10251
rect 18521 10217 18555 10251
rect 21465 10217 21499 10251
rect 29837 10217 29871 10251
rect 31401 10217 31435 10251
rect 34437 10217 34471 10251
rect 43913 10217 43947 10251
rect 47685 10217 47719 10251
rect 47961 10217 47995 10251
rect 49157 10217 49191 10251
rect 50261 10217 50295 10251
rect 54217 10217 54251 10251
rect 56333 10217 56367 10251
rect 5365 10149 5399 10183
rect 7021 10149 7055 10183
rect 8953 10149 8987 10183
rect 24225 10149 24259 10183
rect 32689 10149 32723 10183
rect 46673 10149 46707 10183
rect 53297 10149 53331 10183
rect 3249 10081 3283 10115
rect 7113 10081 7147 10115
rect 9505 10081 9539 10115
rect 9965 10081 9999 10115
rect 10977 10081 11011 10115
rect 11897 10081 11931 10115
rect 11989 10081 12023 10115
rect 13185 10081 13219 10115
rect 13829 10081 13863 10115
rect 16497 10081 16531 10115
rect 16773 10081 16807 10115
rect 17049 10081 17083 10115
rect 17693 10081 17727 10115
rect 17969 10081 18003 10115
rect 22477 10081 22511 10115
rect 22753 10081 22787 10115
rect 23213 10081 23247 10115
rect 23673 10081 23707 10115
rect 24961 10081 24995 10115
rect 27813 10081 27847 10115
rect 28089 10081 28123 10115
rect 28549 10081 28583 10115
rect 29377 10081 29411 10115
rect 30021 10081 30055 10115
rect 32275 10081 32309 10115
rect 32413 10081 32447 10115
rect 33609 10081 33643 10115
rect 33701 10081 33735 10115
rect 37059 10081 37093 10115
rect 37473 10081 37507 10115
rect 38117 10081 38151 10115
rect 38301 10081 38335 10115
rect 38485 10081 38519 10115
rect 39589 10081 39623 10115
rect 40693 10081 40727 10115
rect 40785 10081 40819 10115
rect 42027 10081 42061 10115
rect 42165 10081 42199 10115
rect 42441 10081 42475 10115
rect 43269 10081 43303 10115
rect 44557 10081 44591 10115
rect 45293 10081 45327 10115
rect 47041 10081 47075 10115
rect 50813 10081 50847 10115
rect 52009 10081 52043 10115
rect 52285 10081 52319 10115
rect 52745 10081 52779 10115
rect 57529 10081 57563 10115
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 5824 10013 5858 10047
rect 5917 10013 5951 10047
rect 6284 10013 6318 10047
rect 6377 10013 6411 10047
rect 6892 10013 6926 10047
rect 10333 10013 10367 10047
rect 11805 10013 11839 10047
rect 13277 10013 13311 10047
rect 14105 10013 14139 10047
rect 16635 10013 16669 10047
rect 17509 10013 17543 10047
rect 18061 10013 18095 10047
rect 19441 10013 19475 10047
rect 22201 10013 22235 10047
rect 22339 10013 22373 10047
rect 23397 10013 23431 10047
rect 23857 10013 23891 10047
rect 25237 10013 25271 10047
rect 27537 10013 27571 10047
rect 27696 10013 27730 10047
rect 28733 10013 28767 10047
rect 30288 10013 30322 10047
rect 32137 10013 32171 10047
rect 33149 10013 33183 10047
rect 33333 10013 33367 10047
rect 34713 10013 34747 10047
rect 36921 10013 36955 10047
rect 37197 10013 37231 10047
rect 37933 10013 37967 10047
rect 40049 10013 40083 10047
rect 41889 10013 41923 10047
rect 42901 10013 42935 10047
rect 43085 10013 43119 10047
rect 49433 10013 49467 10047
rect 50629 10013 50663 10047
rect 51733 10013 51767 10047
rect 51892 10013 51926 10047
rect 52929 10013 52963 10047
rect 3065 9945 3099 9979
rect 6009 9945 6043 9979
rect 6745 9945 6779 9979
rect 7481 9945 7515 9979
rect 14372 9945 14406 9979
rect 19708 9945 19742 9979
rect 23765 9945 23799 9979
rect 25482 9945 25516 9979
rect 33793 9945 33827 9979
rect 34980 9945 35014 9979
rect 38577 9945 38611 9979
rect 39037 9945 39071 9979
rect 40601 9945 40635 9979
rect 43545 9945 43579 9979
rect 44005 9945 44039 9979
rect 45560 9945 45594 9979
rect 49985 9945 50019 9979
rect 50721 9945 50755 9979
rect 7849 9877 7883 9911
rect 11437 9877 11471 9911
rect 15853 9877 15887 9911
rect 18153 9877 18187 9911
rect 18981 9877 19015 9911
rect 20821 9877 20855 9911
rect 21557 9877 21591 9911
rect 24409 9877 24443 9911
rect 26617 9877 26651 9911
rect 26893 9877 26927 9911
rect 31493 9877 31527 9911
rect 34161 9877 34195 9911
rect 36093 9877 36127 9911
rect 36277 9877 36311 9911
rect 38945 9877 38979 9911
rect 40233 9877 40267 9911
rect 41245 9877 41279 9911
rect 43453 9877 43487 9911
rect 51089 9877 51123 9911
rect 56977 9877 57011 9911
rect 3341 9673 3375 9707
rect 6101 9673 6135 9707
rect 11805 9673 11839 9707
rect 13277 9673 13311 9707
rect 15761 9673 15795 9707
rect 22385 9673 22419 9707
rect 31953 9673 31987 9707
rect 33701 9673 33735 9707
rect 35265 9673 35299 9707
rect 36645 9673 36679 9707
rect 38485 9673 38519 9707
rect 38577 9673 38611 9707
rect 42809 9673 42843 9707
rect 45109 9673 45143 9707
rect 45845 9673 45879 9707
rect 49709 9673 49743 9707
rect 54217 9673 54251 9707
rect 56885 9673 56919 9707
rect 7757 9605 7791 9639
rect 11345 9605 11379 9639
rect 12541 9605 12575 9639
rect 15669 9605 15703 9639
rect 17816 9605 17850 9639
rect 19656 9605 19690 9639
rect 20453 9605 20487 9639
rect 23520 9605 23554 9639
rect 27261 9605 27295 9639
rect 33793 9605 33827 9639
rect 40233 9605 40267 9639
rect 42257 9605 42291 9639
rect 42717 9605 42751 9639
rect 43361 9605 43395 9639
rect 46765 9605 46799 9639
rect 50822 9605 50856 9639
rect 51549 9605 51583 9639
rect 52745 9605 52779 9639
rect 3249 9537 3283 9571
rect 6469 9537 6503 9571
rect 6745 9537 6779 9571
rect 7113 9537 7147 9571
rect 7849 9537 7883 9571
rect 9873 9537 9907 9571
rect 10793 9537 10827 9571
rect 12725 9537 12759 9571
rect 14096 9537 14130 9571
rect 16313 9537 16347 9571
rect 21281 9537 21315 9571
rect 21373 9537 21407 9571
rect 22109 9537 22143 9571
rect 24501 9537 24535 9571
rect 25053 9537 25087 9571
rect 25320 9537 25354 9571
rect 27629 9537 27663 9571
rect 27896 9537 27930 9571
rect 29101 9537 29135 9571
rect 29837 9537 29871 9571
rect 30104 9537 30138 9571
rect 32137 9537 32171 9571
rect 33057 9537 33091 9571
rect 34345 9537 34379 9571
rect 34529 9537 34563 9571
rect 35173 9537 35207 9571
rect 35909 9537 35943 9571
rect 36093 9537 36127 9571
rect 37841 9537 37875 9571
rect 39129 9537 39163 9571
rect 40785 9537 40819 9571
rect 43913 9537 43947 9571
rect 46397 9537 46431 9571
rect 52285 9537 52319 9571
rect 54309 9537 54343 9571
rect 56149 9537 56183 9571
rect 8033 9469 8067 9503
rect 9413 9469 9447 9503
rect 9965 9469 9999 9503
rect 11897 9469 11931 9503
rect 13829 9469 13863 9503
rect 15945 9469 15979 9503
rect 18061 9469 18095 9503
rect 19901 9469 19935 9503
rect 20545 9469 20579 9503
rect 20637 9469 20671 9503
rect 21557 9469 21591 9503
rect 23765 9469 23799 9503
rect 29653 9469 29687 9503
rect 31309 9469 31343 9503
rect 32689 9469 32723 9503
rect 42625 9469 42659 9503
rect 48145 9469 48179 9503
rect 51089 9469 51123 9503
rect 51273 9469 51307 9503
rect 51457 9469 51491 9503
rect 53297 9469 53331 9503
rect 54033 9469 54067 9503
rect 55321 9469 55355 9503
rect 55505 9469 55539 9503
rect 56977 9469 57011 9503
rect 57069 9469 57103 9503
rect 15209 9401 15243 9435
rect 29009 9401 29043 9435
rect 31217 9401 31251 9435
rect 43177 9401 43211 9435
rect 54677 9401 54711 9435
rect 8769 9333 8803 9367
rect 8861 9333 8895 9367
rect 9689 9333 9723 9367
rect 10609 9333 10643 9367
rect 13737 9333 13771 9367
rect 15301 9333 15335 9367
rect 16681 9333 16715 9367
rect 18337 9333 18371 9367
rect 18521 9333 18555 9367
rect 20085 9333 20119 9367
rect 20913 9333 20947 9367
rect 23857 9333 23891 9367
rect 26433 9333 26467 9367
rect 26709 9333 26743 9367
rect 36921 9333 36955 9367
rect 37565 9333 37599 9367
rect 41153 9333 41187 9367
rect 41613 9333 41647 9367
rect 47225 9333 47259 9367
rect 48053 9333 48087 9367
rect 48789 9333 48823 9367
rect 51917 9333 51951 9367
rect 53849 9333 53883 9367
rect 54769 9333 54803 9367
rect 56517 9333 56551 9367
rect 3157 9129 3191 9163
rect 3525 9129 3559 9163
rect 5825 9129 5859 9163
rect 6561 9129 6595 9163
rect 7021 9129 7055 9163
rect 7849 9129 7883 9163
rect 10701 9129 10735 9163
rect 14749 9129 14783 9163
rect 16129 9129 16163 9163
rect 18153 9129 18187 9163
rect 18521 9129 18555 9163
rect 21373 9129 21407 9163
rect 22385 9129 22419 9163
rect 23305 9129 23339 9163
rect 23857 9129 23891 9163
rect 27721 9129 27755 9163
rect 29745 9129 29779 9163
rect 30113 9129 30147 9163
rect 31309 9129 31343 9163
rect 34437 9129 34471 9163
rect 34897 9129 34931 9163
rect 36277 9129 36311 9163
rect 38209 9129 38243 9163
rect 38485 9129 38519 9163
rect 55597 9129 55631 9163
rect 56333 9129 56367 9163
rect 3893 9061 3927 9095
rect 6193 9061 6227 9095
rect 6653 9061 6687 9095
rect 7481 9061 7515 9095
rect 8677 9061 8711 9095
rect 19901 9061 19935 9095
rect 43085 9061 43119 9095
rect 51549 9061 51583 9095
rect 2697 8993 2731 9027
rect 4261 8993 4295 9027
rect 4629 8993 4663 9027
rect 6745 8993 6779 9027
rect 8309 8993 8343 9027
rect 12081 8993 12115 9027
rect 13737 8993 13771 9027
rect 14289 8993 14323 9027
rect 15393 8993 15427 9027
rect 15577 8993 15611 9027
rect 17509 8993 17543 9027
rect 20453 8993 20487 9027
rect 20821 8993 20855 9027
rect 21741 8993 21775 9027
rect 22661 8993 22695 9027
rect 22845 8993 22879 9027
rect 26341 8993 26375 9027
rect 26985 8993 27019 9027
rect 27629 8993 27663 9027
rect 28273 8993 28307 9027
rect 28549 8993 28583 9027
rect 30757 8993 30791 9027
rect 31677 8993 31711 9027
rect 32781 8993 32815 9027
rect 35909 8993 35943 9027
rect 47041 8993 47075 9027
rect 48145 8993 48179 9027
rect 48513 8993 48547 9027
rect 50169 8993 50203 9027
rect 52193 8993 52227 9027
rect 55781 8993 55815 9027
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 6101 8925 6135 8959
rect 8401 8925 8435 8959
rect 9045 8925 9079 8959
rect 10057 8925 10091 8959
rect 12633 8925 12667 8959
rect 25145 8925 25179 8959
rect 26157 8925 26191 8959
rect 28181 8925 28215 8959
rect 29193 8925 29227 8959
rect 30849 8925 30883 8959
rect 32965 8925 32999 8959
rect 36369 8925 36403 8959
rect 37197 8925 37231 8959
rect 38945 8925 38979 8959
rect 45937 8925 45971 8959
rect 48605 8925 48639 8959
rect 49709 8925 49743 8959
rect 56425 8925 56459 8959
rect 57897 8925 57931 8959
rect 58449 8925 58483 8959
rect 3525 8857 3559 8891
rect 5457 8857 5491 8891
rect 7757 8857 7791 8891
rect 8677 8857 8711 8891
rect 9597 8857 9631 8891
rect 10609 8857 10643 8891
rect 11814 8857 11848 8891
rect 13277 8857 13311 8891
rect 19717 8857 19751 8891
rect 24869 8857 24903 8891
rect 26893 8857 26927 8891
rect 30941 8857 30975 8891
rect 38577 8857 38611 8891
rect 47317 8857 47351 8891
rect 48697 8857 48731 8891
rect 50436 8857 50470 8891
rect 51641 8857 51675 8891
rect 53389 8857 53423 8891
rect 55137 8857 55171 8891
rect 56692 8857 56726 8891
rect 3801 8789 3835 8823
rect 5834 8789 5868 8823
rect 8493 8789 8527 8823
rect 22937 8789 22971 8823
rect 25697 8789 25731 8823
rect 25789 8789 25823 8823
rect 26249 8789 26283 8823
rect 28089 8789 28123 8823
rect 32873 8789 32907 8823
rect 33333 8789 33367 8823
rect 33609 8789 33643 8823
rect 34069 8789 34103 8823
rect 35265 8789 35299 8823
rect 37013 8789 37047 8823
rect 37841 8789 37875 8823
rect 45385 8789 45419 8823
rect 46305 8789 46339 8823
rect 46489 8789 46523 8823
rect 49065 8789 49099 8823
rect 49157 8789 49191 8823
rect 53205 8789 53239 8823
rect 57805 8789 57839 8823
rect 2329 8585 2363 8619
rect 4261 8585 4295 8619
rect 7665 8585 7699 8619
rect 10609 8585 10643 8619
rect 14381 8585 14415 8619
rect 15209 8585 15243 8619
rect 17325 8585 17359 8619
rect 17693 8585 17727 8619
rect 20913 8585 20947 8619
rect 21373 8585 21407 8619
rect 24869 8585 24903 8619
rect 25605 8585 25639 8619
rect 26617 8585 26651 8619
rect 27629 8585 27663 8619
rect 27905 8585 27939 8619
rect 47593 8585 47627 8619
rect 51089 8585 51123 8619
rect 51733 8585 51767 8619
rect 54953 8585 54987 8619
rect 57897 8585 57931 8619
rect 3893 8517 3927 8551
rect 7021 8517 7055 8551
rect 10241 8517 10275 8551
rect 13921 8517 13955 8551
rect 14841 8517 14875 8551
rect 34161 8517 34195 8551
rect 35817 8517 35851 8551
rect 38117 8517 38151 8551
rect 38577 8517 38611 8551
rect 45100 8517 45134 8551
rect 47225 8517 47259 8551
rect 48728 8517 48762 8551
rect 53840 8517 53874 8551
rect 55413 8517 55447 8551
rect 3065 8449 3099 8483
rect 3525 8449 3559 8483
rect 3801 8449 3835 8483
rect 6561 8449 6595 8483
rect 6653 8449 6687 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 8401 8449 8435 8483
rect 8668 8449 8702 8483
rect 10333 8449 10367 8483
rect 10977 8449 11011 8483
rect 11621 8449 11655 8483
rect 11888 8449 11922 8483
rect 13277 8449 13311 8483
rect 16681 8449 16715 8483
rect 25513 8449 25547 8483
rect 26157 8449 26191 8483
rect 26985 8449 27019 8483
rect 28365 8449 28399 8483
rect 32781 8449 32815 8483
rect 34345 8449 34379 8483
rect 34529 8449 34563 8483
rect 35725 8449 35759 8483
rect 36277 8449 36311 8483
rect 40417 8449 40451 8483
rect 44833 8449 44867 8483
rect 46397 8449 46431 8483
rect 51825 8449 51859 8483
rect 53573 8449 53607 8483
rect 56195 8449 56229 8483
rect 57253 8449 57287 8483
rect 3157 8381 3191 8415
rect 7113 8381 7147 8415
rect 8309 8381 8343 8415
rect 11069 8381 11103 8415
rect 11161 8381 11195 8415
rect 15485 8381 15519 8415
rect 15761 8381 15795 8415
rect 22661 8381 22695 8415
rect 23397 8381 23431 8415
rect 29377 8381 29411 8415
rect 30665 8381 30699 8415
rect 31401 8381 31435 8415
rect 33517 8381 33551 8415
rect 35909 8381 35943 8415
rect 37841 8381 37875 8415
rect 38025 8381 38059 8415
rect 39129 8381 39163 8415
rect 39865 8381 39899 8415
rect 43085 8381 43119 8415
rect 44741 8381 44775 8415
rect 48973 8381 49007 8415
rect 50445 8381 50479 8415
rect 53389 8381 53423 8415
rect 56057 8381 56091 8415
rect 56333 8381 56367 8415
rect 57069 8381 57103 8415
rect 58449 8381 58483 8415
rect 9781 8313 9815 8347
rect 13001 8313 13035 8347
rect 22109 8313 22143 8347
rect 24685 8313 24719 8347
rect 29929 8313 29963 8347
rect 31769 8313 31803 8347
rect 33977 8313 34011 8347
rect 35173 8313 35207 8347
rect 35357 8313 35391 8347
rect 36829 8313 36863 8347
rect 38485 8313 38519 8347
rect 41061 8313 41095 8347
rect 44097 8313 44131 8347
rect 55321 8313 55355 8347
rect 56609 8313 56643 8347
rect 7481 8245 7515 8279
rect 16405 8245 16439 8279
rect 22845 8245 22879 8279
rect 28181 8245 28215 8279
rect 28825 8245 28859 8279
rect 30113 8245 30147 8279
rect 30849 8245 30883 8279
rect 32689 8245 32723 8279
rect 37473 8245 37507 8279
rect 39313 8245 39347 8279
rect 42441 8245 42475 8279
rect 43453 8245 43487 8279
rect 46213 8245 46247 8279
rect 49893 8245 49927 8279
rect 52377 8245 52411 8279
rect 52837 8245 52871 8279
rect 3433 8041 3467 8075
rect 7573 8041 7607 8075
rect 8953 8041 8987 8075
rect 15485 8041 15519 8075
rect 19901 8041 19935 8075
rect 21005 8041 21039 8075
rect 21833 8041 21867 8075
rect 22753 8041 22787 8075
rect 24685 8041 24719 8075
rect 25237 8041 25271 8075
rect 28825 8041 28859 8075
rect 29837 8041 29871 8075
rect 30021 8041 30055 8075
rect 36185 8041 36219 8075
rect 36277 8041 36311 8075
rect 37749 8041 37783 8075
rect 44649 8041 44683 8075
rect 45017 8041 45051 8075
rect 49893 8041 49927 8075
rect 50169 8041 50203 8075
rect 51733 8041 51767 8075
rect 57805 8041 57839 8075
rect 3801 7973 3835 8007
rect 24869 7973 24903 8007
rect 27169 7973 27203 8007
rect 43361 7973 43395 8007
rect 47317 7973 47351 8007
rect 49065 7973 49099 8007
rect 57713 7973 57747 8007
rect 6837 7905 6871 7939
rect 8585 7905 8619 7939
rect 10333 7905 10367 7939
rect 11069 7905 11103 7939
rect 12127 7905 12161 7939
rect 12541 7905 12575 7939
rect 13829 7905 13863 7939
rect 16037 7905 16071 7939
rect 16129 7905 16163 7939
rect 17601 7905 17635 7939
rect 17877 7905 17911 7939
rect 19257 7905 19291 7939
rect 22109 7905 22143 7939
rect 25881 7905 25915 7939
rect 26157 7905 26191 7939
rect 27997 7905 28031 7939
rect 28181 7905 28215 7939
rect 28365 7905 28399 7939
rect 30573 7905 30607 7939
rect 31217 7905 31251 7939
rect 32321 7905 32355 7939
rect 33425 7905 33459 7939
rect 44005 7905 44039 7939
rect 45569 7905 45603 7939
rect 47777 7905 47811 7939
rect 48605 7905 48639 7939
rect 50721 7905 50755 7939
rect 52285 7905 52319 7939
rect 52653 7905 52687 7939
rect 53757 7905 53791 7939
rect 58357 7905 58391 7939
rect 3524 7837 3558 7871
rect 3617 7837 3651 7871
rect 4076 7837 4110 7871
rect 4169 7837 4203 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 6377 7837 6411 7871
rect 7205 7837 7239 7871
rect 10885 7837 10919 7871
rect 11989 7837 12023 7871
rect 12265 7837 12299 7871
rect 13001 7837 13035 7871
rect 13185 7837 13219 7871
rect 14105 7837 14139 7871
rect 18153 7837 18187 7871
rect 20729 7837 20763 7871
rect 22385 7837 22419 7871
rect 23857 7837 23891 7871
rect 25605 7837 25639 7871
rect 30849 7837 30883 7871
rect 31953 7837 31987 7871
rect 33057 7837 33091 7871
rect 34345 7837 34379 7871
rect 34805 7837 34839 7871
rect 37657 7837 37691 7871
rect 39129 7837 39163 7871
rect 41061 7837 41095 7871
rect 41245 7837 41279 7871
rect 41981 7837 42015 7871
rect 45385 7837 45419 7871
rect 46765 7837 46799 7871
rect 46903 7837 46937 7871
rect 47041 7837 47075 7871
rect 47961 7837 47995 7871
rect 48421 7837 48455 7871
rect 50997 7837 51031 7871
rect 52837 7837 52871 7871
rect 55873 7837 55907 7871
rect 56333 7837 56367 7871
rect 56600 7837 56634 7871
rect 58173 7837 58207 7871
rect 7849 7769 7883 7803
rect 10066 7769 10100 7803
rect 14372 7769 14406 7803
rect 15945 7769 15979 7803
rect 16681 7769 16715 7803
rect 16773 7769 16807 7803
rect 20913 7769 20947 7803
rect 23121 7769 23155 7803
rect 25053 7769 25087 7803
rect 26433 7769 26467 7803
rect 27353 7769 27387 7803
rect 28457 7769 28491 7803
rect 30389 7769 30423 7803
rect 35072 7769 35106 7803
rect 37412 7769 37446 7803
rect 38884 7769 38918 7803
rect 42248 7769 42282 7803
rect 44741 7769 44775 7803
rect 48513 7769 48547 7803
rect 50537 7769 50571 7803
rect 51641 7769 51675 7803
rect 54024 7769 54058 7803
rect 55321 7769 55355 7803
rect 4537 7701 4571 7735
rect 7573 7701 7607 7735
rect 7757 7701 7791 7735
rect 10517 7701 10551 7735
rect 10977 7701 11011 7735
rect 11345 7701 11379 7735
rect 13277 7701 13311 7735
rect 15577 7701 15611 7735
rect 18061 7701 18095 7735
rect 18521 7701 18555 7735
rect 20085 7701 20119 7735
rect 22293 7701 22327 7735
rect 23305 7701 23339 7735
rect 25697 7701 25731 7735
rect 26341 7701 26375 7735
rect 26801 7701 26835 7735
rect 30481 7701 30515 7735
rect 39405 7701 39439 7735
rect 40509 7701 40543 7735
rect 41889 7701 41923 7735
rect 43453 7701 43487 7735
rect 44465 7701 44499 7735
rect 45477 7701 45511 7735
rect 46121 7701 46155 7735
rect 48053 7701 48087 7735
rect 50629 7701 50663 7735
rect 52745 7701 52779 7735
rect 53205 7701 53239 7735
rect 55137 7701 55171 7735
rect 58265 7701 58299 7735
rect 3709 7497 3743 7531
rect 6009 7497 6043 7531
rect 7941 7497 7975 7531
rect 9045 7497 9079 7531
rect 9965 7497 9999 7531
rect 11805 7497 11839 7531
rect 12357 7497 12391 7531
rect 14197 7497 14231 7531
rect 15025 7497 15059 7531
rect 16313 7497 16347 7531
rect 18889 7497 18923 7531
rect 20177 7497 20211 7531
rect 23213 7497 23247 7531
rect 24961 7497 24995 7531
rect 31217 7497 31251 7531
rect 36369 7497 36403 7531
rect 36461 7497 36495 7531
rect 40969 7497 41003 7531
rect 41061 7497 41095 7531
rect 41521 7497 41555 7531
rect 42717 7497 42751 7531
rect 42809 7497 42843 7531
rect 43177 7497 43211 7531
rect 45661 7497 45695 7531
rect 48329 7497 48363 7531
rect 50629 7497 50663 7531
rect 52193 7497 52227 7531
rect 52745 7497 52779 7531
rect 54769 7497 54803 7531
rect 55781 7497 55815 7531
rect 56701 7497 56735 7531
rect 56793 7497 56827 7531
rect 57713 7497 57747 7531
rect 58541 7497 58575 7531
rect 5273 7429 5307 7463
rect 7205 7429 7239 7463
rect 12817 7429 12851 7463
rect 20269 7429 20303 7463
rect 30104 7429 30138 7463
rect 38025 7429 38059 7463
rect 39856 7429 39890 7463
rect 42257 7429 42291 7463
rect 43729 7429 43763 7463
rect 46029 7429 46063 7463
rect 47133 7429 47167 7463
rect 49516 7429 49550 7463
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 7573 7361 7607 7395
rect 7757 7361 7791 7395
rect 8953 7361 8987 7395
rect 9229 7361 9263 7395
rect 9505 7361 9539 7395
rect 11069 7361 11103 7395
rect 15669 7361 15703 7395
rect 16405 7361 16439 7395
rect 18081 7361 18115 7395
rect 21833 7361 21867 7395
rect 22089 7361 22123 7395
rect 23673 7361 23707 7395
rect 25053 7361 25087 7395
rect 27169 7361 27203 7395
rect 28742 7361 28776 7395
rect 29653 7361 29687 7395
rect 32137 7361 32171 7395
rect 32404 7361 32438 7395
rect 33609 7361 33643 7395
rect 34897 7361 34931 7395
rect 37565 7361 37599 7395
rect 39589 7361 39623 7395
rect 41429 7361 41463 7395
rect 43637 7361 43671 7395
rect 44189 7361 44223 7395
rect 44445 7361 44479 7395
rect 46121 7361 46155 7395
rect 47961 7361 47995 7395
rect 53869 7361 53903 7395
rect 54125 7361 54159 7395
rect 54677 7361 54711 7395
rect 55137 7361 55171 7395
rect 57897 7361 57931 7395
rect 5733 7293 5767 7327
rect 5825 7293 5859 7327
rect 6837 7293 6871 7327
rect 8217 7293 8251 7327
rect 10425 7293 10459 7327
rect 12081 7293 12115 7327
rect 12265 7293 12299 7327
rect 13369 7293 13403 7327
rect 13553 7293 13587 7327
rect 14933 7293 14967 7327
rect 18337 7293 18371 7327
rect 19717 7293 19751 7327
rect 20361 7293 20395 7327
rect 21097 7293 21131 7327
rect 21649 7293 21683 7327
rect 23765 7293 23799 7327
rect 23949 7293 23983 7327
rect 24409 7293 24443 7327
rect 29009 7293 29043 7327
rect 29837 7293 29871 7327
rect 31861 7293 31895 7327
rect 33977 7293 34011 7327
rect 35081 7293 35115 7327
rect 36185 7293 36219 7327
rect 37749 7293 37783 7327
rect 37933 7293 37967 7327
rect 41705 7293 41739 7327
rect 42533 7293 42567 7327
rect 43913 7293 43947 7327
rect 46305 7293 46339 7327
rect 46489 7293 46523 7327
rect 49249 7293 49283 7327
rect 51457 7293 51491 7327
rect 51917 7293 51951 7327
rect 52101 7293 52135 7327
rect 54861 7293 54895 7327
rect 56241 7293 56275 7327
rect 56977 7293 57011 7327
rect 5273 7225 5307 7259
rect 9413 7225 9447 7259
rect 12725 7225 12759 7259
rect 19809 7225 19843 7259
rect 27629 7225 27663 7259
rect 36829 7225 36863 7259
rect 38393 7225 38427 7259
rect 52561 7225 52595 7259
rect 7481 7157 7515 7191
rect 10517 7157 10551 7191
rect 14289 7157 14323 7191
rect 16957 7157 16991 7191
rect 19073 7157 19107 7191
rect 20821 7157 20855 7191
rect 23305 7157 23339 7191
rect 26341 7157 26375 7191
rect 29101 7157 29135 7191
rect 31309 7157 31343 7191
rect 33517 7157 33551 7191
rect 38669 7157 38703 7191
rect 39313 7157 39347 7191
rect 43269 7157 43303 7191
rect 45569 7157 45603 7191
rect 50905 7157 50939 7191
rect 54309 7157 54343 7191
rect 56333 7157 56367 7191
rect 4905 6953 4939 6987
rect 5181 6953 5215 6987
rect 6285 6953 6319 6987
rect 9689 6953 9723 6987
rect 10885 6953 10919 6987
rect 15393 6953 15427 6987
rect 18337 6953 18371 6987
rect 20637 6953 20671 6987
rect 22937 6953 22971 6987
rect 24501 6953 24535 6987
rect 35633 6953 35667 6987
rect 38117 6953 38151 6987
rect 41061 6953 41095 6987
rect 46213 6953 46247 6987
rect 46489 6953 46523 6987
rect 50353 6953 50387 6987
rect 54217 6953 54251 6987
rect 56793 6953 56827 6987
rect 36921 6885 36955 6919
rect 38393 6885 38427 6919
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 6009 6817 6043 6851
rect 6126 6817 6160 6851
rect 7573 6817 7607 6851
rect 10701 6817 10735 6851
rect 11529 6817 11563 6851
rect 14565 6817 14599 6851
rect 14657 6817 14691 6851
rect 15577 6817 15611 6851
rect 16221 6817 16255 6851
rect 16614 6817 16648 6851
rect 16773 6817 16807 6851
rect 17601 6817 17635 6851
rect 19257 6817 19291 6851
rect 21005 6817 21039 6851
rect 22201 6817 22235 6851
rect 22661 6817 22695 6851
rect 22845 6817 22879 6851
rect 23397 6817 23431 6851
rect 23489 6817 23523 6851
rect 26249 6817 26283 6851
rect 26433 6817 26467 6851
rect 26893 6817 26927 6851
rect 27286 6817 27320 6851
rect 27445 6817 27479 6851
rect 28273 6817 28307 6851
rect 32137 6817 32171 6851
rect 32689 6817 32723 6851
rect 34713 6817 34747 6851
rect 35817 6817 35851 6851
rect 36277 6817 36311 6851
rect 36461 6817 36495 6851
rect 37314 6817 37348 6851
rect 37473 6817 37507 6851
rect 38761 6817 38795 6851
rect 39589 6817 39623 6851
rect 40601 6817 40635 6851
rect 42027 6817 42061 6851
rect 42441 6817 42475 6851
rect 42901 6817 42935 6851
rect 43729 6817 43763 6851
rect 45569 6817 45603 6851
rect 47777 6817 47811 6851
rect 49893 6817 49927 6851
rect 51365 6817 51399 6851
rect 51503 6817 51537 6851
rect 51917 6817 51951 6851
rect 52377 6817 52411 6851
rect 53941 6817 53975 6851
rect 54769 6817 54803 6851
rect 56241 6817 56275 6851
rect 57437 6817 57471 6851
rect 58357 6817 58391 6851
rect 2697 6749 2731 6783
rect 2881 6749 2915 6783
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 4261 6749 4295 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7941 6749 7975 6783
rect 8769 6749 8803 6783
rect 10149 6749 10183 6783
rect 11253 6749 11287 6783
rect 11713 6749 11747 6783
rect 13369 6749 13403 6783
rect 14473 6749 14507 6783
rect 15761 6749 15795 6783
rect 16497 6749 16531 6783
rect 17417 6749 17451 6783
rect 18889 6749 18923 6783
rect 19513 6749 19547 6783
rect 21649 6749 21683 6783
rect 21787 6749 21821 6783
rect 21925 6749 21959 6783
rect 25625 6749 25659 6783
rect 25881 6749 25915 6783
rect 27169 6749 27203 6783
rect 28549 6749 28583 6783
rect 31145 6749 31179 6783
rect 31401 6749 31435 6783
rect 32296 6749 32330 6783
rect 32413 6749 32447 6783
rect 33149 6749 33183 6783
rect 33333 6749 33367 6783
rect 33517 6749 33551 6783
rect 35265 6749 35299 6783
rect 37197 6749 37231 6783
rect 41889 6749 41923 6783
rect 42165 6749 42199 6783
rect 43085 6749 43119 6783
rect 47869 6749 47903 6783
rect 48421 6749 48455 6783
rect 49157 6749 49191 6783
rect 51641 6749 51675 6783
rect 52561 6749 52595 6783
rect 53205 6749 53239 6783
rect 57345 6749 57379 6783
rect 57953 6749 57987 6783
rect 3341 6681 3375 6715
rect 3801 6681 3835 6715
rect 3985 6681 4019 6715
rect 4169 6681 4203 6715
rect 5181 6681 5215 6715
rect 9045 6681 9079 6715
rect 9229 6681 9263 6715
rect 11345 6681 11379 6715
rect 12541 6681 12575 6715
rect 17877 6681 17911 6715
rect 34253 6681 34287 6715
rect 36001 6681 36035 6715
rect 38945 6681 38979 6715
rect 40509 6681 40543 6715
rect 45477 6681 45511 6715
rect 46397 6681 46431 6715
rect 56885 6681 56919 6715
rect 57621 6681 57655 6715
rect 58081 6681 58115 6715
rect 58173 6681 58207 6715
rect 58357 6681 58391 6715
rect 2789 6613 2823 6647
rect 4997 6613 5031 6647
rect 5917 6613 5951 6647
rect 10057 6613 10091 6647
rect 13001 6613 13035 6647
rect 13921 6613 13955 6647
rect 14105 6613 14139 6647
rect 17785 6613 17819 6647
rect 18245 6613 18279 6647
rect 23305 6613 23339 6647
rect 24225 6613 24259 6647
rect 28089 6613 28123 6647
rect 28457 6613 28491 6647
rect 28917 6613 28951 6647
rect 30021 6613 30055 6647
rect 31493 6613 31527 6647
rect 40049 6613 40083 6647
rect 40417 6613 40451 6647
rect 41245 6613 41279 6647
rect 43177 6613 43211 6647
rect 47133 6613 47167 6647
rect 48605 6613 48639 6647
rect 50721 6613 50755 6647
rect 52653 6613 52687 6647
rect 53389 6613 53423 6647
rect 55597 6613 55631 6647
rect 56609 6613 56643 6647
rect 3617 6409 3651 6443
rect 6745 6409 6779 6443
rect 8677 6409 8711 6443
rect 11253 6409 11287 6443
rect 12081 6409 12115 6443
rect 14105 6409 14139 6443
rect 14473 6409 14507 6443
rect 18153 6409 18187 6443
rect 21005 6409 21039 6443
rect 21649 6409 21683 6443
rect 23213 6409 23247 6443
rect 26985 6409 27019 6443
rect 27997 6409 28031 6443
rect 28733 6409 28767 6443
rect 31033 6409 31067 6443
rect 31493 6409 31527 6443
rect 35081 6409 35115 6443
rect 36829 6409 36863 6443
rect 37749 6409 37783 6443
rect 41521 6409 41555 6443
rect 47409 6409 47443 6443
rect 47593 6409 47627 6443
rect 51917 6409 51951 6443
rect 56609 6409 56643 6443
rect 57897 6409 57931 6443
rect 14565 6341 14599 6375
rect 17141 6341 17175 6375
rect 17325 6341 17359 6375
rect 22100 6341 22134 6375
rect 25044 6341 25078 6375
rect 50804 6341 50838 6375
rect 52285 6341 52319 6375
rect 56517 6341 56551 6375
rect 1593 6273 1627 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3709 6273 3743 6307
rect 4261 6273 4295 6307
rect 5089 6273 5123 6307
rect 6377 6273 6411 6307
rect 7564 6273 7598 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 9965 6273 9999 6307
rect 12173 6273 12207 6307
rect 14933 6273 14967 6307
rect 15200 6273 15234 6307
rect 17509 6273 17543 6307
rect 18797 6273 18831 6307
rect 19073 6273 19107 6307
rect 19340 6273 19374 6307
rect 20913 6273 20947 6307
rect 21833 6273 21867 6307
rect 23857 6273 23891 6307
rect 24593 6273 24627 6307
rect 26525 6273 26559 6307
rect 28825 6273 28859 6307
rect 31125 6273 31159 6307
rect 32413 6273 32447 6307
rect 32669 6273 32703 6307
rect 34529 6273 34563 6307
rect 36553 6273 36587 6307
rect 37657 6273 37691 6307
rect 38853 6273 38887 6307
rect 39405 6273 39439 6307
rect 39672 6273 39706 6307
rect 41705 6273 41739 6307
rect 42809 6273 42843 6307
rect 46029 6273 46063 6307
rect 46296 6273 46330 6307
rect 47961 6273 47995 6307
rect 48053 6273 48087 6307
rect 49065 6273 49099 6307
rect 49332 6273 49366 6307
rect 50537 6273 50571 6307
rect 1869 6205 1903 6239
rect 4445 6205 4479 6239
rect 5825 6205 5859 6239
rect 7297 6205 7331 6239
rect 10609 6205 10643 6239
rect 14749 6205 14783 6239
rect 17049 6205 17083 6239
rect 21189 6205 21223 6239
rect 24409 6205 24443 6239
rect 24777 6205 24811 6239
rect 27629 6205 27663 6239
rect 30941 6205 30975 6239
rect 31769 6205 31803 6239
rect 37841 6205 37875 6239
rect 40877 6205 40911 6239
rect 42165 6205 42199 6239
rect 42533 6205 42567 6239
rect 42717 6205 42751 6239
rect 43821 6205 43855 6239
rect 48145 6205 48179 6239
rect 55505 6205 55539 6239
rect 56333 6205 56367 6239
rect 57621 6205 57655 6239
rect 58541 6205 58575 6239
rect 5273 6137 5307 6171
rect 5641 6137 5675 6171
rect 9689 6137 9723 6171
rect 20453 6137 20487 6171
rect 26157 6137 26191 6171
rect 33793 6137 33827 6171
rect 40785 6137 40819 6171
rect 41889 6137 41923 6171
rect 43177 6137 43211 6171
rect 56977 6137 57011 6171
rect 3157 6069 3191 6103
rect 4537 6069 4571 6103
rect 5733 6069 5767 6103
rect 6101 6069 6135 6103
rect 6745 6069 6779 6103
rect 6929 6069 6963 6103
rect 9137 6069 9171 6103
rect 13645 6069 13679 6103
rect 16313 6069 16347 6103
rect 18245 6069 18279 6103
rect 20545 6069 20579 6103
rect 23305 6069 23339 6103
rect 33885 6069 33919 6103
rect 37289 6069 37323 6103
rect 38301 6069 38335 6103
rect 39313 6069 39347 6103
rect 43269 6069 43303 6103
rect 50445 6069 50479 6103
rect 54125 6069 54159 6103
rect 54953 6069 54987 6103
rect 55413 6069 55447 6103
rect 56149 6069 56183 6103
rect 57069 6069 57103 6103
rect 2145 5865 2179 5899
rect 2973 5865 3007 5899
rect 6469 5865 6503 5899
rect 8401 5865 8435 5899
rect 12725 5865 12759 5899
rect 15577 5865 15611 5899
rect 16497 5865 16531 5899
rect 17601 5865 17635 5899
rect 19993 5865 20027 5899
rect 21373 5865 21407 5899
rect 31217 5865 31251 5899
rect 32413 5865 32447 5899
rect 33241 5865 33275 5899
rect 38117 5865 38151 5899
rect 39589 5865 39623 5899
rect 39865 5865 39899 5899
rect 40877 5865 40911 5899
rect 43361 5865 43395 5899
rect 47409 5865 47443 5899
rect 49341 5865 49375 5899
rect 50997 5865 51031 5899
rect 55137 5865 55171 5899
rect 58173 5865 58207 5899
rect 26065 5797 26099 5831
rect 34989 5797 35023 5831
rect 36645 5797 36679 5831
rect 41245 5797 41279 5831
rect 43269 5797 43303 5831
rect 50169 5797 50203 5831
rect 58357 5797 58391 5831
rect 2053 5729 2087 5763
rect 3525 5729 3559 5763
rect 9873 5729 9907 5763
rect 14197 5729 14231 5763
rect 16129 5729 16163 5763
rect 16313 5729 16347 5763
rect 17049 5729 17083 5763
rect 20545 5729 20579 5763
rect 20729 5729 20763 5763
rect 23213 5729 23247 5763
rect 24685 5729 24719 5763
rect 26709 5729 26743 5763
rect 26985 5729 27019 5763
rect 30113 5729 30147 5763
rect 30573 5729 30607 5763
rect 32045 5729 32079 5763
rect 32597 5729 32631 5763
rect 33793 5729 33827 5763
rect 33885 5729 33919 5763
rect 35265 5729 35299 5763
rect 37381 5729 37415 5763
rect 43913 5729 43947 5763
rect 46857 5729 46891 5763
rect 49985 5729 50019 5763
rect 50629 5729 50663 5763
rect 50721 5729 50755 5763
rect 51457 5729 51491 5763
rect 51641 5729 51675 5763
rect 1777 5661 1811 5695
rect 1961 5661 1995 5695
rect 2697 5661 2731 5695
rect 4077 5661 4111 5695
rect 4344 5661 4378 5695
rect 7113 5661 7147 5695
rect 8033 5661 8067 5695
rect 9229 5661 9263 5695
rect 11345 5661 11379 5695
rect 13553 5661 13587 5695
rect 14453 5661 14487 5695
rect 16037 5661 16071 5695
rect 18245 5661 18279 5695
rect 22845 5661 22879 5695
rect 26525 5661 26559 5695
rect 27629 5661 27663 5695
rect 28825 5661 28859 5695
rect 32873 5661 32907 5695
rect 33701 5661 33735 5695
rect 37473 5661 37507 5695
rect 38761 5661 38795 5695
rect 40417 5661 40451 5695
rect 41889 5661 41923 5695
rect 45201 5661 45235 5695
rect 46121 5661 46155 5695
rect 46489 5661 46523 5695
rect 50537 5661 50571 5695
rect 53205 5661 53239 5695
rect 55321 5661 55355 5695
rect 56793 5661 56827 5695
rect 57060 5661 57094 5695
rect 58541 5661 58575 5695
rect 1593 5593 1627 5627
rect 7573 5593 7607 5627
rect 8769 5593 8803 5627
rect 10140 5593 10174 5627
rect 11612 5593 11646 5627
rect 12909 5593 12943 5627
rect 24952 5593 24986 5627
rect 26617 5593 26651 5627
rect 32781 5593 32815 5627
rect 35532 5593 35566 5627
rect 36737 5593 36771 5627
rect 42156 5593 42190 5627
rect 44373 5593 44407 5627
rect 55588 5593 55622 5627
rect 5457 5525 5491 5559
rect 9781 5525 9815 5559
rect 11253 5525 11287 5559
rect 13921 5525 13955 5559
rect 15669 5525 15703 5559
rect 17693 5525 17727 5559
rect 19441 5525 19475 5559
rect 22293 5525 22327 5559
rect 26157 5525 26191 5559
rect 28273 5525 28307 5559
rect 29561 5525 29595 5559
rect 33333 5525 33367 5559
rect 34437 5525 34471 5559
rect 38209 5525 38243 5559
rect 39129 5525 39163 5559
rect 41705 5525 41739 5559
rect 44649 5525 44683 5559
rect 45569 5525 45603 5559
rect 51365 5525 51399 5559
rect 52193 5525 52227 5559
rect 52653 5525 52687 5559
rect 54769 5525 54803 5559
rect 56701 5525 56735 5559
rect 3433 5321 3467 5355
rect 3596 5321 3630 5355
rect 3893 5321 3927 5355
rect 12173 5321 12207 5355
rect 22385 5321 22419 5355
rect 25605 5321 25639 5355
rect 26617 5321 26651 5355
rect 32505 5321 32539 5355
rect 33241 5321 33275 5355
rect 33977 5321 34011 5355
rect 35173 5321 35207 5355
rect 36185 5321 36219 5355
rect 42809 5321 42843 5355
rect 45661 5321 45695 5355
rect 49985 5321 50019 5355
rect 51181 5321 51215 5355
rect 51549 5321 51583 5355
rect 51917 5321 51951 5355
rect 52745 5321 52779 5355
rect 53113 5321 53147 5355
rect 55413 5321 55447 5355
rect 55781 5321 55815 5355
rect 57713 5321 57747 5355
rect 2973 5253 3007 5287
rect 3801 5253 3835 5287
rect 7665 5253 7699 5287
rect 9321 5253 9355 5287
rect 14013 5253 14047 5287
rect 15485 5253 15519 5287
rect 17684 5253 17718 5287
rect 22201 5253 22235 5287
rect 22753 5253 22787 5287
rect 28172 5253 28206 5287
rect 31953 5253 31987 5287
rect 36737 5253 36771 5287
rect 39313 5253 39347 5287
rect 45324 5253 45358 5287
rect 46029 5253 46063 5287
rect 47317 5253 47351 5287
rect 4537 5185 4571 5219
rect 7849 5185 7883 5219
rect 8116 5185 8150 5219
rect 10885 5185 10919 5219
rect 11529 5185 11563 5219
rect 12449 5185 12483 5219
rect 15393 5185 15427 5219
rect 16037 5185 16071 5219
rect 16497 5185 16531 5219
rect 20453 5185 20487 5219
rect 22845 5185 22879 5219
rect 26249 5185 26283 5219
rect 33149 5185 33183 5219
rect 33793 5185 33827 5219
rect 34529 5185 34563 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 37013 5185 37047 5219
rect 37381 5185 37415 5219
rect 37648 5185 37682 5219
rect 44097 5185 44131 5219
rect 45569 5185 45603 5219
rect 46857 5185 46891 5219
rect 47041 5185 47075 5219
rect 47593 5185 47627 5219
rect 50537 5185 50571 5219
rect 52193 5185 52227 5219
rect 53205 5185 53239 5219
rect 53849 5185 53883 5219
rect 56333 5185 56367 5219
rect 56589 5185 56623 5219
rect 58449 5185 58483 5219
rect 4997 5117 5031 5151
rect 17417 5117 17451 5151
rect 19441 5117 19475 5151
rect 22937 5117 22971 5151
rect 27905 5117 27939 5151
rect 29561 5117 29595 5151
rect 35541 5117 35575 5151
rect 41061 5117 41095 5151
rect 42257 5117 42291 5151
rect 42901 5117 42935 5151
rect 43085 5117 43119 5151
rect 43545 5117 43579 5151
rect 46121 5117 46155 5151
rect 46305 5117 46339 5151
rect 46765 5117 46799 5151
rect 48145 5117 48179 5151
rect 52469 5117 52503 5151
rect 53297 5117 53331 5151
rect 55229 5117 55263 5151
rect 55873 5117 55907 5151
rect 55965 5117 55999 5151
rect 3341 5049 3375 5083
rect 5365 5049 5399 5083
rect 9229 5049 9263 5083
rect 17233 5049 17267 5083
rect 18797 5049 18831 5083
rect 29285 5049 29319 5083
rect 42441 5049 42475 5083
rect 44189 5049 44223 5083
rect 52009 5049 52043 5083
rect 54217 5049 54251 5083
rect 2789 4981 2823 5015
rect 2973 4981 3007 5015
rect 3617 4981 3651 5015
rect 7021 4981 7055 5015
rect 7389 4981 7423 5015
rect 14841 4981 14875 5015
rect 18889 4981 18923 5015
rect 19901 4981 19935 5015
rect 21005 4981 21039 5015
rect 21373 4981 21407 5015
rect 23397 4981 23431 5015
rect 23857 4981 23891 5015
rect 30205 4981 30239 5015
rect 32413 4981 32447 5015
rect 34897 4981 34931 5015
rect 38761 4981 38795 5015
rect 39037 4981 39071 5015
rect 41429 4981 41463 5015
rect 41613 4981 41647 5015
rect 47041 4981 47075 5015
rect 49709 4981 49743 5015
rect 50445 4981 50479 5015
rect 54585 4981 54619 5015
rect 54861 4981 54895 5015
rect 57897 4981 57931 5015
rect 3801 4777 3835 4811
rect 5089 4777 5123 4811
rect 9137 4777 9171 4811
rect 11161 4777 11195 4811
rect 11621 4777 11655 4811
rect 13093 4777 13127 4811
rect 15117 4777 15151 4811
rect 17693 4777 17727 4811
rect 19349 4777 19383 4811
rect 21557 4777 21591 4811
rect 24869 4777 24903 4811
rect 25145 4777 25179 4811
rect 28089 4777 28123 4811
rect 28273 4777 28307 4811
rect 34805 4777 34839 4811
rect 37289 4777 37323 4811
rect 38485 4777 38519 4811
rect 40049 4777 40083 4811
rect 54677 4777 54711 4811
rect 56057 4777 56091 4811
rect 4537 4709 4571 4743
rect 10057 4709 10091 4743
rect 16773 4709 16807 4743
rect 32689 4709 32723 4743
rect 42257 4709 42291 4743
rect 46029 4709 46063 4743
rect 3341 4641 3375 4675
rect 4445 4641 4479 4675
rect 7297 4641 7331 4675
rect 9781 4641 9815 4675
rect 10701 4641 10735 4675
rect 18153 4641 18187 4675
rect 18337 4641 18371 4675
rect 26801 4641 26835 4675
rect 27721 4641 27755 4675
rect 28825 4641 28859 4675
rect 32137 4641 32171 4675
rect 34529 4641 34563 4675
rect 35449 4641 35483 4675
rect 35541 4641 35575 4675
rect 37841 4641 37875 4675
rect 38761 4641 38795 4675
rect 40325 4641 40359 4675
rect 40693 4641 40727 4675
rect 40877 4641 40911 4675
rect 42349 4641 42383 4675
rect 46581 4641 46615 4675
rect 49249 4641 49283 4675
rect 56333 4641 56367 4675
rect 56885 4641 56919 4675
rect 4537 4573 4571 4607
rect 4809 4573 4843 4607
rect 4913 4573 4947 4607
rect 5641 4573 5675 4607
rect 5825 4573 5859 4607
rect 6009 4573 6043 4607
rect 6101 4573 6135 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 8677 4573 8711 4607
rect 10425 4573 10459 4607
rect 14657 4573 14691 4607
rect 16037 4573 16071 4607
rect 17601 4573 17635 4607
rect 18521 4573 18555 4607
rect 18705 4573 18739 4607
rect 18981 4573 19015 4607
rect 19533 4573 19567 4607
rect 20269 4573 20303 4607
rect 20637 4573 20671 4607
rect 20729 4573 20763 4607
rect 20913 4573 20947 4607
rect 21281 4573 21315 4607
rect 22017 4573 22051 4607
rect 23857 4573 23891 4607
rect 24409 4573 24443 4607
rect 25329 4573 25363 4607
rect 26341 4573 26375 4607
rect 26525 4573 26559 4607
rect 28641 4573 28675 4607
rect 29745 4573 29779 4607
rect 30389 4573 30423 4607
rect 31861 4573 31895 4607
rect 32781 4573 32815 4607
rect 35914 4573 35948 4607
rect 36093 4573 36127 4607
rect 36829 4573 36863 4607
rect 38117 4573 38151 4607
rect 39589 4573 39623 4607
rect 39865 4573 39899 4607
rect 41144 4573 41178 4607
rect 43085 4573 43119 4607
rect 43269 4573 43303 4607
rect 43361 4573 43395 4607
rect 43545 4573 43579 4607
rect 43821 4573 43855 4607
rect 44741 4573 44775 4607
rect 45201 4573 45235 4607
rect 46305 4573 46339 4607
rect 46848 4573 46882 4607
rect 48237 4573 48271 4607
rect 49525 4573 49559 4607
rect 49709 4573 49743 4607
rect 49893 4573 49927 4607
rect 50169 4573 50203 4607
rect 51917 4573 51951 4607
rect 52193 4573 52227 4607
rect 53757 4573 53791 4607
rect 55045 4573 55079 4607
rect 55781 4573 55815 4607
rect 55873 4573 55907 4607
rect 56057 4573 56091 4607
rect 57161 4573 57195 4607
rect 4721 4505 4755 4539
rect 7665 4505 7699 4539
rect 8033 4505 8067 4539
rect 14105 4505 14139 4539
rect 17141 4505 17175 4539
rect 18061 4505 18095 4539
rect 19809 4505 19843 4539
rect 20821 4505 20855 4539
rect 26157 4505 26191 4539
rect 28733 4505 28767 4539
rect 31493 4505 31527 4539
rect 32321 4505 32355 4539
rect 33609 4505 33643 4539
rect 35541 4505 35575 4539
rect 35725 4505 35759 4539
rect 35817 4505 35851 4539
rect 36369 4505 36403 4539
rect 43177 4505 43211 4539
rect 44097 4505 44131 4539
rect 52460 4505 52494 4539
rect 58357 4505 58391 4539
rect 2145 4437 2179 4471
rect 2789 4437 2823 4471
rect 5549 4437 5583 4471
rect 8125 4437 8159 4471
rect 10517 4437 10551 4471
rect 12173 4437 12207 4471
rect 13553 4437 13587 4471
rect 13921 4437 13955 4471
rect 15485 4437 15519 4471
rect 16405 4437 16439 4471
rect 18613 4437 18647 4471
rect 18797 4437 18831 4471
rect 21097 4437 21131 4471
rect 22385 4437 22419 4471
rect 24133 4437 24167 4471
rect 24593 4437 24627 4471
rect 26433 4437 26467 4471
rect 27445 4437 27479 4471
rect 29377 4437 29411 4471
rect 31125 4437 31159 4471
rect 32229 4437 32263 4471
rect 33885 4437 33919 4471
rect 37565 4437 37599 4471
rect 38025 4437 38059 4471
rect 39313 4437 39347 4471
rect 42993 4437 43027 4471
rect 43453 4437 43487 4471
rect 43637 4437 43671 4471
rect 45569 4437 45603 4471
rect 47961 4437 47995 4471
rect 48697 4437 48731 4471
rect 49801 4437 49835 4471
rect 53573 4437 53607 4471
rect 54309 4437 54343 4471
rect 55597 4437 55631 4471
rect 6377 4233 6411 4267
rect 10977 4233 11011 4267
rect 15025 4233 15059 4267
rect 21005 4233 21039 4267
rect 23397 4233 23431 4267
rect 27997 4233 28031 4267
rect 30205 4233 30239 4267
rect 34253 4233 34287 4267
rect 36277 4233 36311 4267
rect 48605 4233 48639 4267
rect 50169 4233 50203 4267
rect 53573 4233 53607 4267
rect 2688 4165 2722 4199
rect 4629 4165 4663 4199
rect 8493 4165 8527 4199
rect 13553 4165 13587 4199
rect 13829 4165 13863 4199
rect 15669 4165 15703 4199
rect 17877 4165 17911 4199
rect 18153 4165 18187 4199
rect 24593 4165 24627 4199
rect 28549 4165 28583 4199
rect 29929 4165 29963 4199
rect 30113 4165 30147 4199
rect 33272 4165 33306 4199
rect 34796 4165 34830 4199
rect 38301 4165 38335 4199
rect 38485 4165 38519 4199
rect 40049 4165 40083 4199
rect 40141 4165 40175 4199
rect 41245 4165 41279 4199
rect 42257 4165 42291 4199
rect 43729 4165 43763 4199
rect 44373 4165 44407 4199
rect 45385 4165 45419 4199
rect 45477 4165 45511 4199
rect 46949 4165 46983 4199
rect 47133 4165 47167 4199
rect 47225 4165 47259 4199
rect 51089 4165 51123 4199
rect 52929 4165 52963 4199
rect 57069 4165 57103 4199
rect 57345 4165 57379 4199
rect 1409 4097 1443 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 4077 4097 4111 4131
rect 4353 4097 4387 4131
rect 4721 4097 4755 4131
rect 4813 4097 4847 4131
rect 5917 4097 5951 4131
rect 7113 4097 7147 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 7941 4097 7975 4131
rect 8120 4087 8154 4121
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 9321 4097 9355 4131
rect 9505 4097 9539 4131
rect 9689 4097 9723 4131
rect 13456 4097 13490 4131
rect 13645 4097 13679 4131
rect 13927 4097 13961 4131
rect 14105 4097 14139 4131
rect 14197 4097 14231 4131
rect 14933 4097 14967 4131
rect 15117 4097 15151 4131
rect 15296 4087 15330 4121
rect 15393 4097 15427 4131
rect 15485 4097 15519 4131
rect 17601 4097 17635 4131
rect 18337 4097 18371 4131
rect 18429 4097 18463 4131
rect 18526 4097 18560 4131
rect 18705 4097 18739 4131
rect 19717 4097 19751 4131
rect 19901 4097 19935 4131
rect 19993 4097 20027 4131
rect 20090 4097 20124 4131
rect 21189 4097 21223 4131
rect 21373 4097 21407 4131
rect 21465 4097 21499 4131
rect 21649 4097 21683 4131
rect 21925 4097 21959 4131
rect 22192 4097 22226 4131
rect 24317 4097 24351 4131
rect 24925 4097 24959 4131
rect 25053 4097 25087 4131
rect 25145 4097 25179 4131
rect 25329 4097 25363 4131
rect 26801 4097 26835 4131
rect 26985 4097 27019 4131
rect 28181 4097 28215 4131
rect 28360 4097 28394 4131
rect 28457 4097 28491 4131
rect 28733 4097 28767 4131
rect 29709 4087 29743 4121
rect 29837 4097 29871 4131
rect 30389 4097 30423 4131
rect 30665 4097 30699 4131
rect 30757 4097 30791 4131
rect 30941 4097 30975 4131
rect 31217 4097 31251 4131
rect 33517 4097 33551 4131
rect 34529 4097 34563 4131
rect 36369 4097 36403 4131
rect 36645 4097 36679 4131
rect 36829 4097 36863 4131
rect 37289 4097 37323 4131
rect 38081 4097 38115 4131
rect 38209 4097 38243 4131
rect 38577 4097 38611 4131
rect 38761 4097 38795 4131
rect 38853 4097 38887 4131
rect 39773 4097 39807 4131
rect 40325 4097 40359 4131
rect 40417 4097 40451 4131
rect 40545 4097 40579 4131
rect 41429 4097 41463 4131
rect 41853 4097 41887 4131
rect 41981 4097 42015 4131
rect 42073 4097 42107 4131
rect 43269 4097 43303 4131
rect 44097 4097 44131 4131
rect 45288 4087 45322 4121
rect 45661 4097 45695 4131
rect 45753 4097 45787 4131
rect 45937 4097 45971 4131
rect 46029 4097 46063 4131
rect 46581 4097 46615 4131
rect 47337 4103 47371 4137
rect 48053 4097 48087 4131
rect 48237 4097 48271 4131
rect 49433 4097 49467 4131
rect 49893 4097 49927 4131
rect 50905 4097 50939 4131
rect 51181 4097 51215 4131
rect 51309 4097 51343 4131
rect 52285 4097 52319 4131
rect 52377 4097 52411 4131
rect 52561 4097 52595 4131
rect 53205 4097 53239 4131
rect 53389 4097 53423 4131
rect 54125 4097 54159 4131
rect 54309 4097 54343 4131
rect 54493 4097 54527 4131
rect 54769 4097 54803 4131
rect 55229 4097 55263 4131
rect 55413 4097 55447 4131
rect 55597 4097 55631 4131
rect 56333 4097 56367 4131
rect 56517 4097 56551 4131
rect 56609 4097 56643 4131
rect 56721 4119 56755 4153
rect 56972 4097 57006 4131
rect 57161 4097 57195 4131
rect 57437 4097 57471 4131
rect 2421 4029 2455 4063
rect 4997 4029 5031 4063
rect 6929 4029 6963 4063
rect 8401 4029 8435 4063
rect 8585 4029 8619 4063
rect 10241 4029 10275 4063
rect 11529 4029 11563 4063
rect 13277 4029 13311 4063
rect 13737 4029 13771 4063
rect 14841 4029 14875 4063
rect 15577 4029 15611 4063
rect 16313 4029 16347 4063
rect 17233 4029 17267 4063
rect 17785 4029 17819 4063
rect 19257 4029 19291 4063
rect 19809 4029 19843 4063
rect 20361 4029 20395 4063
rect 23949 4029 23983 4063
rect 24409 4029 24443 4063
rect 25237 4029 25271 4063
rect 25973 4029 26007 4063
rect 27445 4029 27479 4063
rect 27813 4029 27847 4063
rect 28641 4029 28675 4063
rect 29377 4029 29411 4063
rect 30481 4029 30515 4063
rect 33609 4029 33643 4063
rect 37933 4029 37967 4063
rect 38393 4029 38427 4063
rect 39497 4029 39531 4063
rect 39865 4029 39899 4063
rect 42165 4029 42199 4063
rect 42441 4029 42475 4063
rect 43085 4029 43119 4063
rect 44189 4029 44223 4063
rect 44465 4029 44499 4063
rect 45017 4029 45051 4063
rect 47225 4029 47259 4063
rect 48973 4029 49007 4063
rect 49617 4029 49651 4063
rect 50813 4029 50847 4063
rect 50997 4029 51031 4063
rect 51641 4029 51675 4063
rect 55045 4029 55079 4063
rect 56241 4029 56275 4063
rect 56425 4029 56459 4063
rect 57253 4029 57287 4063
rect 57897 4029 57931 4063
rect 1593 3961 1627 3995
rect 3801 3961 3835 3995
rect 7205 3961 7239 3995
rect 12633 3961 12667 3995
rect 14105 3961 14139 3995
rect 15761 3961 15795 3995
rect 17417 3961 17451 3995
rect 18153 3961 18187 3995
rect 23305 3961 23339 3995
rect 25421 3961 25455 3995
rect 27169 3961 27203 3995
rect 28825 3961 28859 3995
rect 30113 3961 30147 3995
rect 32137 3961 32171 3995
rect 35909 3961 35943 3995
rect 36553 3961 36587 3995
rect 40141 3961 40175 3995
rect 45661 3961 45695 3995
rect 49249 3961 49283 3995
rect 1869 3893 1903 3927
rect 2145 3893 2179 3927
rect 5365 3893 5399 3927
rect 7573 3893 7607 3927
rect 7757 3893 7791 3927
rect 9229 3893 9263 3927
rect 9505 3893 9539 3927
rect 11253 3893 11287 3927
rect 12173 3893 12207 3927
rect 12449 3893 12483 3927
rect 14381 3893 14415 3927
rect 16681 3893 16715 3927
rect 17601 3893 17635 3927
rect 21373 3893 21407 3927
rect 21649 3893 21683 3927
rect 24133 3893 24167 3927
rect 24409 3893 24443 3927
rect 26433 3893 26467 3927
rect 26617 3893 26651 3927
rect 30665 3893 30699 3927
rect 30757 3893 30791 3927
rect 31677 3893 31711 3927
rect 36829 3893 36863 3927
rect 38761 3893 38795 3927
rect 39589 3893 39623 3927
rect 39957 3893 39991 3927
rect 40877 3893 40911 3927
rect 41613 3893 41647 3927
rect 43453 3893 43487 3927
rect 43913 3893 43947 3927
rect 44189 3893 44223 3927
rect 45937 3893 45971 3927
rect 47777 3893 47811 3927
rect 48237 3893 48271 3927
rect 49617 3893 49651 3927
rect 52377 3893 52411 3927
rect 54309 3893 54343 3927
rect 54585 3893 54619 3927
rect 55413 3893 55447 3927
rect 57621 3893 57655 3927
rect 58541 3893 58575 3927
rect 3157 3689 3191 3723
rect 6193 3689 6227 3723
rect 6285 3689 6319 3723
rect 6653 3689 6687 3723
rect 10517 3689 10551 3723
rect 13921 3689 13955 3723
rect 17601 3689 17635 3723
rect 19073 3689 19107 3723
rect 20913 3689 20947 3723
rect 22477 3689 22511 3723
rect 22753 3689 22787 3723
rect 25881 3689 25915 3723
rect 30941 3689 30975 3723
rect 37657 3689 37691 3723
rect 43361 3689 43395 3723
rect 44833 3689 44867 3723
rect 54585 3689 54619 3723
rect 55045 3689 55079 3723
rect 56885 3689 56919 3723
rect 58541 3689 58575 3723
rect 14197 3621 14231 3655
rect 15025 3621 15059 3655
rect 34529 3621 34563 3655
rect 39313 3621 39347 3655
rect 45017 3621 45051 3655
rect 46949 3621 46983 3655
rect 49249 3621 49283 3655
rect 2973 3553 3007 3587
rect 14565 3553 14599 3587
rect 17693 3553 17727 3587
rect 21097 3553 21131 3587
rect 31493 3553 31527 3587
rect 33149 3553 33183 3587
rect 34805 3553 34839 3587
rect 35449 3553 35483 3587
rect 36277 3553 36311 3587
rect 43453 3553 43487 3587
rect 45293 3553 45327 3587
rect 47777 3553 47811 3587
rect 50169 3553 50203 3587
rect 54493 3553 54527 3587
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 4813 3485 4847 3519
rect 6469 3485 6503 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 8309 3485 8343 3519
rect 8953 3485 8987 3519
rect 10890 3495 10924 3529
rect 12449 3485 12483 3519
rect 12541 3485 12575 3519
rect 14381 3485 14415 3519
rect 14479 3485 14513 3519
rect 14657 3485 14691 3519
rect 14841 3485 14875 3519
rect 15301 3485 15335 3519
rect 15557 3485 15591 3519
rect 17049 3485 17083 3519
rect 20370 3485 20404 3519
rect 20637 3485 20671 3519
rect 20729 3485 20763 3519
rect 22569 3485 22603 3519
rect 22845 3485 22879 3519
rect 24501 3485 24535 3519
rect 25973 3485 26007 3519
rect 27629 3485 27663 3519
rect 27813 3485 27847 3519
rect 27905 3485 27939 3519
rect 29561 3485 29595 3519
rect 29828 3485 29862 3519
rect 31217 3485 31251 3519
rect 31401 3485 31435 3519
rect 35822 3485 35856 3519
rect 36185 3485 36219 3519
rect 37933 3485 37967 3519
rect 39681 3485 39715 3519
rect 39865 3485 39899 3519
rect 42717 3485 42751 3519
rect 43085 3485 43119 3519
rect 43177 3485 43211 3519
rect 43709 3485 43743 3519
rect 45201 3485 45235 3519
rect 45560 3485 45594 3519
rect 47133 3485 47167 3519
rect 48044 3485 48078 3519
rect 49801 3485 49835 3519
rect 50425 3485 50459 3519
rect 52754 3485 52788 3519
rect 53021 3485 53055 3519
rect 54226 3485 54260 3519
rect 54861 3485 54895 3519
rect 55137 3485 55171 3519
rect 55321 3485 55355 3519
rect 58265 3485 58299 3519
rect 58357 3485 58391 3519
rect 58553 3485 58587 3519
rect 2728 3417 2762 3451
rect 3801 3417 3835 3451
rect 5080 3417 5114 3451
rect 7104 3417 7138 3451
rect 8585 3417 8619 3451
rect 9220 3417 9254 3451
rect 10517 3417 10551 3451
rect 10701 3417 10735 3451
rect 10793 3417 10827 3451
rect 12182 3417 12216 3451
rect 12808 3417 12842 3451
rect 17960 3417 17994 3451
rect 21364 3417 21398 3451
rect 23090 3417 23124 3451
rect 24746 3417 24780 3451
rect 26240 3417 26274 3451
rect 28150 3417 28184 3451
rect 31309 3417 31343 3451
rect 31738 3417 31772 3451
rect 33416 3417 33450 3451
rect 35449 3417 35483 3451
rect 35633 3417 35667 3451
rect 35725 3417 35759 3451
rect 36544 3417 36578 3451
rect 38200 3417 38234 3451
rect 40132 3417 40166 3451
rect 42472 3417 42506 3451
rect 43361 3417 43395 3451
rect 47409 3417 47443 3451
rect 55566 3417 55600 3451
rect 58020 3417 58054 3451
rect 1593 3349 1627 3383
rect 3525 3349 3559 3383
rect 4721 3349 4755 3383
rect 8217 3349 8251 3383
rect 10333 3349 10367 3383
rect 11069 3349 11103 3383
rect 16681 3349 16715 3383
rect 19257 3349 19291 3383
rect 24225 3349 24259 3383
rect 27353 3349 27387 3383
rect 27721 3349 27755 3383
rect 29285 3349 29319 3383
rect 32873 3349 32907 3383
rect 35357 3349 35391 3383
rect 36001 3349 36035 3383
rect 39497 3349 39531 3383
rect 41245 3349 41279 3383
rect 41337 3349 41371 3383
rect 42901 3349 42935 3383
rect 46673 3349 46707 3383
rect 49157 3349 49191 3383
rect 51549 3349 51583 3383
rect 51641 3349 51675 3383
rect 53113 3349 53147 3383
rect 56701 3349 56735 3383
rect 1685 3145 1719 3179
rect 2145 3145 2179 3179
rect 2513 3145 2547 3179
rect 3985 3145 4019 3179
rect 7849 3145 7883 3179
rect 8309 3145 8343 3179
rect 9137 3145 9171 3179
rect 11621 3145 11655 3179
rect 13553 3145 13587 3179
rect 14473 3145 14507 3179
rect 15945 3145 15979 3179
rect 16957 3145 16991 3179
rect 17969 3145 18003 3179
rect 19165 3145 19199 3179
rect 20913 3145 20947 3179
rect 21833 3145 21867 3179
rect 24041 3145 24075 3179
rect 25697 3145 25731 3179
rect 26985 3145 27019 3179
rect 31033 3145 31067 3179
rect 32229 3145 32263 3179
rect 33701 3145 33735 3179
rect 36093 3145 36127 3179
rect 37013 3145 37047 3179
rect 39037 3145 39071 3179
rect 42441 3145 42475 3179
rect 43361 3145 43395 3179
rect 46949 3145 46983 3179
rect 47593 3145 47627 3179
rect 52285 3145 52319 3179
rect 58541 3145 58575 3179
rect 9597 3077 9631 3111
rect 9781 3077 9815 3111
rect 9873 3077 9907 3111
rect 10793 3077 10827 3111
rect 14810 3077 14844 3111
rect 16037 3077 16071 3111
rect 21373 3077 21407 3111
rect 22661 3077 22695 3111
rect 22845 3077 22879 3111
rect 22937 3077 22971 3111
rect 33149 3077 33183 3111
rect 39589 3077 39623 3111
rect 46581 3077 46615 3111
rect 46765 3077 46799 3111
rect 48329 3077 48363 3111
rect 48513 3077 48547 3111
rect 48605 3077 48639 3111
rect 51457 3077 51491 3111
rect 51733 3077 51767 3111
rect 53481 3077 53515 3111
rect 53665 3077 53699 3111
rect 53757 3077 53791 3111
rect 1593 3009 1627 3043
rect 2605 3009 2639 3043
rect 4261 3009 4295 3043
rect 4629 3009 4663 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 7021 3009 7055 3043
rect 7113 3009 7147 3043
rect 7665 3009 7699 3043
rect 8401 3009 8435 3043
rect 9229 3009 9263 3043
rect 9970 3009 10004 3043
rect 10149 3009 10183 3043
rect 10517 3009 10551 3043
rect 11069 3009 11103 3043
rect 11805 3009 11839 3043
rect 12081 3009 12115 3043
rect 13737 3009 13771 3043
rect 14565 3009 14599 3043
rect 16221 3009 16255 3043
rect 16313 3009 16347 3043
rect 16410 3009 16444 3043
rect 17141 3009 17175 3043
rect 18153 3009 18187 3043
rect 18429 3009 18463 3043
rect 19257 3009 19291 3043
rect 21097 3009 21131 3043
rect 21260 3009 21294 3043
rect 21465 3009 21499 3043
rect 21649 3009 21683 3043
rect 23034 3009 23068 3043
rect 23949 3009 23983 3043
rect 24133 3009 24167 3043
rect 24225 3009 24259 3043
rect 26709 3009 26743 3043
rect 27721 3009 27755 3043
rect 29285 3009 29319 3043
rect 30941 3009 30975 3043
rect 31217 3009 31251 3043
rect 33415 3009 33449 3043
rect 33517 3009 33551 3043
rect 33885 3009 33919 3043
rect 34621 3009 34655 3043
rect 35909 3009 35943 3043
rect 36277 3009 36311 3043
rect 36369 3009 36403 3043
rect 36553 3009 36587 3043
rect 36829 3009 36863 3043
rect 37565 3009 37599 3043
rect 39221 3009 39255 3043
rect 39476 3009 39510 3043
rect 39681 3009 39715 3043
rect 39865 3009 39899 3043
rect 40969 3009 41003 3043
rect 43913 3009 43947 3043
rect 45293 3009 45327 3043
rect 46361 3009 46395 3043
rect 46489 3009 46523 3043
rect 47133 3009 47167 3043
rect 47225 3009 47259 3043
rect 48717 3031 48751 3065
rect 49157 3009 49191 3043
rect 51641 3009 51675 3043
rect 51861 3009 51895 3043
rect 52469 3009 52503 3043
rect 52745 3009 52779 3043
rect 53885 2999 53919 3033
rect 54033 3009 54067 3043
rect 57713 3009 57747 3043
rect 1869 2941 1903 2975
rect 2237 2941 2271 2975
rect 2354 2941 2388 2975
rect 3249 2941 3283 2975
rect 3433 2941 3467 2975
rect 6377 2941 6411 2975
rect 7389 2941 7423 2975
rect 8033 2941 8067 2975
rect 8125 2941 8159 2975
rect 8953 2941 8987 2975
rect 9873 2941 9907 2975
rect 10885 2941 10919 2975
rect 12541 2941 12575 2975
rect 13829 2941 13863 2975
rect 16129 2941 16163 2975
rect 17233 2941 17267 2975
rect 17877 2941 17911 2975
rect 18245 2941 18279 2975
rect 18613 2941 18647 2975
rect 19717 2941 19751 2975
rect 22385 2941 22419 2975
rect 22753 2941 22787 2975
rect 23765 2941 23799 2975
rect 24685 2941 24719 2975
rect 26249 2941 26283 2975
rect 27629 2941 27663 2975
rect 28273 2941 28307 2975
rect 28549 2941 28583 2975
rect 29653 2941 29687 2975
rect 31401 2941 31435 2975
rect 32873 2941 32907 2975
rect 34437 2941 34471 2975
rect 34897 2941 34931 2975
rect 35265 2941 35299 2975
rect 36461 2941 36495 2975
rect 37933 2941 37967 2975
rect 39773 2941 39807 2975
rect 40509 2941 40543 2975
rect 41245 2941 41279 2975
rect 42993 2941 43027 2975
rect 44281 2941 44315 2975
rect 45569 2941 45603 2975
rect 48145 2941 48179 2975
rect 48605 2941 48639 2975
rect 49525 2941 49559 2975
rect 50537 2941 50571 2975
rect 51457 2941 51491 2975
rect 53297 2941 53331 2975
rect 53757 2941 53791 2975
rect 54493 2941 54527 2975
rect 55505 2941 55539 2975
rect 57253 2941 57287 2975
rect 57989 2941 58023 2975
rect 6193 2873 6227 2907
rect 10333 2873 10367 2907
rect 21649 2873 21683 2907
rect 26525 2873 26559 2907
rect 30757 2873 30791 2907
rect 46213 2873 46247 2907
rect 5181 2805 5215 2839
rect 8217 2805 8251 2839
rect 10701 2805 10735 2839
rect 10793 2805 10827 2839
rect 11253 2805 11287 2839
rect 18429 2805 18463 2839
rect 23213 2805 23247 2839
rect 29101 2805 29135 2839
rect 31953 2805 31987 2839
rect 39957 2805 39991 2839
rect 46765 2805 46799 2839
rect 47409 2805 47443 2839
rect 51181 2805 51215 2839
rect 56149 2805 56183 2839
rect 4721 2601 4755 2635
rect 6561 2601 6595 2635
rect 7297 2601 7331 2635
rect 9781 2601 9815 2635
rect 12173 2601 12207 2635
rect 12265 2601 12299 2635
rect 14381 2601 14415 2635
rect 17509 2601 17543 2635
rect 20177 2601 20211 2635
rect 21833 2601 21867 2635
rect 24409 2601 24443 2635
rect 25329 2601 25363 2635
rect 27445 2601 27479 2635
rect 29101 2601 29135 2635
rect 29745 2601 29779 2635
rect 30481 2601 30515 2635
rect 33977 2601 34011 2635
rect 37105 2601 37139 2635
rect 39405 2601 39439 2635
rect 39681 2601 39715 2635
rect 41337 2601 41371 2635
rect 42073 2601 42107 2635
rect 43913 2601 43947 2635
rect 45017 2601 45051 2635
rect 47225 2601 47259 2635
rect 49801 2601 49835 2635
rect 50169 2601 50203 2635
rect 52193 2601 52227 2635
rect 55137 2601 55171 2635
rect 57253 2601 57287 2635
rect 57897 2601 57931 2635
rect 3985 2533 4019 2567
rect 14289 2533 14323 2567
rect 19441 2533 19475 2567
rect 32321 2533 32355 2567
rect 36369 2533 36403 2567
rect 44649 2533 44683 2567
rect 49709 2533 49743 2567
rect 55413 2533 55447 2567
rect 57529 2533 57563 2567
rect 1869 2465 1903 2499
rect 2789 2465 2823 2499
rect 10333 2465 10367 2499
rect 13461 2465 13495 2499
rect 15853 2465 15887 2499
rect 18061 2465 18095 2499
rect 20821 2465 20855 2499
rect 23029 2465 23063 2499
rect 25881 2465 25915 2499
rect 27997 2465 28031 2499
rect 31033 2465 31067 2499
rect 37749 2465 37783 2499
rect 40325 2465 40359 2499
rect 42901 2465 42935 2499
rect 45569 2465 45603 2499
rect 48053 2465 48087 2499
rect 53205 2465 53239 2499
rect 2053 2397 2087 2431
rect 2145 2397 2179 2431
rect 3801 2397 3835 2431
rect 4169 2397 4203 2431
rect 6193 2397 6227 2431
rect 6377 2397 6411 2431
rect 6745 2397 6779 2431
rect 8677 2397 8711 2431
rect 9229 2397 9263 2431
rect 10057 2397 10091 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 12449 2397 12483 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 15025 2397 15059 2431
rect 15209 2397 15243 2431
rect 16957 2397 16991 2431
rect 17601 2397 17635 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 22385 2397 22419 2431
rect 22569 2397 22603 2431
rect 24593 2397 24627 2431
rect 24777 2397 24811 2431
rect 25513 2397 25547 2431
rect 27072 2397 27106 2431
rect 27261 2397 27295 2431
rect 27445 2397 27479 2431
rect 27537 2397 27571 2431
rect 29285 2397 29319 2431
rect 29561 2397 29595 2431
rect 29929 2397 29963 2431
rect 30757 2397 30791 2431
rect 32137 2397 32171 2431
rect 33701 2397 33735 2431
rect 34161 2397 34195 2431
rect 34381 2397 34415 2431
rect 35909 2397 35943 2431
rect 36185 2397 36219 2431
rect 36553 2397 36587 2431
rect 37289 2397 37323 2431
rect 38761 2397 38795 2431
rect 39497 2397 39531 2431
rect 39681 2397 39715 2431
rect 39957 2397 39991 2431
rect 41889 2397 41923 2431
rect 42257 2397 42291 2431
rect 42441 2397 42475 2431
rect 44465 2397 44499 2431
rect 44833 2397 44867 2431
rect 46949 2397 46983 2431
rect 47409 2397 47443 2431
rect 47777 2397 47811 2431
rect 49065 2397 49099 2431
rect 49985 2397 50019 2431
rect 50353 2397 50387 2431
rect 52101 2397 52135 2431
rect 52377 2397 52411 2431
rect 52745 2397 52779 2431
rect 54217 2397 54251 2431
rect 54861 2397 54895 2431
rect 54953 2397 54987 2431
rect 55597 2397 55631 2431
rect 56885 2397 56919 2431
rect 57437 2397 57471 2431
rect 57713 2397 57747 2431
rect 58449 2397 58483 2431
rect 5273 2329 5307 2363
rect 7573 2329 7607 2363
rect 27169 2329 27203 2363
rect 32689 2329 32723 2363
rect 33977 2329 34011 2363
rect 34253 2329 34287 2363
rect 34897 2329 34931 2363
rect 45937 2329 45971 2363
rect 51089 2329 51123 2363
rect 55873 2329 55907 2363
<< metal1 >>
rect 1104 27770 58880 27792
rect 1104 27718 8172 27770
rect 8224 27718 8236 27770
rect 8288 27718 8300 27770
rect 8352 27718 8364 27770
rect 8416 27718 8428 27770
rect 8480 27718 22616 27770
rect 22668 27718 22680 27770
rect 22732 27718 22744 27770
rect 22796 27718 22808 27770
rect 22860 27718 22872 27770
rect 22924 27718 37060 27770
rect 37112 27718 37124 27770
rect 37176 27718 37188 27770
rect 37240 27718 37252 27770
rect 37304 27718 37316 27770
rect 37368 27718 51504 27770
rect 51556 27718 51568 27770
rect 51620 27718 51632 27770
rect 51684 27718 51696 27770
rect 51748 27718 51760 27770
rect 51812 27718 58880 27770
rect 1104 27696 58880 27718
rect 51350 27412 51356 27464
rect 51408 27452 51414 27464
rect 51629 27455 51687 27461
rect 51629 27452 51641 27455
rect 51408 27424 51641 27452
rect 51408 27412 51414 27424
rect 51629 27421 51641 27424
rect 51675 27421 51687 27455
rect 51629 27415 51687 27421
rect 51902 27276 51908 27328
rect 51960 27316 51966 27328
rect 52273 27319 52331 27325
rect 52273 27316 52285 27319
rect 51960 27288 52285 27316
rect 51960 27276 51966 27288
rect 52273 27285 52285 27288
rect 52319 27285 52331 27319
rect 52273 27279 52331 27285
rect 1104 27226 59040 27248
rect 1104 27174 15394 27226
rect 15446 27174 15458 27226
rect 15510 27174 15522 27226
rect 15574 27174 15586 27226
rect 15638 27174 15650 27226
rect 15702 27174 29838 27226
rect 29890 27174 29902 27226
rect 29954 27174 29966 27226
rect 30018 27174 30030 27226
rect 30082 27174 30094 27226
rect 30146 27174 44282 27226
rect 44334 27174 44346 27226
rect 44398 27174 44410 27226
rect 44462 27174 44474 27226
rect 44526 27174 44538 27226
rect 44590 27174 58726 27226
rect 58778 27174 58790 27226
rect 58842 27174 58854 27226
rect 58906 27174 58918 27226
rect 58970 27174 58982 27226
rect 59034 27174 59040 27226
rect 1104 27152 59040 27174
rect 30374 27004 30380 27056
rect 30432 27044 30438 27056
rect 31481 27047 31539 27053
rect 31481 27044 31493 27047
rect 30432 27016 31493 27044
rect 30432 27004 30438 27016
rect 31481 27013 31493 27016
rect 31527 27013 31539 27047
rect 31481 27007 31539 27013
rect 17310 26868 17316 26920
rect 17368 26908 17374 26920
rect 18601 26911 18659 26917
rect 18601 26908 18613 26911
rect 17368 26880 18613 26908
rect 17368 26868 17374 26880
rect 18601 26877 18613 26880
rect 18647 26877 18659 26911
rect 18601 26871 18659 26877
rect 28350 26868 28356 26920
rect 28408 26868 28414 26920
rect 28718 26868 28724 26920
rect 28776 26868 28782 26920
rect 29273 26911 29331 26917
rect 29273 26877 29285 26911
rect 29319 26908 29331 26911
rect 30190 26908 30196 26920
rect 29319 26880 30196 26908
rect 29319 26877 29331 26880
rect 29273 26871 29331 26877
rect 30190 26868 30196 26880
rect 30248 26868 30254 26920
rect 30282 26868 30288 26920
rect 30340 26908 30346 26920
rect 30745 26911 30803 26917
rect 30745 26908 30757 26911
rect 30340 26880 30757 26908
rect 30340 26868 30346 26880
rect 30745 26877 30757 26880
rect 30791 26877 30803 26911
rect 30745 26871 30803 26877
rect 45186 26868 45192 26920
rect 45244 26868 45250 26920
rect 46290 26868 46296 26920
rect 46348 26908 46354 26920
rect 46477 26911 46535 26917
rect 46477 26908 46489 26911
rect 46348 26880 46489 26908
rect 46348 26868 46354 26880
rect 46477 26877 46489 26880
rect 46523 26877 46535 26911
rect 46477 26871 46535 26877
rect 46658 26868 46664 26920
rect 46716 26868 46722 26920
rect 48130 26868 48136 26920
rect 48188 26868 48194 26920
rect 49234 26868 49240 26920
rect 49292 26868 49298 26920
rect 50798 26868 50804 26920
rect 50856 26868 50862 26920
rect 51074 26868 51080 26920
rect 51132 26868 51138 26920
rect 51994 26868 52000 26920
rect 52052 26908 52058 26920
rect 52273 26911 52331 26917
rect 52273 26908 52285 26911
rect 52052 26880 52285 26908
rect 52052 26868 52058 26880
rect 52273 26877 52285 26880
rect 52319 26877 52331 26911
rect 52273 26871 52331 26877
rect 54662 26868 54668 26920
rect 54720 26868 54726 26920
rect 45462 26800 45468 26852
rect 45520 26840 45526 26852
rect 45925 26843 45983 26849
rect 45925 26840 45937 26843
rect 45520 26812 45937 26840
rect 45520 26800 45526 26812
rect 45925 26809 45937 26812
rect 45971 26809 45983 26843
rect 45925 26803 45983 26809
rect 48222 26800 48228 26852
rect 48280 26840 48286 26852
rect 48685 26843 48743 26849
rect 48685 26840 48697 26843
rect 48280 26812 48697 26840
rect 48280 26800 48286 26812
rect 48685 26809 48697 26812
rect 48731 26809 48743 26843
rect 51721 26843 51779 26849
rect 51721 26840 51733 26843
rect 48685 26803 48743 26809
rect 51046 26812 51733 26840
rect 18509 26775 18567 26781
rect 18509 26741 18521 26775
rect 18555 26772 18567 26775
rect 18690 26772 18696 26784
rect 18555 26744 18696 26772
rect 18555 26741 18567 26744
rect 18509 26735 18567 26741
rect 18690 26732 18696 26744
rect 18748 26732 18754 26784
rect 18966 26732 18972 26784
rect 19024 26772 19030 26784
rect 19245 26775 19303 26781
rect 19245 26772 19257 26775
rect 19024 26744 19257 26772
rect 19024 26732 19030 26744
rect 19245 26741 19257 26744
rect 19291 26741 19303 26775
rect 19245 26735 19303 26741
rect 27798 26732 27804 26784
rect 27856 26732 27862 26784
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 30193 26775 30251 26781
rect 30193 26772 30205 26775
rect 30156 26744 30205 26772
rect 30156 26732 30162 26744
rect 30193 26741 30205 26744
rect 30239 26741 30251 26775
rect 30193 26735 30251 26741
rect 31202 26732 31208 26784
rect 31260 26732 31266 26784
rect 45830 26732 45836 26784
rect 45888 26732 45894 26784
rect 47302 26732 47308 26784
rect 47360 26732 47366 26784
rect 47578 26732 47584 26784
rect 47636 26732 47642 26784
rect 48593 26775 48651 26781
rect 48593 26741 48605 26775
rect 48639 26772 48651 26775
rect 48774 26772 48780 26784
rect 48639 26744 48780 26772
rect 48639 26741 48651 26744
rect 48593 26735 48651 26741
rect 48774 26732 48780 26744
rect 48832 26732 48838 26784
rect 50246 26732 50252 26784
rect 50304 26732 50310 26784
rect 50706 26732 50712 26784
rect 50764 26772 50770 26784
rect 51046 26772 51074 26812
rect 51721 26809 51733 26812
rect 51767 26809 51779 26843
rect 51721 26803 51779 26809
rect 50764 26744 51074 26772
rect 51629 26775 51687 26781
rect 50764 26732 50770 26744
rect 51629 26741 51641 26775
rect 51675 26772 51687 26775
rect 52086 26772 52092 26784
rect 51675 26744 52092 26772
rect 51675 26741 51687 26744
rect 51629 26735 51687 26741
rect 52086 26732 52092 26744
rect 52144 26732 52150 26784
rect 53834 26732 53840 26784
rect 53892 26772 53898 26784
rect 54113 26775 54171 26781
rect 54113 26772 54125 26775
rect 53892 26744 54125 26772
rect 53892 26732 53898 26744
rect 54113 26741 54125 26744
rect 54159 26741 54171 26775
rect 54113 26735 54171 26741
rect 1104 26682 58880 26704
rect 1104 26630 8172 26682
rect 8224 26630 8236 26682
rect 8288 26630 8300 26682
rect 8352 26630 8364 26682
rect 8416 26630 8428 26682
rect 8480 26630 22616 26682
rect 22668 26630 22680 26682
rect 22732 26630 22744 26682
rect 22796 26630 22808 26682
rect 22860 26630 22872 26682
rect 22924 26630 37060 26682
rect 37112 26630 37124 26682
rect 37176 26630 37188 26682
rect 37240 26630 37252 26682
rect 37304 26630 37316 26682
rect 37368 26630 51504 26682
rect 51556 26630 51568 26682
rect 51620 26630 51632 26682
rect 51684 26630 51696 26682
rect 51748 26630 51760 26682
rect 51812 26630 58880 26682
rect 1104 26608 58880 26630
rect 17310 26528 17316 26580
rect 17368 26528 17374 26580
rect 47857 26571 47915 26577
rect 47857 26537 47869 26571
rect 47903 26568 47915 26571
rect 48130 26568 48136 26580
rect 47903 26540 48136 26568
rect 47903 26537 47915 26540
rect 47857 26531 47915 26537
rect 48130 26528 48136 26540
rect 48188 26528 48194 26580
rect 48332 26540 48820 26568
rect 31205 26503 31263 26509
rect 31205 26469 31217 26503
rect 31251 26469 31263 26503
rect 31205 26463 31263 26469
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 18616 26404 19257 26432
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26333 15439 26367
rect 15381 26327 15439 26333
rect 18437 26367 18495 26373
rect 18437 26333 18449 26367
rect 18483 26364 18495 26367
rect 18616 26364 18644 26404
rect 19245 26401 19257 26404
rect 19291 26401 19303 26435
rect 31220 26432 31248 26463
rect 31849 26435 31907 26441
rect 31849 26432 31861 26435
rect 31220 26404 31861 26432
rect 19245 26395 19303 26401
rect 31849 26401 31861 26404
rect 31895 26401 31907 26435
rect 31849 26395 31907 26401
rect 48133 26435 48191 26441
rect 48133 26401 48145 26435
rect 48179 26432 48191 26435
rect 48332 26432 48360 26540
rect 48792 26512 48820 26540
rect 51350 26528 51356 26580
rect 51408 26568 51414 26580
rect 51537 26571 51595 26577
rect 51537 26568 51549 26571
rect 51408 26540 51549 26568
rect 51408 26528 51414 26540
rect 51537 26537 51549 26540
rect 51583 26537 51595 26571
rect 51537 26531 51595 26537
rect 48685 26503 48743 26509
rect 48685 26469 48697 26503
rect 48731 26469 48743 26503
rect 48685 26463 48743 26469
rect 48179 26404 48360 26432
rect 48700 26432 48728 26463
rect 48774 26460 48780 26512
rect 48832 26460 48838 26512
rect 53561 26503 53619 26509
rect 53561 26469 53573 26503
rect 53607 26500 53619 26503
rect 54662 26500 54668 26512
rect 53607 26472 54668 26500
rect 53607 26469 53619 26472
rect 53561 26463 53619 26469
rect 54662 26460 54668 26472
rect 54720 26460 54726 26512
rect 49329 26435 49387 26441
rect 49329 26432 49341 26435
rect 48700 26404 49341 26432
rect 48179 26401 48191 26404
rect 48133 26395 48191 26401
rect 49329 26401 49341 26404
rect 49375 26401 49387 26435
rect 49329 26395 49387 26401
rect 18483 26336 18644 26364
rect 18693 26367 18751 26373
rect 18483 26333 18495 26336
rect 18437 26327 18495 26333
rect 18693 26333 18705 26367
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 15102 26188 15108 26240
rect 15160 26228 15166 26240
rect 15396 26228 15424 26327
rect 15648 26299 15706 26305
rect 15648 26265 15660 26299
rect 15694 26296 15706 26299
rect 15838 26296 15844 26308
rect 15694 26268 15844 26296
rect 15694 26265 15706 26268
rect 15648 26259 15706 26265
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 17129 26299 17187 26305
rect 17129 26265 17141 26299
rect 17175 26296 17187 26299
rect 17862 26296 17868 26308
rect 17175 26268 17868 26296
rect 17175 26265 17187 26268
rect 17129 26259 17187 26265
rect 17862 26256 17868 26268
rect 17920 26256 17926 26308
rect 18708 26296 18736 26327
rect 19794 26324 19800 26376
rect 19852 26324 19858 26376
rect 27893 26367 27951 26373
rect 27893 26333 27905 26367
rect 27939 26364 27951 26367
rect 29638 26364 29644 26376
rect 27939 26336 29644 26364
rect 27939 26333 27951 26336
rect 27893 26327 27951 26333
rect 22462 26296 22468 26308
rect 18708 26268 22468 26296
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 15160 26200 15424 26228
rect 15160 26188 15166 26200
rect 16758 26188 16764 26240
rect 16816 26188 16822 26240
rect 17310 26188 17316 26240
rect 17368 26228 17374 26240
rect 18969 26231 19027 26237
rect 18969 26228 18981 26231
rect 17368 26200 18981 26228
rect 17368 26188 17374 26200
rect 18969 26197 18981 26200
rect 19015 26197 19027 26231
rect 18969 26191 19027 26197
rect 27614 26188 27620 26240
rect 27672 26228 27678 26240
rect 27908 26228 27936 26327
rect 29638 26324 29644 26336
rect 29696 26364 29702 26376
rect 30098 26373 30104 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29696 26336 29837 26364
rect 29696 26324 29702 26336
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 30092 26364 30104 26373
rect 30059 26336 30104 26364
rect 29825 26327 29883 26333
rect 30092 26327 30104 26336
rect 30098 26324 30104 26327
rect 30156 26324 30162 26376
rect 45005 26367 45063 26373
rect 45005 26333 45017 26367
rect 45051 26364 45063 26367
rect 46477 26367 46535 26373
rect 46477 26364 46489 26367
rect 45051 26336 46489 26364
rect 45051 26333 45063 26336
rect 45005 26327 45063 26333
rect 46477 26333 46489 26336
rect 46523 26364 46535 26367
rect 46566 26364 46572 26376
rect 46523 26336 46572 26364
rect 46523 26333 46535 26336
rect 46477 26327 46535 26333
rect 46566 26324 46572 26336
rect 46624 26324 46630 26376
rect 46744 26367 46802 26373
rect 46744 26333 46756 26367
rect 46790 26364 46802 26367
rect 47302 26364 47308 26376
rect 46790 26336 47308 26364
rect 46790 26333 46802 26336
rect 46744 26327 46802 26333
rect 47302 26324 47308 26336
rect 47360 26324 47366 26376
rect 48222 26324 48228 26376
rect 48280 26364 48286 26376
rect 48317 26367 48375 26373
rect 48317 26364 48329 26367
rect 48280 26336 48329 26364
rect 48280 26324 48286 26336
rect 48317 26333 48329 26336
rect 48363 26333 48375 26367
rect 48317 26327 48375 26333
rect 49878 26324 49884 26376
rect 49936 26364 49942 26376
rect 50157 26367 50215 26373
rect 50157 26364 50169 26367
rect 49936 26336 50169 26364
rect 49936 26324 49942 26336
rect 50157 26333 50169 26336
rect 50203 26364 50215 26367
rect 52181 26367 52239 26373
rect 52181 26364 52193 26367
rect 50203 26336 52193 26364
rect 50203 26333 50215 26336
rect 50157 26327 50215 26333
rect 52181 26333 52193 26336
rect 52227 26364 52239 26367
rect 52227 26336 52408 26364
rect 52227 26333 52239 26336
rect 52181 26327 52239 26333
rect 28160 26299 28218 26305
rect 28160 26265 28172 26299
rect 28206 26296 28218 26299
rect 28442 26296 28448 26308
rect 28206 26268 28448 26296
rect 28206 26265 28218 26268
rect 28160 26259 28218 26265
rect 28442 26256 28448 26268
rect 28500 26256 28506 26308
rect 44174 26256 44180 26308
rect 44232 26296 44238 26308
rect 44729 26299 44787 26305
rect 44729 26296 44741 26299
rect 44232 26268 44741 26296
rect 44232 26256 44238 26268
rect 44729 26265 44741 26268
rect 44775 26296 44787 26299
rect 45272 26299 45330 26305
rect 44775 26268 45232 26296
rect 44775 26265 44787 26268
rect 44729 26259 44787 26265
rect 27672 26200 27936 26228
rect 27672 26188 27678 26200
rect 29270 26188 29276 26240
rect 29328 26188 29334 26240
rect 30834 26188 30840 26240
rect 30892 26228 30898 26240
rect 31297 26231 31355 26237
rect 31297 26228 31309 26231
rect 30892 26200 31309 26228
rect 30892 26188 30898 26200
rect 31297 26197 31309 26200
rect 31343 26197 31355 26231
rect 31297 26191 31355 26197
rect 31570 26188 31576 26240
rect 31628 26228 31634 26240
rect 32217 26231 32275 26237
rect 32217 26228 32229 26231
rect 31628 26200 32229 26228
rect 31628 26188 31634 26200
rect 32217 26197 32229 26200
rect 32263 26197 32275 26231
rect 45204 26228 45232 26268
rect 45272 26265 45284 26299
rect 45318 26296 45330 26299
rect 45370 26296 45376 26308
rect 45318 26268 45376 26296
rect 45318 26265 45330 26268
rect 45272 26259 45330 26265
rect 45370 26256 45376 26268
rect 45428 26256 45434 26308
rect 48130 26256 48136 26308
rect 48188 26296 48194 26308
rect 48777 26299 48835 26305
rect 48777 26296 48789 26299
rect 48188 26268 48789 26296
rect 48188 26256 48194 26268
rect 48777 26265 48789 26268
rect 48823 26265 48835 26299
rect 48777 26259 48835 26265
rect 50424 26299 50482 26305
rect 50424 26265 50436 26299
rect 50470 26296 50482 26299
rect 50706 26296 50712 26308
rect 50470 26268 50712 26296
rect 50470 26265 50482 26268
rect 50424 26259 50482 26265
rect 50706 26256 50712 26268
rect 50764 26256 50770 26308
rect 52380 26240 52408 26336
rect 54202 26324 54208 26376
rect 54260 26324 54266 26376
rect 54386 26324 54392 26376
rect 54444 26324 54450 26376
rect 52448 26299 52506 26305
rect 52448 26265 52460 26299
rect 52494 26296 52506 26299
rect 53653 26299 53711 26305
rect 53653 26296 53665 26299
rect 52494 26268 53665 26296
rect 52494 26265 52506 26268
rect 52448 26259 52506 26265
rect 53653 26265 53665 26268
rect 53699 26265 53711 26299
rect 53653 26259 53711 26265
rect 45738 26228 45744 26240
rect 45204 26200 45744 26228
rect 32217 26191 32275 26197
rect 45738 26188 45744 26200
rect 45796 26188 45802 26240
rect 46382 26188 46388 26240
rect 46440 26188 46446 26240
rect 46842 26188 46848 26240
rect 46900 26228 46906 26240
rect 48225 26231 48283 26237
rect 48225 26228 48237 26231
rect 46900 26200 48237 26228
rect 46900 26188 46906 26200
rect 48225 26197 48237 26200
rect 48271 26197 48283 26231
rect 48225 26191 48283 26197
rect 48590 26188 48596 26240
rect 48648 26228 48654 26240
rect 51350 26228 51356 26240
rect 48648 26200 51356 26228
rect 48648 26188 48654 26200
rect 51350 26188 51356 26200
rect 51408 26228 51414 26240
rect 51813 26231 51871 26237
rect 51813 26228 51825 26231
rect 51408 26200 51825 26228
rect 51408 26188 51414 26200
rect 51813 26197 51825 26200
rect 51859 26197 51871 26231
rect 51813 26191 51871 26197
rect 52362 26188 52368 26240
rect 52420 26188 52426 26240
rect 54570 26188 54576 26240
rect 54628 26228 54634 26240
rect 55033 26231 55091 26237
rect 55033 26228 55045 26231
rect 54628 26200 55045 26228
rect 54628 26188 54634 26200
rect 55033 26197 55045 26200
rect 55079 26197 55091 26231
rect 55033 26191 55091 26197
rect 1104 26138 59040 26160
rect 1104 26086 15394 26138
rect 15446 26086 15458 26138
rect 15510 26086 15522 26138
rect 15574 26086 15586 26138
rect 15638 26086 15650 26138
rect 15702 26086 29838 26138
rect 29890 26086 29902 26138
rect 29954 26086 29966 26138
rect 30018 26086 30030 26138
rect 30082 26086 30094 26138
rect 30146 26086 44282 26138
rect 44334 26086 44346 26138
rect 44398 26086 44410 26138
rect 44462 26086 44474 26138
rect 44526 26086 44538 26138
rect 44590 26086 58726 26138
rect 58778 26086 58790 26138
rect 58842 26086 58854 26138
rect 58906 26086 58918 26138
rect 58970 26086 58982 26138
rect 59034 26086 59040 26138
rect 1104 26064 59040 26086
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 19429 26027 19487 26033
rect 16540 25996 19104 26024
rect 16540 25984 16546 25996
rect 19076 25965 19104 25996
rect 19429 25993 19441 26027
rect 19475 26024 19487 26027
rect 19794 26024 19800 26036
rect 19475 25996 19800 26024
rect 19475 25993 19487 25996
rect 19429 25987 19487 25993
rect 19794 25984 19800 25996
rect 19852 25984 19858 26036
rect 28902 25984 28908 26036
rect 28960 26024 28966 26036
rect 29638 26024 29644 26036
rect 28960 25996 29644 26024
rect 28960 25984 28966 25996
rect 29638 25984 29644 25996
rect 29696 25984 29702 26036
rect 29822 25984 29828 26036
rect 29880 26024 29886 26036
rect 31481 26027 31539 26033
rect 31481 26024 31493 26027
rect 29880 25996 31493 26024
rect 29880 25984 29886 25996
rect 31481 25993 31493 25996
rect 31527 25993 31539 26027
rect 31481 25987 31539 25993
rect 44177 26027 44235 26033
rect 44177 25993 44189 26027
rect 44223 26024 44235 26027
rect 45186 26024 45192 26036
rect 44223 25996 45192 26024
rect 44223 25993 44235 25996
rect 44177 25987 44235 25993
rect 45186 25984 45192 25996
rect 45244 25984 45250 26036
rect 45830 25984 45836 26036
rect 45888 26024 45894 26036
rect 46017 26027 46075 26033
rect 46017 26024 46029 26027
rect 45888 25996 46029 26024
rect 45888 25984 45894 25996
rect 46017 25993 46029 25996
rect 46063 25993 46075 26027
rect 46017 25987 46075 25993
rect 46290 25984 46296 26036
rect 46348 26024 46354 26036
rect 46385 26027 46443 26033
rect 46385 26024 46397 26027
rect 46348 25996 46397 26024
rect 46348 25984 46354 25996
rect 46385 25993 46397 25996
rect 46431 25993 46443 26027
rect 46385 25987 46443 25993
rect 46477 26027 46535 26033
rect 46477 25993 46489 26027
rect 46523 26024 46535 26027
rect 46658 26024 46664 26036
rect 46523 25996 46664 26024
rect 46523 25993 46535 25996
rect 46477 25987 46535 25993
rect 46658 25984 46664 25996
rect 46716 25984 46722 26036
rect 46842 25984 46848 26036
rect 46900 25984 46906 26036
rect 46937 26027 46995 26033
rect 46937 25993 46949 26027
rect 46983 26024 46995 26027
rect 47578 26024 47584 26036
rect 46983 25996 47584 26024
rect 46983 25993 46995 25996
rect 46937 25987 46995 25993
rect 47578 25984 47584 25996
rect 47636 25984 47642 26036
rect 48961 26027 49019 26033
rect 48961 25993 48973 26027
rect 49007 26024 49019 26027
rect 49234 26024 49240 26036
rect 49007 25996 49240 26024
rect 49007 25993 49019 25996
rect 48961 25987 49019 25993
rect 49234 25984 49240 25996
rect 49292 25984 49298 26036
rect 51074 25984 51080 26036
rect 51132 26024 51138 26036
rect 51169 26027 51227 26033
rect 51169 26024 51181 26027
rect 51132 25996 51181 26024
rect 51132 25984 51138 25996
rect 51169 25993 51181 25996
rect 51215 25993 51227 26027
rect 51169 25987 51227 25993
rect 51994 25984 52000 26036
rect 52052 25984 52058 26036
rect 54113 26027 54171 26033
rect 54113 25993 54125 26027
rect 54159 25993 54171 26027
rect 54113 25987 54171 25993
rect 54205 26027 54263 26033
rect 54205 25993 54217 26027
rect 54251 26024 54263 26027
rect 54478 26024 54484 26036
rect 54251 25996 54484 26024
rect 54251 25993 54263 25996
rect 54205 25987 54263 25993
rect 27798 25965 27804 25968
rect 14921 25959 14979 25965
rect 14921 25925 14933 25959
rect 14967 25956 14979 25959
rect 15258 25959 15316 25965
rect 15258 25956 15270 25959
rect 14967 25928 15270 25956
rect 14967 25925 14979 25928
rect 14921 25919 14979 25925
rect 15258 25925 15270 25928
rect 15304 25925 15316 25959
rect 15258 25919 15316 25925
rect 19061 25959 19119 25965
rect 19061 25925 19073 25959
rect 19107 25956 19119 25959
rect 27792 25956 27804 25965
rect 19107 25928 19840 25956
rect 27759 25928 27804 25956
rect 19107 25925 19119 25928
rect 19061 25919 19119 25925
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25888 15071 25891
rect 15102 25888 15108 25900
rect 15059 25860 15108 25888
rect 15059 25857 15071 25860
rect 15013 25851 15071 25857
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 19812 25897 19840 25928
rect 27792 25919 27804 25928
rect 27798 25916 27804 25919
rect 27856 25916 27862 25968
rect 45312 25959 45370 25965
rect 45312 25925 45324 25959
rect 45358 25956 45370 25959
rect 45462 25956 45468 25968
rect 45358 25928 45468 25956
rect 45358 25925 45370 25928
rect 45312 25919 45370 25925
rect 45462 25916 45468 25928
rect 45520 25916 45526 25968
rect 46566 25956 46572 25968
rect 45572 25928 46572 25956
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 18969 25891 19027 25897
rect 18969 25888 18981 25891
rect 18371 25860 18981 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 18969 25857 18981 25860
rect 19015 25888 19027 25891
rect 19797 25891 19855 25897
rect 19015 25860 19288 25888
rect 19015 25857 19027 25860
rect 18969 25851 19027 25857
rect 19260 25832 19288 25860
rect 19797 25857 19809 25891
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25888 27583 25891
rect 27614 25888 27620 25900
rect 27571 25860 27620 25888
rect 27571 25857 27583 25860
rect 27525 25851 27583 25857
rect 27614 25848 27620 25860
rect 27672 25848 27678 25900
rect 29914 25848 29920 25900
rect 29972 25848 29978 25900
rect 30006 25848 30012 25900
rect 30064 25897 30070 25900
rect 45572 25897 45600 25928
rect 46566 25916 46572 25928
rect 46624 25956 46630 25968
rect 50056 25959 50114 25965
rect 46624 25928 49832 25956
rect 46624 25916 46630 25928
rect 30064 25891 30113 25897
rect 30064 25857 30067 25891
rect 30101 25857 30113 25891
rect 31113 25891 31171 25897
rect 31113 25888 31125 25891
rect 30064 25851 30113 25857
rect 30852 25860 31125 25888
rect 30064 25848 30070 25851
rect 30852 25832 30880 25860
rect 31113 25857 31125 25860
rect 31159 25857 31171 25891
rect 31573 25891 31631 25897
rect 31573 25888 31585 25891
rect 31113 25851 31171 25857
rect 31220 25860 31585 25888
rect 7006 25780 7012 25832
rect 7064 25780 7070 25832
rect 7742 25780 7748 25832
rect 7800 25780 7806 25832
rect 8018 25780 8024 25832
rect 8076 25820 8082 25832
rect 8481 25823 8539 25829
rect 8481 25820 8493 25823
rect 8076 25792 8493 25820
rect 8076 25780 8082 25792
rect 8481 25789 8493 25792
rect 8527 25789 8539 25823
rect 8481 25783 8539 25789
rect 10962 25780 10968 25832
rect 11020 25780 11026 25832
rect 13814 25780 13820 25832
rect 13872 25780 13878 25832
rect 14366 25780 14372 25832
rect 14424 25780 14430 25832
rect 17310 25780 17316 25832
rect 17368 25780 17374 25832
rect 17402 25780 17408 25832
rect 17460 25829 17466 25832
rect 17460 25823 17509 25829
rect 17460 25789 17463 25823
rect 17497 25789 17509 25823
rect 17460 25783 17509 25789
rect 17460 25780 17466 25783
rect 17586 25780 17592 25832
rect 17644 25780 17650 25832
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 11793 25755 11851 25761
rect 11793 25721 11805 25755
rect 11839 25752 11851 25755
rect 12434 25752 12440 25764
rect 11839 25724 12440 25752
rect 11839 25721 11851 25724
rect 11793 25715 11851 25721
rect 12434 25712 12440 25724
rect 12492 25712 12498 25764
rect 13170 25752 13176 25764
rect 12820 25724 13176 25752
rect 6454 25644 6460 25696
rect 6512 25644 6518 25696
rect 7190 25644 7196 25696
rect 7248 25644 7254 25696
rect 7926 25644 7932 25696
rect 7984 25644 7990 25696
rect 8846 25644 8852 25696
rect 8904 25644 8910 25696
rect 10410 25644 10416 25696
rect 10468 25644 10474 25696
rect 12161 25687 12219 25693
rect 12161 25653 12173 25687
rect 12207 25684 12219 25687
rect 12820 25684 12848 25724
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 17862 25712 17868 25764
rect 17920 25712 17926 25764
rect 18524 25752 18552 25783
rect 18690 25780 18696 25832
rect 18748 25820 18754 25832
rect 19153 25823 19211 25829
rect 19153 25820 19165 25823
rect 18748 25792 19165 25820
rect 18748 25780 18754 25792
rect 19153 25789 19165 25792
rect 19199 25789 19211 25823
rect 19153 25783 19211 25789
rect 19242 25780 19248 25832
rect 19300 25780 19306 25832
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25789 19947 25823
rect 19889 25783 19947 25789
rect 20073 25823 20131 25829
rect 20073 25789 20085 25823
rect 20119 25820 20131 25823
rect 20119 25792 20484 25820
rect 20119 25789 20131 25792
rect 20073 25783 20131 25789
rect 18966 25752 18972 25764
rect 18524 25724 18972 25752
rect 18966 25712 18972 25724
rect 19024 25752 19030 25764
rect 19904 25752 19932 25783
rect 19024 25724 19932 25752
rect 19024 25712 19030 25724
rect 20456 25696 20484 25792
rect 28718 25780 28724 25832
rect 28776 25780 28782 25832
rect 29546 25780 29552 25832
rect 29604 25820 29610 25832
rect 30193 25823 30251 25829
rect 30193 25820 30205 25823
rect 29604 25792 30205 25820
rect 29604 25780 29610 25792
rect 30193 25789 30205 25792
rect 30239 25789 30251 25823
rect 30193 25783 30251 25789
rect 30834 25780 30840 25832
rect 30892 25780 30898 25832
rect 30929 25823 30987 25829
rect 30929 25789 30941 25823
rect 30975 25820 30987 25823
rect 31220 25820 31248 25860
rect 31573 25857 31585 25860
rect 31619 25888 31631 25891
rect 45557 25891 45615 25897
rect 31619 25860 31708 25888
rect 31619 25857 31631 25860
rect 31573 25851 31631 25857
rect 30975 25792 31248 25820
rect 30975 25789 30987 25792
rect 30929 25783 30987 25789
rect 31294 25780 31300 25832
rect 31352 25780 31358 25832
rect 28736 25752 28764 25780
rect 28905 25755 28963 25761
rect 28905 25752 28917 25755
rect 28736 25724 28917 25752
rect 28905 25721 28917 25724
rect 28951 25721 28963 25755
rect 28905 25715 28963 25721
rect 30469 25755 30527 25761
rect 30469 25721 30481 25755
rect 30515 25752 30527 25755
rect 31570 25752 31576 25764
rect 30515 25724 31576 25752
rect 30515 25721 30527 25724
rect 30469 25715 30527 25721
rect 31570 25712 31576 25724
rect 31628 25712 31634 25764
rect 31680 25696 31708 25860
rect 45557 25857 45569 25891
rect 45603 25857 45615 25891
rect 45557 25851 45615 25857
rect 45646 25848 45652 25900
rect 45704 25888 45710 25900
rect 45925 25891 45983 25897
rect 45925 25888 45937 25891
rect 45704 25860 45937 25888
rect 45704 25848 45710 25860
rect 45925 25857 45937 25860
rect 45971 25888 45983 25891
rect 46842 25888 46848 25900
rect 45971 25860 46848 25888
rect 45971 25857 45983 25860
rect 45925 25851 45983 25857
rect 46842 25848 46848 25860
rect 46900 25848 46906 25900
rect 47596 25897 47624 25928
rect 47581 25891 47639 25897
rect 47581 25857 47593 25891
rect 47627 25857 47639 25891
rect 47581 25851 47639 25857
rect 47848 25891 47906 25897
rect 47848 25857 47860 25891
rect 47894 25888 47906 25891
rect 48130 25888 48136 25900
rect 47894 25860 48136 25888
rect 47894 25857 47906 25860
rect 47848 25851 47906 25857
rect 48130 25848 48136 25860
rect 48188 25848 48194 25900
rect 48590 25848 48596 25900
rect 48648 25848 48654 25900
rect 49804 25897 49832 25928
rect 50056 25925 50068 25959
rect 50102 25956 50114 25959
rect 50246 25956 50252 25968
rect 50102 25928 50252 25956
rect 50102 25925 50114 25928
rect 50056 25919 50114 25925
rect 50246 25916 50252 25928
rect 50304 25916 50310 25968
rect 53000 25959 53058 25965
rect 51552 25928 52491 25956
rect 49789 25891 49847 25897
rect 49789 25857 49801 25891
rect 49835 25888 49847 25891
rect 49878 25888 49884 25900
rect 49835 25860 49884 25888
rect 49835 25857 49847 25860
rect 49789 25851 49847 25857
rect 49878 25848 49884 25860
rect 49936 25848 49942 25900
rect 50890 25848 50896 25900
rect 50948 25888 50954 25900
rect 51552 25897 51580 25928
rect 51537 25891 51595 25897
rect 51537 25888 51549 25891
rect 50948 25860 51549 25888
rect 50948 25848 50954 25860
rect 51537 25857 51549 25860
rect 51583 25857 51595 25891
rect 51537 25851 51595 25857
rect 51629 25891 51687 25897
rect 51629 25857 51641 25891
rect 51675 25888 51687 25891
rect 51902 25888 51908 25900
rect 51675 25860 51908 25888
rect 51675 25857 51687 25860
rect 51629 25851 51687 25857
rect 51902 25848 51908 25860
rect 51960 25888 51966 25900
rect 52270 25888 52276 25900
rect 51960 25860 52276 25888
rect 51960 25848 51966 25860
rect 52270 25848 52276 25860
rect 52328 25848 52334 25900
rect 52365 25891 52423 25897
rect 52365 25857 52377 25891
rect 52411 25857 52423 25891
rect 52463 25888 52491 25928
rect 53000 25925 53012 25959
rect 53046 25956 53058 25959
rect 53834 25956 53840 25968
rect 53046 25928 53840 25956
rect 53046 25925 53058 25928
rect 53000 25919 53058 25925
rect 53834 25916 53840 25928
rect 53892 25916 53898 25968
rect 54128 25956 54156 25987
rect 54478 25984 54484 25996
rect 54536 25984 54542 26036
rect 54386 25956 54392 25968
rect 54128 25928 54392 25956
rect 54386 25916 54392 25928
rect 54444 25916 54450 25968
rect 52463 25860 53788 25888
rect 52365 25851 52423 25857
rect 32677 25823 32735 25829
rect 32677 25820 32689 25823
rect 31956 25792 32689 25820
rect 31956 25761 31984 25792
rect 32677 25789 32689 25792
rect 32723 25789 32735 25823
rect 32677 25783 32735 25789
rect 45738 25780 45744 25832
rect 45796 25780 45802 25832
rect 46658 25780 46664 25832
rect 46716 25820 46722 25832
rect 47029 25823 47087 25829
rect 47029 25820 47041 25823
rect 46716 25792 47041 25820
rect 46716 25780 46722 25792
rect 47029 25789 47041 25792
rect 47075 25789 47087 25823
rect 47029 25783 47087 25789
rect 31941 25755 31999 25761
rect 31941 25721 31953 25755
rect 31987 25721 31999 25755
rect 31941 25715 31999 25721
rect 12207 25656 12848 25684
rect 12207 25653 12219 25656
rect 12161 25647 12219 25653
rect 12894 25644 12900 25696
rect 12952 25684 12958 25696
rect 13265 25687 13323 25693
rect 13265 25684 13277 25687
rect 12952 25656 13277 25684
rect 12952 25644 12958 25656
rect 13265 25653 13277 25656
rect 13311 25653 13323 25687
rect 13265 25647 13323 25653
rect 16393 25687 16451 25693
rect 16393 25653 16405 25687
rect 16439 25684 16451 25687
rect 16574 25684 16580 25696
rect 16439 25656 16580 25684
rect 16439 25653 16451 25656
rect 16393 25647 16451 25653
rect 16574 25644 16580 25656
rect 16632 25644 16638 25696
rect 16669 25687 16727 25693
rect 16669 25653 16681 25687
rect 16715 25684 16727 25687
rect 17494 25684 17500 25696
rect 16715 25656 17500 25684
rect 16715 25653 16727 25656
rect 16669 25647 16727 25653
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 18598 25644 18604 25696
rect 18656 25644 18662 25696
rect 20438 25644 20444 25696
rect 20496 25644 20502 25696
rect 29273 25687 29331 25693
rect 29273 25653 29285 25687
rect 29319 25684 29331 25687
rect 30650 25684 30656 25696
rect 29319 25656 30656 25684
rect 29319 25653 29331 25656
rect 29273 25647 29331 25653
rect 30650 25644 30656 25656
rect 30708 25644 30714 25696
rect 31662 25644 31668 25696
rect 31720 25644 31726 25696
rect 32122 25644 32128 25696
rect 32180 25644 32186 25696
rect 46014 25644 46020 25696
rect 46072 25684 46078 25696
rect 48608 25684 48636 25848
rect 51258 25780 51264 25832
rect 51316 25780 51322 25832
rect 51350 25780 51356 25832
rect 51408 25780 51414 25832
rect 51994 25780 52000 25832
rect 52052 25820 52058 25832
rect 52380 25820 52408 25851
rect 52052 25792 52408 25820
rect 52733 25823 52791 25829
rect 52052 25780 52058 25792
rect 52733 25789 52745 25823
rect 52779 25789 52791 25823
rect 53760 25820 53788 25860
rect 54570 25848 54576 25900
rect 54628 25848 54634 25900
rect 54665 25823 54723 25829
rect 54665 25820 54677 25823
rect 53760 25792 54677 25820
rect 52733 25783 52791 25789
rect 54665 25789 54677 25792
rect 54711 25789 54723 25823
rect 54665 25783 54723 25789
rect 54757 25823 54815 25829
rect 54757 25789 54769 25823
rect 54803 25820 54815 25823
rect 55217 25823 55275 25829
rect 55217 25820 55229 25823
rect 54803 25792 55229 25820
rect 54803 25789 54815 25792
rect 54757 25783 54815 25789
rect 55217 25789 55229 25792
rect 55263 25789 55275 25823
rect 55217 25783 55275 25789
rect 51276 25752 51304 25780
rect 52362 25752 52368 25764
rect 51276 25724 52368 25752
rect 52362 25712 52368 25724
rect 52420 25752 52426 25764
rect 52748 25752 52776 25783
rect 54772 25752 54800 25783
rect 52420 25724 52776 25752
rect 54680 25724 54800 25752
rect 52420 25712 52426 25724
rect 46072 25656 48636 25684
rect 46072 25644 46078 25656
rect 48774 25644 48780 25696
rect 48832 25684 48838 25696
rect 54680 25684 54708 25724
rect 48832 25656 54708 25684
rect 48832 25644 48838 25656
rect 1104 25594 58880 25616
rect 1104 25542 8172 25594
rect 8224 25542 8236 25594
rect 8288 25542 8300 25594
rect 8352 25542 8364 25594
rect 8416 25542 8428 25594
rect 8480 25542 22616 25594
rect 22668 25542 22680 25594
rect 22732 25542 22744 25594
rect 22796 25542 22808 25594
rect 22860 25542 22872 25594
rect 22924 25542 37060 25594
rect 37112 25542 37124 25594
rect 37176 25542 37188 25594
rect 37240 25542 37252 25594
rect 37304 25542 37316 25594
rect 37368 25542 51504 25594
rect 51556 25542 51568 25594
rect 51620 25542 51632 25594
rect 51684 25542 51696 25594
rect 51748 25542 51760 25594
rect 51812 25542 58880 25594
rect 1104 25520 58880 25542
rect 7742 25440 7748 25492
rect 7800 25440 7806 25492
rect 7929 25483 7987 25489
rect 7929 25449 7941 25483
rect 7975 25480 7987 25483
rect 8018 25480 8024 25492
rect 7975 25452 8024 25480
rect 7975 25449 7987 25452
rect 7929 25443 7987 25449
rect 8018 25440 8024 25452
rect 8076 25440 8082 25492
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10962 25480 10968 25492
rect 10643 25452 10968 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 14274 25480 14280 25492
rect 12360 25452 14280 25480
rect 10505 25415 10563 25421
rect 10505 25381 10517 25415
rect 10551 25412 10563 25415
rect 12360 25412 12388 25452
rect 14274 25440 14280 25452
rect 14332 25440 14338 25492
rect 14366 25440 14372 25492
rect 14424 25480 14430 25492
rect 15197 25483 15255 25489
rect 15197 25480 15209 25483
rect 14424 25452 15209 25480
rect 14424 25440 14430 25452
rect 15197 25449 15209 25452
rect 15243 25449 15255 25483
rect 17954 25480 17960 25492
rect 15197 25443 15255 25449
rect 16592 25452 17960 25480
rect 10551 25384 12388 25412
rect 13725 25415 13783 25421
rect 10551 25381 10563 25384
rect 10505 25375 10563 25381
rect 8018 25304 8024 25356
rect 8076 25344 8082 25356
rect 8481 25347 8539 25353
rect 8481 25344 8493 25347
rect 8076 25316 8493 25344
rect 8076 25304 8082 25316
rect 8481 25313 8493 25316
rect 8527 25344 8539 25347
rect 8846 25344 8852 25356
rect 8527 25316 8852 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 8846 25304 8852 25316
rect 8904 25304 8910 25356
rect 11256 25353 11284 25384
rect 13725 25381 13737 25415
rect 13771 25412 13783 25415
rect 16592 25412 16620 25452
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 19242 25440 19248 25492
rect 19300 25440 19306 25492
rect 27801 25483 27859 25489
rect 27801 25449 27813 25483
rect 27847 25480 27859 25483
rect 28350 25480 28356 25492
rect 27847 25452 28356 25480
rect 27847 25449 27859 25452
rect 27801 25443 27859 25449
rect 28350 25440 28356 25452
rect 28408 25440 28414 25492
rect 28460 25452 29224 25480
rect 17586 25412 17592 25424
rect 13771 25384 14136 25412
rect 13771 25381 13783 25384
rect 13725 25375 13783 25381
rect 14108 25353 14136 25384
rect 15028 25384 16620 25412
rect 11241 25347 11299 25353
rect 11241 25313 11253 25347
rect 11287 25344 11299 25347
rect 14093 25347 14151 25353
rect 11287 25316 11321 25344
rect 11287 25313 11299 25316
rect 11241 25307 11299 25313
rect 14093 25313 14105 25347
rect 14139 25313 14151 25347
rect 14093 25307 14151 25313
rect 5534 25236 5540 25288
rect 5592 25236 5598 25288
rect 6362 25236 6368 25288
rect 6420 25236 6426 25288
rect 6454 25236 6460 25288
rect 6512 25276 6518 25288
rect 6621 25279 6679 25285
rect 6621 25276 6633 25279
rect 6512 25248 6633 25276
rect 6512 25236 6518 25248
rect 6621 25245 6633 25248
rect 6667 25245 6679 25279
rect 6621 25239 6679 25245
rect 9490 25236 9496 25288
rect 9548 25236 9554 25288
rect 11422 25236 11428 25288
rect 11480 25236 11486 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 12434 25276 12440 25288
rect 12391 25248 12440 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 12434 25236 12440 25248
rect 12492 25236 12498 25288
rect 12612 25279 12670 25285
rect 12612 25245 12624 25279
rect 12658 25276 12670 25279
rect 12894 25276 12900 25288
rect 12658 25248 12900 25276
rect 12658 25245 12670 25248
rect 12612 25239 12670 25245
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 8297 25211 8355 25217
rect 8297 25177 8309 25211
rect 8343 25208 8355 25211
rect 8570 25208 8576 25220
rect 8343 25180 8576 25208
rect 8343 25177 8355 25180
rect 8297 25171 8355 25177
rect 8570 25168 8576 25180
rect 8628 25208 8634 25220
rect 15028 25217 15056 25384
rect 15746 25304 15752 25356
rect 15804 25304 15810 25356
rect 16482 25344 16488 25356
rect 16316 25316 16488 25344
rect 15657 25279 15715 25285
rect 15657 25245 15669 25279
rect 15703 25276 15715 25279
rect 16114 25276 16120 25288
rect 15703 25248 16120 25276
rect 15703 25245 15715 25248
rect 15657 25239 15715 25245
rect 16114 25236 16120 25248
rect 16172 25276 16178 25288
rect 16316 25276 16344 25316
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 16592 25353 16620 25384
rect 17512 25384 17592 25412
rect 16577 25347 16635 25353
rect 16577 25313 16589 25347
rect 16623 25313 16635 25347
rect 16577 25307 16635 25313
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 16853 25347 16911 25353
rect 16853 25344 16865 25347
rect 16816 25316 16865 25344
rect 16816 25304 16822 25316
rect 16853 25313 16865 25316
rect 16899 25313 16911 25347
rect 16853 25307 16911 25313
rect 17512 25285 17540 25384
rect 17586 25372 17592 25384
rect 17644 25372 17650 25424
rect 18969 25415 19027 25421
rect 18969 25381 18981 25415
rect 19015 25412 19027 25415
rect 19015 25384 19840 25412
rect 19015 25381 19027 25384
rect 18969 25375 19027 25381
rect 19812 25353 19840 25384
rect 27706 25372 27712 25424
rect 27764 25412 27770 25424
rect 28460 25412 28488 25452
rect 27764 25384 28488 25412
rect 28629 25415 28687 25421
rect 27764 25372 27770 25384
rect 28629 25381 28641 25415
rect 28675 25412 28687 25415
rect 28994 25412 29000 25424
rect 28675 25384 29000 25412
rect 28675 25381 28687 25384
rect 28629 25375 28687 25381
rect 28994 25372 29000 25384
rect 29052 25372 29058 25424
rect 29196 25353 29224 25452
rect 29914 25440 29920 25492
rect 29972 25480 29978 25492
rect 30374 25480 30380 25492
rect 29972 25452 30380 25480
rect 29972 25440 29978 25452
rect 30374 25440 30380 25452
rect 30432 25440 30438 25492
rect 31662 25440 31668 25492
rect 31720 25440 31726 25492
rect 45830 25440 45836 25492
rect 45888 25480 45894 25492
rect 46842 25480 46848 25492
rect 45888 25452 46848 25480
rect 45888 25440 45894 25452
rect 46842 25440 46848 25452
rect 46900 25440 46906 25492
rect 46934 25440 46940 25492
rect 46992 25480 46998 25492
rect 48225 25483 48283 25489
rect 48225 25480 48237 25483
rect 46992 25452 48237 25480
rect 46992 25440 46998 25452
rect 48225 25449 48237 25452
rect 48271 25449 48283 25483
rect 48225 25443 48283 25449
rect 49878 25440 49884 25492
rect 49936 25440 49942 25492
rect 50341 25483 50399 25489
rect 50341 25449 50353 25483
rect 50387 25480 50399 25483
rect 50798 25480 50804 25492
rect 50387 25452 50804 25480
rect 50387 25449 50399 25452
rect 50341 25443 50399 25449
rect 50798 25440 50804 25452
rect 50856 25440 50862 25492
rect 50890 25440 50896 25492
rect 50948 25480 50954 25492
rect 54021 25483 54079 25489
rect 50948 25452 52868 25480
rect 50948 25440 50954 25452
rect 46014 25412 46020 25424
rect 45664 25384 46020 25412
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25313 19855 25347
rect 28353 25347 28411 25353
rect 28353 25344 28365 25347
rect 19797 25307 19855 25313
rect 27264 25316 28365 25344
rect 16172 25248 16344 25276
rect 16393 25279 16451 25285
rect 16172 25236 16178 25248
rect 16393 25245 16405 25279
rect 16439 25276 16451 25279
rect 17497 25279 17555 25285
rect 17497 25276 17509 25279
rect 16439 25248 17509 25276
rect 16439 25245 16451 25248
rect 16393 25239 16451 25245
rect 17497 25245 17509 25248
rect 17543 25245 17555 25279
rect 17497 25239 17555 25245
rect 17589 25279 17647 25285
rect 17589 25245 17601 25279
rect 17635 25276 17647 25279
rect 18782 25276 18788 25288
rect 17635 25248 18788 25276
rect 17635 25245 17647 25248
rect 17589 25239 17647 25245
rect 18782 25236 18788 25248
rect 18840 25236 18846 25288
rect 26234 25236 26240 25288
rect 26292 25236 26298 25288
rect 8941 25211 8999 25217
rect 8941 25208 8953 25211
rect 8628 25180 8953 25208
rect 8628 25168 8634 25180
rect 8941 25177 8953 25180
rect 8987 25177 8999 25211
rect 8941 25171 8999 25177
rect 10965 25211 11023 25217
rect 10965 25177 10977 25211
rect 11011 25208 11023 25211
rect 12069 25211 12127 25217
rect 12069 25208 12081 25211
rect 11011 25180 12081 25208
rect 11011 25177 11023 25180
rect 10965 25171 11023 25177
rect 12069 25177 12081 25180
rect 12115 25177 12127 25211
rect 15013 25211 15071 25217
rect 15013 25208 15025 25211
rect 12069 25171 12127 25177
rect 13924 25180 15025 25208
rect 4890 25100 4896 25152
rect 4948 25100 4954 25152
rect 7098 25100 7104 25152
rect 7156 25140 7162 25152
rect 8389 25143 8447 25149
rect 8389 25140 8401 25143
rect 7156 25112 8401 25140
rect 7156 25100 7162 25112
rect 8389 25109 8401 25112
rect 8435 25109 8447 25143
rect 8389 25103 8447 25109
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11698 25140 11704 25152
rect 11103 25112 11704 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11698 25100 11704 25112
rect 11756 25100 11762 25152
rect 12084 25140 12112 25171
rect 13924 25152 13952 25180
rect 15013 25177 15025 25180
rect 15059 25177 15071 25211
rect 15013 25171 15071 25177
rect 15565 25211 15623 25217
rect 15565 25177 15577 25211
rect 15611 25208 15623 25211
rect 17402 25208 17408 25220
rect 15611 25180 17408 25208
rect 15611 25177 15623 25180
rect 15565 25171 15623 25177
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 17856 25211 17914 25217
rect 17856 25177 17868 25211
rect 17902 25208 17914 25211
rect 18230 25208 18236 25220
rect 17902 25180 18236 25208
rect 17902 25177 17914 25180
rect 17856 25171 17914 25177
rect 18230 25168 18236 25180
rect 18288 25168 18294 25220
rect 27264 25152 27292 25316
rect 28353 25313 28365 25316
rect 28399 25313 28411 25347
rect 28353 25307 28411 25313
rect 29181 25347 29239 25353
rect 29181 25313 29193 25347
rect 29227 25313 29239 25347
rect 29181 25307 29239 25313
rect 31573 25347 31631 25353
rect 31573 25313 31585 25347
rect 31619 25344 31631 25347
rect 38378 25344 38384 25356
rect 31619 25316 38384 25344
rect 31619 25313 31631 25316
rect 31573 25307 31631 25313
rect 38378 25304 38384 25316
rect 38436 25304 38442 25356
rect 44821 25347 44879 25353
rect 44821 25313 44833 25347
rect 44867 25344 44879 25347
rect 44910 25344 44916 25356
rect 44867 25316 44916 25344
rect 44867 25313 44879 25316
rect 44821 25307 44879 25313
rect 44910 25304 44916 25316
rect 44968 25344 44974 25356
rect 45664 25353 45692 25384
rect 46014 25372 46020 25384
rect 46072 25372 46078 25424
rect 47305 25415 47363 25421
rect 47305 25381 47317 25415
rect 47351 25412 47363 25415
rect 47351 25384 48728 25412
rect 47351 25381 47363 25384
rect 47305 25375 47363 25381
rect 45649 25347 45707 25353
rect 45649 25344 45661 25347
rect 44968 25316 45661 25344
rect 44968 25304 44974 25316
rect 45649 25313 45661 25316
rect 45695 25313 45707 25347
rect 45649 25307 45707 25313
rect 45922 25304 45928 25356
rect 45980 25344 45986 25356
rect 47029 25347 47087 25353
rect 47029 25344 47041 25347
rect 45980 25316 47041 25344
rect 45980 25304 45986 25316
rect 47029 25313 47041 25316
rect 47075 25313 47087 25347
rect 47029 25307 47087 25313
rect 47578 25304 47584 25356
rect 47636 25304 47642 25356
rect 47765 25347 47823 25353
rect 47765 25313 47777 25347
rect 47811 25344 47823 25347
rect 48222 25344 48228 25356
rect 47811 25316 48228 25344
rect 47811 25313 47823 25316
rect 47765 25307 47823 25313
rect 48222 25304 48228 25316
rect 48280 25304 48286 25356
rect 30190 25276 30196 25288
rect 28920 25248 30196 25276
rect 28169 25211 28227 25217
rect 28169 25177 28181 25211
rect 28215 25208 28227 25211
rect 28920 25208 28948 25248
rect 30190 25236 30196 25248
rect 30248 25236 30254 25288
rect 31317 25279 31375 25285
rect 31317 25245 31329 25279
rect 31363 25276 31375 25279
rect 32122 25276 32128 25288
rect 31363 25248 32128 25276
rect 31363 25245 31375 25248
rect 31317 25239 31375 25245
rect 32122 25236 32128 25248
rect 32180 25236 32186 25288
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25245 32275 25279
rect 32217 25239 32275 25245
rect 45373 25279 45431 25285
rect 45373 25245 45385 25279
rect 45419 25276 45431 25279
rect 45940 25276 45968 25304
rect 45419 25248 45968 25276
rect 45419 25245 45431 25248
rect 45373 25239 45431 25245
rect 28215 25180 28948 25208
rect 28997 25211 29055 25217
rect 28215 25177 28227 25180
rect 28169 25171 28227 25177
rect 28997 25177 29009 25211
rect 29043 25208 29055 25211
rect 29546 25208 29552 25220
rect 29043 25180 29552 25208
rect 29043 25177 29055 25180
rect 28997 25171 29055 25177
rect 29546 25168 29552 25180
rect 29604 25168 29610 25220
rect 32232 25208 32260 25239
rect 46750 25236 46756 25288
rect 46808 25236 46814 25288
rect 46842 25236 46848 25288
rect 46900 25285 46906 25288
rect 46900 25279 46949 25285
rect 46900 25245 46903 25279
rect 46937 25245 46949 25279
rect 47596 25276 47624 25304
rect 47949 25279 48007 25285
rect 47949 25276 47961 25279
rect 47596 25248 47961 25276
rect 46900 25239 46949 25245
rect 47949 25245 47961 25248
rect 47995 25245 48007 25279
rect 47949 25239 48007 25245
rect 46900 25236 46906 25239
rect 30208 25180 32260 25208
rect 45465 25211 45523 25217
rect 12618 25140 12624 25152
rect 12084 25112 12624 25140
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 13906 25100 13912 25152
rect 13964 25100 13970 25152
rect 14734 25100 14740 25152
rect 14792 25100 14798 25152
rect 16022 25100 16028 25152
rect 16080 25100 16086 25152
rect 25130 25100 25136 25152
rect 25188 25100 25194 25152
rect 25590 25100 25596 25152
rect 25648 25100 25654 25152
rect 27246 25100 27252 25152
rect 27304 25100 27310 25152
rect 28261 25143 28319 25149
rect 28261 25109 28273 25143
rect 28307 25140 28319 25143
rect 29086 25140 29092 25152
rect 28307 25112 29092 25140
rect 28307 25109 28319 25112
rect 28261 25103 28319 25109
rect 29086 25100 29092 25112
rect 29144 25100 29150 25152
rect 30208 25149 30236 25180
rect 45465 25177 45477 25211
rect 45511 25208 45523 25211
rect 45646 25208 45652 25220
rect 45511 25180 45652 25208
rect 45511 25177 45523 25180
rect 45465 25171 45523 25177
rect 45646 25168 45652 25180
rect 45704 25168 45710 25220
rect 30193 25143 30251 25149
rect 30193 25109 30205 25143
rect 30239 25109 30251 25143
rect 30193 25103 30251 25109
rect 45002 25100 45008 25152
rect 45060 25100 45066 25152
rect 46109 25143 46167 25149
rect 46109 25109 46121 25143
rect 46155 25140 46167 25143
rect 48038 25140 48044 25152
rect 46155 25112 48044 25140
rect 46155 25109 46167 25112
rect 46109 25103 46167 25109
rect 48038 25100 48044 25112
rect 48096 25100 48102 25152
rect 48700 25149 48728 25384
rect 49896 25344 49924 25440
rect 50893 25347 50951 25353
rect 50893 25344 50905 25347
rect 49896 25316 50905 25344
rect 50893 25313 50905 25316
rect 50939 25313 50951 25347
rect 52086 25344 52092 25356
rect 50893 25307 50951 25313
rect 51460 25316 52092 25344
rect 50709 25279 50767 25285
rect 50709 25245 50721 25279
rect 50755 25276 50767 25279
rect 51460 25276 51488 25316
rect 52086 25304 52092 25316
rect 52144 25353 52150 25356
rect 52144 25347 52193 25353
rect 52144 25313 52147 25347
rect 52181 25313 52193 25347
rect 52144 25307 52193 25313
rect 52144 25304 52150 25307
rect 52270 25304 52276 25356
rect 52328 25304 52334 25356
rect 52546 25304 52552 25356
rect 52604 25304 52610 25356
rect 50755 25248 51488 25276
rect 50755 25245 50767 25248
rect 50709 25239 50767 25245
rect 51994 25236 52000 25288
rect 52052 25236 52058 25288
rect 52840 25276 52868 25452
rect 54021 25449 54033 25483
rect 54067 25480 54079 25483
rect 54202 25480 54208 25492
rect 54067 25452 54208 25480
rect 54067 25449 54079 25452
rect 54021 25443 54079 25449
rect 54202 25440 54208 25452
rect 54260 25440 54266 25492
rect 54570 25412 54576 25424
rect 53024 25384 54576 25412
rect 53024 25353 53052 25384
rect 54570 25372 54576 25384
rect 54628 25372 54634 25424
rect 53009 25347 53067 25353
rect 53009 25313 53021 25347
rect 53055 25313 53067 25347
rect 53009 25307 53067 25313
rect 53374 25304 53380 25356
rect 53432 25304 53438 25356
rect 54662 25304 54668 25356
rect 54720 25304 54726 25356
rect 53193 25279 53251 25285
rect 52840 25248 53052 25276
rect 53024 25208 53052 25248
rect 53193 25245 53205 25279
rect 53239 25276 53251 25279
rect 53239 25248 53604 25276
rect 53239 25245 53251 25248
rect 53193 25239 53251 25245
rect 53576 25217 53604 25248
rect 53561 25211 53619 25217
rect 53024 25180 53328 25208
rect 48685 25143 48743 25149
rect 48685 25109 48697 25143
rect 48731 25140 48743 25143
rect 48774 25140 48780 25152
rect 48731 25112 48780 25140
rect 48731 25109 48743 25112
rect 48685 25103 48743 25109
rect 48774 25100 48780 25112
rect 48832 25100 48838 25152
rect 50798 25100 50804 25152
rect 50856 25100 50862 25152
rect 51353 25143 51411 25149
rect 51353 25109 51365 25143
rect 51399 25140 51411 25143
rect 53190 25140 53196 25152
rect 51399 25112 53196 25140
rect 51399 25109 51411 25112
rect 51353 25103 51411 25109
rect 53190 25100 53196 25112
rect 53248 25100 53254 25152
rect 53300 25140 53328 25180
rect 53561 25177 53573 25211
rect 53607 25208 53619 25211
rect 54113 25211 54171 25217
rect 54113 25208 54125 25211
rect 53607 25180 54125 25208
rect 53607 25177 53619 25180
rect 53561 25171 53619 25177
rect 54113 25177 54125 25180
rect 54159 25177 54171 25211
rect 54113 25171 54171 25177
rect 53653 25143 53711 25149
rect 53653 25140 53665 25143
rect 53300 25112 53665 25140
rect 53653 25109 53665 25112
rect 53699 25109 53711 25143
rect 53653 25103 53711 25109
rect 1104 25050 59040 25072
rect 1104 24998 15394 25050
rect 15446 24998 15458 25050
rect 15510 24998 15522 25050
rect 15574 24998 15586 25050
rect 15638 24998 15650 25050
rect 15702 24998 29838 25050
rect 29890 24998 29902 25050
rect 29954 24998 29966 25050
rect 30018 24998 30030 25050
rect 30082 24998 30094 25050
rect 30146 24998 44282 25050
rect 44334 24998 44346 25050
rect 44398 24998 44410 25050
rect 44462 24998 44474 25050
rect 44526 24998 44538 25050
rect 44590 24998 58726 25050
rect 58778 24998 58790 25050
rect 58842 24998 58854 25050
rect 58906 24998 58918 25050
rect 58970 24998 58982 25050
rect 59034 24998 59040 25050
rect 1104 24976 59040 24998
rect 5445 24939 5503 24945
rect 5445 24905 5457 24939
rect 5491 24905 5503 24939
rect 5445 24899 5503 24905
rect 6733 24939 6791 24945
rect 6733 24905 6745 24939
rect 6779 24936 6791 24939
rect 7006 24936 7012 24948
rect 6779 24908 7012 24936
rect 6779 24905 6791 24908
rect 6733 24899 6791 24905
rect 4332 24871 4390 24877
rect 4332 24837 4344 24871
rect 4378 24868 4390 24871
rect 4890 24868 4896 24880
rect 4378 24840 4896 24868
rect 4378 24837 4390 24840
rect 4332 24831 4390 24837
rect 4890 24828 4896 24840
rect 4948 24828 4954 24880
rect 5460 24800 5488 24899
rect 7006 24896 7012 24908
rect 7064 24896 7070 24948
rect 7098 24896 7104 24948
rect 7156 24896 7162 24948
rect 7190 24896 7196 24948
rect 7248 24896 7254 24948
rect 8941 24939 8999 24945
rect 8941 24905 8953 24939
rect 8987 24936 8999 24939
rect 9490 24936 9496 24948
rect 8987 24908 9496 24936
rect 8987 24905 8999 24908
rect 8941 24899 8999 24905
rect 9490 24896 9496 24908
rect 9548 24896 9554 24948
rect 11241 24939 11299 24945
rect 11241 24905 11253 24939
rect 11287 24936 11299 24939
rect 11422 24936 11428 24948
rect 11287 24908 11428 24936
rect 11287 24905 11299 24908
rect 11241 24899 11299 24905
rect 11422 24896 11428 24908
rect 11480 24896 11486 24948
rect 11992 24908 13584 24936
rect 5537 24803 5595 24809
rect 5537 24800 5549 24803
rect 5460 24772 5549 24800
rect 5537 24769 5549 24772
rect 5583 24769 5595 24803
rect 5537 24763 5595 24769
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 7116 24800 7144 24896
rect 7828 24871 7886 24877
rect 7828 24837 7840 24871
rect 7874 24868 7886 24871
rect 7926 24868 7932 24880
rect 7874 24840 7932 24868
rect 7874 24837 7886 24840
rect 7828 24831 7886 24837
rect 7926 24828 7932 24840
rect 7984 24828 7990 24880
rect 10128 24871 10186 24877
rect 10128 24837 10140 24871
rect 10174 24868 10186 24871
rect 10410 24868 10416 24880
rect 10174 24840 10416 24868
rect 10174 24837 10186 24840
rect 10128 24831 10186 24837
rect 10410 24828 10416 24840
rect 10468 24828 10474 24880
rect 11992 24800 12020 24908
rect 13556 24800 13584 24908
rect 13814 24896 13820 24948
rect 13872 24896 13878 24948
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 14734 24936 14740 24948
rect 14323 24908 14740 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 14292 24868 14320 24899
rect 14734 24896 14740 24908
rect 14792 24896 14798 24948
rect 17313 24939 17371 24945
rect 17313 24905 17325 24939
rect 17359 24936 17371 24939
rect 17402 24936 17408 24948
rect 17359 24908 17408 24936
rect 17359 24905 17371 24908
rect 17313 24899 17371 24905
rect 17402 24896 17408 24908
rect 17460 24896 17466 24948
rect 18230 24896 18236 24948
rect 18288 24896 18294 24948
rect 29546 24896 29552 24948
rect 29604 24936 29610 24948
rect 29825 24939 29883 24945
rect 29825 24936 29837 24939
rect 29604 24908 29837 24936
rect 29604 24896 29610 24908
rect 29825 24905 29837 24908
rect 29871 24905 29883 24939
rect 29825 24899 29883 24905
rect 30653 24939 30711 24945
rect 30653 24905 30665 24939
rect 30699 24936 30711 24939
rect 30834 24936 30840 24948
rect 30699 24908 30840 24936
rect 30699 24905 30711 24908
rect 30653 24899 30711 24905
rect 30834 24896 30840 24908
rect 30892 24896 30898 24948
rect 43257 24939 43315 24945
rect 43257 24905 43269 24939
rect 43303 24905 43315 24939
rect 43257 24899 43315 24905
rect 14108 24840 14320 24868
rect 5960 24772 7144 24800
rect 7392 24772 8708 24800
rect 5960 24760 5966 24772
rect 7392 24741 7420 24772
rect 8680 24744 8708 24772
rect 9232 24772 12020 24800
rect 13464 24772 13584 24800
rect 13725 24803 13783 24809
rect 4065 24735 4123 24741
rect 4065 24732 4077 24735
rect 3988 24704 4077 24732
rect 3988 24608 4016 24704
rect 4065 24701 4077 24704
rect 4111 24701 4123 24735
rect 4065 24695 4123 24701
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24701 7435 24735
rect 7377 24695 7435 24701
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24701 7619 24735
rect 7561 24695 7619 24701
rect 6362 24664 6368 24676
rect 5368 24636 6368 24664
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 5368 24596 5396 24636
rect 6362 24624 6368 24636
rect 6420 24664 6426 24676
rect 7576 24664 7604 24695
rect 8662 24692 8668 24744
rect 8720 24732 8726 24744
rect 9232 24741 9260 24772
rect 9217 24735 9275 24741
rect 9217 24732 9229 24735
rect 8720 24704 9229 24732
rect 8720 24692 8726 24704
rect 9217 24701 9229 24704
rect 9263 24701 9275 24735
rect 9217 24695 9275 24701
rect 9858 24692 9864 24744
rect 9916 24692 9922 24744
rect 12526 24692 12532 24744
rect 12584 24692 12590 24744
rect 12618 24692 12624 24744
rect 12676 24741 12682 24744
rect 12676 24735 12725 24741
rect 12676 24701 12679 24735
rect 12713 24701 12725 24735
rect 12676 24695 12725 24701
rect 12805 24735 12863 24741
rect 12805 24701 12817 24735
rect 12851 24732 12863 24735
rect 12851 24704 13032 24732
rect 12851 24701 12863 24704
rect 12805 24695 12863 24701
rect 12676 24692 12682 24695
rect 6420 24636 7604 24664
rect 6420 24624 6426 24636
rect 4028 24568 5396 24596
rect 4028 24556 4034 24568
rect 6178 24556 6184 24608
rect 6236 24556 6242 24608
rect 7576 24596 7604 24636
rect 9876 24596 9904 24692
rect 7576 24568 9904 24596
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 11701 24599 11759 24605
rect 11701 24596 11713 24599
rect 11296 24568 11713 24596
rect 11296 24556 11302 24568
rect 11701 24565 11713 24568
rect 11747 24565 11759 24599
rect 11701 24559 11759 24565
rect 11882 24556 11888 24608
rect 11940 24556 11946 24608
rect 12342 24556 12348 24608
rect 12400 24596 12406 24608
rect 13004 24596 13032 24704
rect 13081 24667 13139 24673
rect 13081 24633 13093 24667
rect 13127 24664 13139 24667
rect 13170 24664 13176 24676
rect 13127 24636 13176 24664
rect 13127 24633 13139 24636
rect 13081 24627 13139 24633
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 13464 24664 13492 24772
rect 13725 24769 13737 24803
rect 13771 24800 13783 24803
rect 14108 24800 14136 24840
rect 17862 24828 17868 24880
rect 17920 24868 17926 24880
rect 19794 24868 19800 24880
rect 17920 24840 19800 24868
rect 17920 24828 17926 24840
rect 19794 24828 19800 24840
rect 19852 24828 19858 24880
rect 27706 24868 27712 24880
rect 26160 24840 27712 24868
rect 13771 24772 14136 24800
rect 14185 24803 14243 24809
rect 13771 24769 13783 24772
rect 13725 24763 13783 24769
rect 14185 24769 14197 24803
rect 14231 24769 14243 24803
rect 14185 24763 14243 24769
rect 13538 24692 13544 24744
rect 13596 24692 13602 24744
rect 13630 24692 13636 24744
rect 13688 24732 13694 24744
rect 14200 24732 14228 24763
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14332 24772 15025 24800
rect 14332 24760 14338 24772
rect 15013 24769 15025 24772
rect 15059 24800 15071 24803
rect 15746 24800 15752 24812
rect 15059 24772 15752 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 15838 24760 15844 24812
rect 15896 24760 15902 24812
rect 16022 24760 16028 24812
rect 16080 24800 16086 24812
rect 16393 24803 16451 24809
rect 16393 24800 16405 24803
rect 16080 24772 16405 24800
rect 16080 24760 16086 24772
rect 16393 24769 16405 24772
rect 16439 24769 16451 24803
rect 16393 24763 16451 24769
rect 16574 24760 16580 24812
rect 16632 24800 16638 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16632 24772 16681 24800
rect 16632 24760 16638 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 18598 24760 18604 24812
rect 18656 24800 18662 24812
rect 18785 24803 18843 24809
rect 18785 24800 18797 24803
rect 18656 24772 18797 24800
rect 18656 24760 18662 24772
rect 18785 24769 18797 24772
rect 18831 24769 18843 24803
rect 18785 24763 18843 24769
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 24029 24803 24087 24809
rect 24029 24800 24041 24803
rect 19392 24772 24041 24800
rect 19392 24760 19398 24772
rect 24029 24769 24041 24772
rect 24075 24800 24087 24803
rect 25314 24800 25320 24812
rect 24075 24772 25320 24800
rect 24075 24769 24087 24772
rect 24029 24763 24087 24769
rect 25314 24760 25320 24772
rect 25372 24800 25378 24812
rect 26160 24800 26188 24840
rect 27706 24828 27712 24840
rect 27764 24828 27770 24880
rect 29086 24828 29092 24880
rect 29144 24868 29150 24880
rect 29730 24868 29736 24880
rect 29144 24840 29736 24868
rect 29144 24828 29150 24840
rect 29730 24828 29736 24840
rect 29788 24868 29794 24880
rect 30561 24871 30619 24877
rect 30561 24868 30573 24871
rect 29788 24840 30573 24868
rect 29788 24828 29794 24840
rect 30561 24837 30573 24840
rect 30607 24837 30619 24871
rect 30561 24831 30619 24837
rect 25372 24772 26188 24800
rect 26257 24803 26315 24809
rect 25372 24760 25378 24772
rect 26257 24769 26269 24803
rect 26303 24800 26315 24803
rect 26303 24772 26464 24800
rect 26303 24769 26315 24772
rect 26257 24763 26315 24769
rect 13688 24704 14228 24732
rect 14369 24735 14427 24741
rect 13688 24692 13694 24704
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 15764 24732 15792 24760
rect 20073 24735 20131 24741
rect 20073 24732 20085 24735
rect 15764 24704 20085 24732
rect 14369 24695 14427 24701
rect 20073 24701 20085 24704
rect 20119 24732 20131 24735
rect 20806 24732 20812 24744
rect 20119 24704 20812 24732
rect 20119 24701 20131 24704
rect 20073 24695 20131 24701
rect 14384 24664 14412 24695
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 24210 24692 24216 24744
rect 24268 24692 24274 24744
rect 26436 24732 26464 24772
rect 26510 24760 26516 24812
rect 26568 24800 26574 24812
rect 27614 24800 27620 24812
rect 26568 24772 27620 24800
rect 26568 24760 26574 24772
rect 27614 24760 27620 24772
rect 27672 24760 27678 24812
rect 28442 24760 28448 24812
rect 28500 24760 28506 24812
rect 28994 24760 29000 24812
rect 29052 24760 29058 24812
rect 29270 24760 29276 24812
rect 29328 24760 29334 24812
rect 42702 24760 42708 24812
rect 42760 24800 42766 24812
rect 42760 24772 42840 24800
rect 42760 24760 42766 24772
rect 26973 24735 27031 24741
rect 26973 24732 26985 24735
rect 26436 24704 26985 24732
rect 26973 24701 26985 24704
rect 27019 24701 27031 24735
rect 26973 24695 27031 24701
rect 27525 24735 27583 24741
rect 27525 24701 27537 24735
rect 27571 24732 27583 24735
rect 27982 24732 27988 24744
rect 27571 24704 27988 24732
rect 27571 24701 27583 24704
rect 27525 24695 27583 24701
rect 27982 24692 27988 24704
rect 28040 24692 28046 24744
rect 30834 24692 30840 24744
rect 30892 24732 30898 24744
rect 42812 24741 42840 24772
rect 42886 24760 42892 24812
rect 42944 24760 42950 24812
rect 43272 24800 43300 24899
rect 45922 24896 45928 24948
rect 45980 24896 45986 24948
rect 51166 24896 51172 24948
rect 51224 24936 51230 24948
rect 51994 24936 52000 24948
rect 51224 24908 52000 24936
rect 51224 24896 51230 24908
rect 51994 24896 52000 24908
rect 52052 24896 52058 24948
rect 52546 24896 52552 24948
rect 52604 24896 52610 24948
rect 53193 24939 53251 24945
rect 53193 24905 53205 24939
rect 53239 24936 53251 24939
rect 53374 24936 53380 24948
rect 53239 24908 53380 24936
rect 53239 24905 53251 24908
rect 53193 24899 53251 24905
rect 52564 24868 52592 24896
rect 50632 24840 52592 24868
rect 50632 24812 50660 24840
rect 43901 24803 43959 24809
rect 43901 24800 43913 24803
rect 43272 24772 43913 24800
rect 43901 24769 43913 24772
rect 43947 24769 43959 24803
rect 43901 24763 43959 24769
rect 45002 24760 45008 24812
rect 45060 24800 45066 24812
rect 45189 24803 45247 24809
rect 45189 24800 45201 24803
rect 45060 24772 45201 24800
rect 45060 24760 45066 24772
rect 45189 24769 45201 24772
rect 45235 24769 45247 24803
rect 45189 24763 45247 24769
rect 45370 24760 45376 24812
rect 45428 24800 45434 24812
rect 45833 24803 45891 24809
rect 45833 24800 45845 24803
rect 45428 24772 45845 24800
rect 45428 24760 45434 24772
rect 45833 24769 45845 24772
rect 45879 24769 45891 24803
rect 45833 24763 45891 24769
rect 46382 24760 46388 24812
rect 46440 24800 46446 24812
rect 46477 24803 46535 24809
rect 46477 24800 46489 24803
rect 46440 24772 46489 24800
rect 46440 24760 46446 24772
rect 46477 24769 46489 24772
rect 46523 24769 46535 24803
rect 50341 24803 50399 24809
rect 46477 24763 46535 24769
rect 46584 24772 47992 24800
rect 31205 24735 31263 24741
rect 31205 24732 31217 24735
rect 30892 24704 31217 24732
rect 30892 24692 30898 24704
rect 31205 24701 31217 24704
rect 31251 24701 31263 24735
rect 31205 24695 31263 24701
rect 42613 24735 42671 24741
rect 42613 24701 42625 24735
rect 42659 24701 42671 24735
rect 42613 24695 42671 24701
rect 42797 24735 42855 24741
rect 42797 24701 42809 24735
rect 42843 24732 42855 24735
rect 44085 24735 44143 24741
rect 44085 24732 44097 24735
rect 42843 24704 44097 24732
rect 42843 24701 42855 24704
rect 42797 24695 42855 24701
rect 44085 24701 44097 24704
rect 44131 24701 44143 24735
rect 44085 24695 44143 24701
rect 15381 24667 15439 24673
rect 15381 24664 15393 24667
rect 13464 24636 15393 24664
rect 15381 24633 15393 24636
rect 15427 24664 15439 24667
rect 16206 24664 16212 24676
rect 15427 24636 16212 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 24765 24667 24823 24673
rect 24765 24633 24777 24667
rect 24811 24664 24823 24667
rect 25222 24664 25228 24676
rect 24811 24636 25228 24664
rect 24811 24633 24823 24636
rect 24765 24627 24823 24633
rect 25222 24624 25228 24636
rect 25280 24624 25286 24676
rect 12400 24568 13032 24596
rect 25133 24599 25191 24605
rect 12400 24556 12406 24568
rect 25133 24565 25145 24599
rect 25179 24596 25191 24599
rect 26234 24596 26240 24608
rect 25179 24568 26240 24596
rect 25179 24565 25191 24568
rect 25133 24559 25191 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 30193 24599 30251 24605
rect 30193 24565 30205 24599
rect 30239 24596 30251 24599
rect 30282 24596 30288 24608
rect 30239 24568 30288 24596
rect 30239 24565 30251 24568
rect 30193 24559 30251 24565
rect 30282 24556 30288 24568
rect 30340 24556 30346 24608
rect 42242 24556 42248 24608
rect 42300 24596 42306 24608
rect 42628 24596 42656 24695
rect 44634 24692 44640 24744
rect 44692 24692 44698 24744
rect 42702 24624 42708 24676
rect 42760 24664 42766 24676
rect 46584 24664 46612 24772
rect 47964 24732 47992 24772
rect 50341 24769 50353 24803
rect 50387 24800 50399 24803
rect 50614 24800 50620 24812
rect 50387 24772 50620 24800
rect 50387 24769 50399 24772
rect 50341 24763 50399 24769
rect 50614 24760 50620 24772
rect 50672 24760 50678 24812
rect 50709 24803 50767 24809
rect 50709 24769 50721 24803
rect 50755 24800 50767 24803
rect 52546 24800 52552 24812
rect 50755 24772 52552 24800
rect 50755 24769 50767 24772
rect 50709 24763 50767 24769
rect 50724 24732 50752 24763
rect 52546 24760 52552 24772
rect 52604 24760 52610 24812
rect 47964 24704 50752 24732
rect 42760 24636 46612 24664
rect 42760 24624 42766 24636
rect 46658 24624 46664 24676
rect 46716 24664 46722 24676
rect 53208 24664 53236 24899
rect 53374 24896 53380 24908
rect 53432 24896 53438 24948
rect 46716 24636 53236 24664
rect 46716 24624 46722 24636
rect 42794 24596 42800 24608
rect 42300 24568 42800 24596
rect 42300 24556 42306 24568
rect 42794 24556 42800 24568
rect 42852 24556 42858 24608
rect 42978 24556 42984 24608
rect 43036 24596 43042 24608
rect 46952 24605 46980 24636
rect 43349 24599 43407 24605
rect 43349 24596 43361 24599
rect 43036 24568 43361 24596
rect 43036 24556 43042 24568
rect 43349 24565 43361 24568
rect 43395 24565 43407 24599
rect 43349 24559 43407 24565
rect 46937 24599 46995 24605
rect 46937 24565 46949 24599
rect 46983 24565 46995 24599
rect 46937 24559 46995 24565
rect 47486 24556 47492 24608
rect 47544 24596 47550 24608
rect 47765 24599 47823 24605
rect 47765 24596 47777 24599
rect 47544 24568 47777 24596
rect 47544 24556 47550 24568
rect 47765 24565 47777 24568
rect 47811 24565 47823 24599
rect 47765 24559 47823 24565
rect 51258 24556 51264 24608
rect 51316 24556 51322 24608
rect 1104 24506 58880 24528
rect 1104 24454 8172 24506
rect 8224 24454 8236 24506
rect 8288 24454 8300 24506
rect 8352 24454 8364 24506
rect 8416 24454 8428 24506
rect 8480 24454 22616 24506
rect 22668 24454 22680 24506
rect 22732 24454 22744 24506
rect 22796 24454 22808 24506
rect 22860 24454 22872 24506
rect 22924 24454 37060 24506
rect 37112 24454 37124 24506
rect 37176 24454 37188 24506
rect 37240 24454 37252 24506
rect 37304 24454 37316 24506
rect 37368 24454 51504 24506
rect 51556 24454 51568 24506
rect 51620 24454 51632 24506
rect 51684 24454 51696 24506
rect 51748 24454 51760 24506
rect 51812 24454 58880 24506
rect 1104 24432 58880 24454
rect 5445 24395 5503 24401
rect 5445 24361 5457 24395
rect 5491 24392 5503 24395
rect 5534 24392 5540 24404
rect 5491 24364 5540 24392
rect 5491 24361 5503 24364
rect 5445 24355 5503 24361
rect 5534 24352 5540 24364
rect 5592 24352 5598 24404
rect 6178 24352 6184 24404
rect 6236 24352 6242 24404
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 7248 24364 7880 24392
rect 7248 24352 7254 24364
rect 3970 24216 3976 24268
rect 4028 24216 4034 24268
rect 5902 24216 5908 24268
rect 5960 24216 5966 24268
rect 6086 24216 6092 24268
rect 6144 24216 6150 24268
rect 6196 24256 6224 24352
rect 7193 24259 7251 24265
rect 7193 24256 7205 24259
rect 6196 24228 7205 24256
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24188 5871 24191
rect 6196 24188 6224 24228
rect 7193 24225 7205 24228
rect 7239 24225 7251 24259
rect 7193 24219 7251 24225
rect 7466 24216 7472 24268
rect 7524 24216 7530 24268
rect 5859 24160 6224 24188
rect 5859 24157 5871 24160
rect 5813 24151 5871 24157
rect 6914 24148 6920 24200
rect 6972 24148 6978 24200
rect 7006 24148 7012 24200
rect 7064 24197 7070 24200
rect 7064 24191 7113 24197
rect 7064 24157 7067 24191
rect 7101 24157 7113 24191
rect 7852 24188 7880 24364
rect 11882 24352 11888 24404
rect 11940 24392 11946 24404
rect 11940 24364 13492 24392
rect 11940 24352 11946 24364
rect 13464 24324 13492 24364
rect 13538 24352 13544 24404
rect 13596 24392 13602 24404
rect 14093 24395 14151 24401
rect 14093 24392 14105 24395
rect 13596 24364 14105 24392
rect 13596 24352 13602 24364
rect 14093 24361 14105 24364
rect 14139 24361 14151 24395
rect 14093 24355 14151 24361
rect 26510 24352 26516 24404
rect 26568 24352 26574 24404
rect 41601 24395 41659 24401
rect 41601 24361 41613 24395
rect 41647 24392 41659 24395
rect 42702 24392 42708 24404
rect 41647 24364 42708 24392
rect 41647 24361 41659 24364
rect 41601 24355 41659 24361
rect 42702 24352 42708 24364
rect 42760 24352 42766 24404
rect 42794 24352 42800 24404
rect 42852 24392 42858 24404
rect 43809 24395 43867 24401
rect 42852 24364 43392 24392
rect 42852 24352 42858 24364
rect 13909 24327 13967 24333
rect 13464 24296 13860 24324
rect 7929 24259 7987 24265
rect 7929 24225 7941 24259
rect 7975 24256 7987 24259
rect 8570 24256 8576 24268
rect 7975 24228 8576 24256
rect 7975 24225 7987 24228
rect 7929 24219 7987 24225
rect 8570 24216 8576 24228
rect 8628 24216 8634 24268
rect 11238 24216 11244 24268
rect 11296 24256 11302 24268
rect 11977 24259 12035 24265
rect 11977 24256 11989 24259
rect 11296 24228 11989 24256
rect 11296 24216 11302 24228
rect 11977 24225 11989 24228
rect 12023 24256 12035 24259
rect 12023 24228 12664 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 8113 24191 8171 24197
rect 8113 24188 8125 24191
rect 7852 24160 8125 24188
rect 7064 24151 7113 24157
rect 8113 24157 8125 24160
rect 8159 24157 8171 24191
rect 8113 24151 8171 24157
rect 7064 24148 7070 24151
rect 9858 24148 9864 24200
rect 9916 24188 9922 24200
rect 9953 24191 10011 24197
rect 9953 24188 9965 24191
rect 9916 24160 9965 24188
rect 9916 24148 9922 24160
rect 9953 24157 9965 24160
rect 9999 24188 10011 24191
rect 12434 24188 12440 24200
rect 9999 24160 12440 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 12434 24148 12440 24160
rect 12492 24188 12498 24200
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12492 24160 12541 24188
rect 12492 24148 12498 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12636 24188 12664 24228
rect 13832 24200 13860 24296
rect 13909 24293 13921 24327
rect 13955 24324 13967 24327
rect 43364 24324 43392 24364
rect 43809 24361 43821 24395
rect 43855 24392 43867 24395
rect 44634 24392 44640 24404
rect 43855 24364 44640 24392
rect 43855 24361 43867 24364
rect 43809 24355 43867 24361
rect 44634 24352 44640 24364
rect 44692 24352 44698 24404
rect 46658 24352 46664 24404
rect 46716 24352 46722 24404
rect 46676 24324 46704 24352
rect 13955 24296 14688 24324
rect 43364 24296 46704 24324
rect 13955 24293 13967 24296
rect 13909 24287 13967 24293
rect 14660 24265 14688 24296
rect 14645 24259 14703 24265
rect 14645 24225 14657 24259
rect 14691 24225 14703 24259
rect 14645 24219 14703 24225
rect 24489 24259 24547 24265
rect 24489 24225 24501 24259
rect 24535 24256 24547 24259
rect 24854 24256 24860 24268
rect 24535 24228 24860 24256
rect 24535 24225 24547 24228
rect 24489 24219 24547 24225
rect 24854 24216 24860 24228
rect 24912 24256 24918 24268
rect 24912 24228 26096 24256
rect 24912 24216 24918 24228
rect 26068 24200 26096 24228
rect 13078 24188 13084 24200
rect 12636 24160 13084 24188
rect 12529 24151 12587 24157
rect 13078 24148 13084 24160
rect 13136 24188 13142 24200
rect 13722 24188 13728 24200
rect 13136 24160 13728 24188
rect 13136 24148 13142 24160
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 13814 24148 13820 24200
rect 13872 24148 13878 24200
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 15381 24191 15439 24197
rect 15381 24188 15393 24191
rect 14148 24160 15393 24188
rect 14148 24148 14154 24160
rect 15381 24157 15393 24160
rect 15427 24157 15439 24191
rect 15381 24151 15439 24157
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 4240 24123 4298 24129
rect 4240 24089 4252 24123
rect 4286 24120 4298 24123
rect 4522 24120 4528 24132
rect 4286 24092 4528 24120
rect 4286 24089 4298 24092
rect 4240 24083 4298 24089
rect 4522 24080 4528 24092
rect 4580 24080 4586 24132
rect 10220 24123 10278 24129
rect 10220 24089 10232 24123
rect 10266 24120 10278 24123
rect 10686 24120 10692 24132
rect 10266 24092 10692 24120
rect 10266 24089 10278 24092
rect 10220 24083 10278 24089
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 11793 24123 11851 24129
rect 11793 24089 11805 24123
rect 11839 24120 11851 24123
rect 12342 24120 12348 24132
rect 11839 24092 12348 24120
rect 11839 24089 11851 24092
rect 11793 24083 11851 24089
rect 12342 24080 12348 24092
rect 12400 24080 12406 24132
rect 12452 24120 12480 24148
rect 12618 24120 12624 24132
rect 12452 24092 12624 24120
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 12796 24123 12854 24129
rect 12796 24089 12808 24123
rect 12842 24120 12854 24123
rect 14829 24123 14887 24129
rect 14829 24120 14841 24123
rect 12842 24092 14841 24120
rect 12842 24089 12854 24092
rect 12796 24083 12854 24089
rect 14829 24089 14841 24092
rect 14875 24089 14887 24123
rect 20088 24120 20116 24151
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 20806 24148 20812 24200
rect 20864 24148 20870 24200
rect 20898 24148 20904 24200
rect 20956 24148 20962 24200
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22244 24160 22661 24188
rect 22244 24148 22250 24160
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 25004 24160 25053 24188
rect 25004 24148 25010 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25130 24148 25136 24200
rect 25188 24188 25194 24200
rect 25225 24191 25283 24197
rect 25225 24188 25237 24191
rect 25188 24160 25237 24188
rect 25188 24148 25194 24160
rect 25225 24157 25237 24160
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 26050 24148 26056 24200
rect 26108 24148 26114 24200
rect 27062 24148 27068 24200
rect 27120 24148 27126 24200
rect 33502 24148 33508 24200
rect 33560 24148 33566 24200
rect 33686 24148 33692 24200
rect 33744 24148 33750 24200
rect 35986 24148 35992 24200
rect 36044 24148 36050 24200
rect 37550 24148 37556 24200
rect 37608 24148 37614 24200
rect 37734 24148 37740 24200
rect 37792 24148 37798 24200
rect 40402 24148 40408 24200
rect 40460 24148 40466 24200
rect 41138 24148 41144 24200
rect 41196 24148 41202 24200
rect 42334 24148 42340 24200
rect 42392 24148 42398 24200
rect 42429 24191 42487 24197
rect 42429 24157 42441 24191
rect 42475 24188 42487 24191
rect 42518 24188 42524 24200
rect 42475 24160 42524 24188
rect 42475 24157 42487 24160
rect 42429 24151 42487 24157
rect 42518 24148 42524 24160
rect 42576 24148 42582 24200
rect 42696 24191 42754 24197
rect 42696 24157 42708 24191
rect 42742 24188 42754 24191
rect 42978 24188 42984 24200
rect 42742 24160 42984 24188
rect 42742 24157 42754 24160
rect 42696 24151 42754 24157
rect 42978 24148 42984 24160
rect 43036 24148 43042 24200
rect 43990 24148 43996 24200
rect 44048 24148 44054 24200
rect 46474 24148 46480 24200
rect 46532 24148 46538 24200
rect 46750 24148 46756 24200
rect 46808 24148 46814 24200
rect 48130 24148 48136 24200
rect 48188 24148 48194 24200
rect 50982 24148 50988 24200
rect 51040 24148 51046 24200
rect 51902 24148 51908 24200
rect 51960 24148 51966 24200
rect 52638 24148 52644 24200
rect 52696 24148 52702 24200
rect 53282 24148 53288 24200
rect 53340 24148 53346 24200
rect 54386 24148 54392 24200
rect 54444 24148 54450 24200
rect 55306 24148 55312 24200
rect 55364 24148 55370 24200
rect 56870 24148 56876 24200
rect 56928 24188 56934 24200
rect 57149 24191 57207 24197
rect 57149 24188 57161 24191
rect 56928 24160 57161 24188
rect 56928 24148 56934 24160
rect 57149 24157 57161 24160
rect 57195 24157 57207 24191
rect 57149 24151 57207 24157
rect 57238 24148 57244 24200
rect 57296 24188 57302 24200
rect 57885 24191 57943 24197
rect 57885 24188 57897 24191
rect 57296 24160 57897 24188
rect 57296 24148 57302 24160
rect 57885 24157 57897 24160
rect 57931 24157 57943 24191
rect 57885 24151 57943 24157
rect 20254 24120 20260 24132
rect 20088 24092 20260 24120
rect 14829 24083 14887 24089
rect 20254 24080 20260 24092
rect 20312 24080 20318 24132
rect 20824 24120 20852 24148
rect 23201 24123 23259 24129
rect 23201 24120 23213 24123
rect 20824 24092 23213 24120
rect 23201 24089 23213 24092
rect 23247 24089 23259 24123
rect 23201 24083 23259 24089
rect 23290 24080 23296 24132
rect 23348 24120 23354 24132
rect 27522 24120 27528 24132
rect 23348 24092 27528 24120
rect 23348 24080 23354 24092
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 47305 24123 47363 24129
rect 47305 24089 47317 24123
rect 47351 24120 47363 24123
rect 47351 24092 48360 24120
rect 47351 24089 47363 24092
rect 47305 24083 47363 24089
rect 48332 24064 48360 24092
rect 5350 24012 5356 24064
rect 5408 24012 5414 24064
rect 6273 24055 6331 24061
rect 6273 24021 6285 24055
rect 6319 24052 6331 24055
rect 7558 24052 7564 24064
rect 6319 24024 7564 24052
rect 6319 24021 6331 24024
rect 6273 24015 6331 24021
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 7650 24012 7656 24064
rect 7708 24052 7714 24064
rect 8389 24055 8447 24061
rect 8389 24052 8401 24055
rect 7708 24024 8401 24052
rect 7708 24012 7714 24024
rect 8389 24021 8401 24024
rect 8435 24021 8447 24055
rect 8389 24015 8447 24021
rect 11330 24012 11336 24064
rect 11388 24012 11394 24064
rect 11422 24012 11428 24064
rect 11480 24012 11486 24064
rect 11698 24012 11704 24064
rect 11756 24052 11762 24064
rect 11885 24055 11943 24061
rect 11885 24052 11897 24055
rect 11756 24024 11897 24052
rect 11756 24012 11762 24024
rect 11885 24021 11897 24024
rect 11931 24052 11943 24055
rect 13630 24052 13636 24064
rect 11931 24024 13636 24052
rect 11931 24021 11943 24024
rect 11885 24015 11943 24021
rect 13630 24012 13636 24024
rect 13688 24012 13694 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 20809 24055 20867 24061
rect 20809 24021 20821 24055
rect 20855 24052 20867 24055
rect 21266 24052 21272 24064
rect 20855 24024 21272 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 21266 24012 21272 24024
rect 21324 24012 21330 24064
rect 21450 24012 21456 24064
rect 21508 24052 21514 24064
rect 21545 24055 21603 24061
rect 21545 24052 21557 24055
rect 21508 24024 21557 24052
rect 21508 24012 21514 24024
rect 21545 24021 21557 24024
rect 21591 24021 21603 24055
rect 21545 24015 21603 24021
rect 22094 24012 22100 24064
rect 22152 24012 22158 24064
rect 23382 24012 23388 24064
rect 23440 24012 23446 24064
rect 25038 24012 25044 24064
rect 25096 24052 25102 24064
rect 26510 24052 26516 24064
rect 25096 24024 26516 24052
rect 25096 24012 25102 24024
rect 26510 24012 26516 24024
rect 26568 24012 26574 24064
rect 27709 24055 27767 24061
rect 27709 24021 27721 24055
rect 27755 24052 27767 24055
rect 27798 24052 27804 24064
rect 27755 24024 27804 24052
rect 27755 24021 27767 24024
rect 27709 24015 27767 24021
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 32950 24012 32956 24064
rect 33008 24012 33014 24064
rect 34330 24012 34336 24064
rect 34388 24012 34394 24064
rect 35434 24012 35440 24064
rect 35492 24012 35498 24064
rect 36814 24012 36820 24064
rect 36872 24052 36878 24064
rect 37001 24055 37059 24061
rect 37001 24052 37013 24055
rect 36872 24024 37013 24052
rect 36872 24012 36878 24024
rect 37001 24021 37013 24024
rect 37047 24021 37059 24055
rect 37001 24015 37059 24021
rect 38381 24055 38439 24061
rect 38381 24021 38393 24055
rect 38427 24052 38439 24055
rect 38930 24052 38936 24064
rect 38427 24024 38936 24052
rect 38427 24021 38439 24024
rect 38381 24015 38439 24021
rect 38930 24012 38936 24024
rect 38988 24012 38994 24064
rect 39666 24012 39672 24064
rect 39724 24012 39730 24064
rect 39850 24012 39856 24064
rect 39908 24012 39914 24064
rect 40586 24012 40592 24064
rect 40644 24012 40650 24064
rect 41690 24012 41696 24064
rect 41748 24012 41754 24064
rect 44634 24012 44640 24064
rect 44692 24012 44698 24064
rect 45922 24012 45928 24064
rect 45980 24012 45986 24064
rect 47394 24012 47400 24064
rect 47452 24052 47458 24064
rect 47489 24055 47547 24061
rect 47489 24052 47501 24055
rect 47452 24024 47501 24052
rect 47452 24012 47458 24024
rect 47489 24021 47501 24024
rect 47535 24021 47547 24055
rect 47489 24015 47547 24021
rect 48314 24012 48320 24064
rect 48372 24012 48378 24064
rect 50430 24012 50436 24064
rect 50488 24012 50494 24064
rect 51261 24055 51319 24061
rect 51261 24021 51273 24055
rect 51307 24052 51319 24055
rect 51350 24052 51356 24064
rect 51307 24024 51356 24052
rect 51307 24021 51319 24024
rect 51261 24015 51319 24021
rect 51350 24012 51356 24024
rect 51408 24012 51414 24064
rect 51997 24055 52055 24061
rect 51997 24021 52009 24055
rect 52043 24052 52055 24055
rect 52454 24052 52460 24064
rect 52043 24024 52460 24052
rect 52043 24021 52055 24024
rect 51997 24015 52055 24021
rect 52454 24012 52460 24024
rect 52512 24012 52518 24064
rect 52730 24012 52736 24064
rect 52788 24012 52794 24064
rect 53650 24012 53656 24064
rect 53708 24012 53714 24064
rect 53834 24012 53840 24064
rect 53892 24012 53898 24064
rect 54570 24012 54576 24064
rect 54628 24052 54634 24064
rect 54757 24055 54815 24061
rect 54757 24052 54769 24055
rect 54628 24024 54769 24052
rect 54628 24012 54634 24024
rect 54757 24021 54769 24024
rect 54803 24021 54815 24055
rect 54757 24015 54815 24021
rect 55214 24012 55220 24064
rect 55272 24052 55278 24064
rect 55953 24055 56011 24061
rect 55953 24052 55965 24055
rect 55272 24024 55965 24052
rect 55272 24012 55278 24024
rect 55953 24021 55965 24024
rect 55999 24052 56011 24055
rect 56042 24052 56048 24064
rect 55999 24024 56048 24052
rect 55999 24021 56011 24024
rect 55953 24015 56011 24021
rect 56042 24012 56048 24024
rect 56100 24012 56106 24064
rect 56594 24012 56600 24064
rect 56652 24012 56658 24064
rect 57330 24012 57336 24064
rect 57388 24012 57394 24064
rect 1104 23962 59040 23984
rect 1104 23910 15394 23962
rect 15446 23910 15458 23962
rect 15510 23910 15522 23962
rect 15574 23910 15586 23962
rect 15638 23910 15650 23962
rect 15702 23910 29838 23962
rect 29890 23910 29902 23962
rect 29954 23910 29966 23962
rect 30018 23910 30030 23962
rect 30082 23910 30094 23962
rect 30146 23910 44282 23962
rect 44334 23910 44346 23962
rect 44398 23910 44410 23962
rect 44462 23910 44474 23962
rect 44526 23910 44538 23962
rect 44590 23910 58726 23962
rect 58778 23910 58790 23962
rect 58842 23910 58854 23962
rect 58906 23910 58918 23962
rect 58970 23910 58982 23962
rect 59034 23910 59040 23962
rect 1104 23888 59040 23910
rect 5169 23851 5227 23857
rect 5169 23817 5181 23851
rect 5215 23848 5227 23851
rect 5534 23848 5540 23860
rect 5215 23820 5540 23848
rect 5215 23817 5227 23820
rect 5169 23811 5227 23817
rect 5534 23808 5540 23820
rect 5592 23848 5598 23860
rect 5902 23848 5908 23860
rect 5592 23820 5908 23848
rect 5592 23808 5598 23820
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 7006 23848 7012 23860
rect 6196 23820 7012 23848
rect 5350 23740 5356 23792
rect 5408 23740 5414 23792
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23681 5135 23715
rect 5368 23712 5396 23740
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 5368 23684 5549 23712
rect 5077 23675 5135 23681
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 5537 23675 5595 23681
rect 5092 23576 5120 23675
rect 5350 23604 5356 23656
rect 5408 23604 5414 23656
rect 6196 23585 6224 23820
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 10686 23808 10692 23860
rect 10744 23808 10750 23860
rect 11422 23808 11428 23860
rect 11480 23808 11486 23860
rect 13538 23808 13544 23860
rect 13596 23848 13602 23860
rect 13725 23851 13783 23857
rect 13725 23848 13737 23851
rect 13596 23820 13737 23848
rect 13596 23808 13602 23820
rect 13725 23817 13737 23820
rect 13771 23817 13783 23851
rect 13725 23811 13783 23817
rect 14090 23808 14096 23860
rect 14148 23808 14154 23860
rect 17954 23808 17960 23860
rect 18012 23848 18018 23860
rect 18601 23851 18659 23857
rect 18601 23848 18613 23851
rect 18012 23820 18613 23848
rect 18012 23808 18018 23820
rect 18601 23817 18613 23820
rect 18647 23848 18659 23851
rect 19334 23848 19340 23860
rect 18647 23820 19340 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 19426 23808 19432 23860
rect 19484 23808 19490 23860
rect 20162 23808 20168 23860
rect 20220 23808 20226 23860
rect 20254 23808 20260 23860
rect 20312 23808 20318 23860
rect 23290 23808 23296 23860
rect 23348 23808 23354 23860
rect 23569 23851 23627 23857
rect 23569 23817 23581 23851
rect 23615 23848 23627 23851
rect 23934 23848 23940 23860
rect 23615 23820 23940 23848
rect 23615 23817 23627 23820
rect 23569 23811 23627 23817
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 25222 23848 25228 23860
rect 24780 23820 25228 23848
rect 11238 23780 11244 23792
rect 6564 23752 11244 23780
rect 6181 23579 6239 23585
rect 6181 23576 6193 23579
rect 5092 23548 6193 23576
rect 6181 23545 6193 23548
rect 6227 23545 6239 23579
rect 6181 23539 6239 23545
rect 4706 23468 4712 23520
rect 4764 23468 4770 23520
rect 6086 23468 6092 23520
rect 6144 23508 6150 23520
rect 6564 23517 6592 23752
rect 11238 23740 11244 23752
rect 11296 23740 11302 23792
rect 11333 23715 11391 23721
rect 11333 23681 11345 23715
rect 11379 23712 11391 23715
rect 11440 23712 11468 23808
rect 11517 23783 11575 23789
rect 11517 23749 11529 23783
rect 11563 23780 11575 23783
rect 14182 23780 14188 23792
rect 11563 23752 14188 23780
rect 11563 23749 11575 23752
rect 11517 23743 11575 23749
rect 14182 23740 14188 23752
rect 14240 23780 14246 23792
rect 14369 23783 14427 23789
rect 14369 23780 14381 23783
rect 14240 23752 14381 23780
rect 14240 23740 14246 23752
rect 14369 23749 14381 23752
rect 14415 23749 14427 23783
rect 14369 23743 14427 23749
rect 19052 23783 19110 23789
rect 19052 23749 19064 23783
rect 19098 23780 19110 23783
rect 19444 23780 19472 23808
rect 21545 23783 21603 23789
rect 21545 23780 21557 23783
rect 19098 23752 19472 23780
rect 20548 23752 21557 23780
rect 19098 23749 19110 23752
rect 19052 23743 19110 23749
rect 11379 23684 11468 23712
rect 11379 23681 11391 23684
rect 11333 23675 11391 23681
rect 13630 23672 13636 23724
rect 13688 23672 13694 23724
rect 18690 23712 18696 23724
rect 15120 23684 18696 23712
rect 13262 23604 13268 23656
rect 13320 23644 13326 23656
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 13320 23616 13461 23644
rect 13320 23604 13326 23616
rect 13449 23613 13461 23616
rect 13495 23644 13507 23647
rect 15120 23644 15148 23684
rect 18690 23672 18696 23684
rect 18748 23712 18754 23724
rect 20548 23712 20576 23752
rect 21545 23749 21557 23752
rect 21591 23749 21603 23783
rect 21545 23743 21603 23749
rect 18748 23684 20576 23712
rect 20625 23715 20683 23721
rect 18748 23672 18754 23684
rect 20625 23681 20637 23715
rect 20671 23712 20683 23715
rect 21266 23712 21272 23724
rect 20671 23684 21272 23712
rect 20671 23681 20683 23684
rect 20625 23675 20683 23681
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 21560 23712 21588 23743
rect 22094 23740 22100 23792
rect 22152 23780 22158 23792
rect 22189 23783 22247 23789
rect 22189 23780 22201 23783
rect 22152 23752 22201 23780
rect 22152 23740 22158 23752
rect 22189 23749 22201 23752
rect 22235 23749 22247 23783
rect 22189 23743 22247 23749
rect 23308 23712 23336 23808
rect 24780 23780 24808 23820
rect 25222 23808 25228 23820
rect 25280 23848 25286 23860
rect 26789 23851 26847 23857
rect 25280 23820 25912 23848
rect 25280 23808 25286 23820
rect 25884 23792 25912 23820
rect 26789 23817 26801 23851
rect 26835 23848 26847 23851
rect 27062 23848 27068 23860
rect 26835 23820 27068 23848
rect 26835 23817 26847 23820
rect 26789 23811 26847 23817
rect 27062 23808 27068 23820
rect 27120 23808 27126 23860
rect 27522 23808 27528 23860
rect 27580 23848 27586 23860
rect 31294 23848 31300 23860
rect 27580 23820 31300 23848
rect 27580 23808 27586 23820
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 31570 23808 31576 23860
rect 31628 23808 31634 23860
rect 33134 23848 33140 23860
rect 32048 23820 33140 23848
rect 23952 23752 24808 23780
rect 23952 23721 23980 23752
rect 24854 23740 24860 23792
rect 24912 23740 24918 23792
rect 25314 23780 25320 23792
rect 24964 23752 25320 23780
rect 21560 23684 23336 23712
rect 23937 23715 23995 23721
rect 13495 23616 15148 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 15194 23604 15200 23656
rect 15252 23644 15258 23656
rect 15381 23647 15439 23653
rect 15381 23644 15393 23647
rect 15252 23616 15393 23644
rect 15252 23604 15258 23616
rect 15381 23613 15393 23616
rect 15427 23613 15439 23647
rect 15381 23607 15439 23613
rect 16390 23604 16396 23656
rect 16448 23604 16454 23656
rect 17402 23604 17408 23656
rect 17460 23604 17466 23656
rect 18782 23604 18788 23656
rect 18840 23604 18846 23656
rect 20717 23647 20775 23653
rect 20717 23613 20729 23647
rect 20763 23613 20775 23647
rect 20717 23607 20775 23613
rect 16224 23548 18828 23576
rect 16224 23520 16252 23548
rect 6549 23511 6607 23517
rect 6549 23508 6561 23511
rect 6144 23480 6561 23508
rect 6144 23468 6150 23480
rect 6549 23477 6561 23480
rect 6595 23477 6607 23511
rect 6549 23471 6607 23477
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 7064 23480 8217 23508
rect 7064 23468 7070 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8205 23471 8263 23477
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 12989 23511 13047 23517
rect 12989 23508 13001 23511
rect 12676 23480 13001 23508
rect 12676 23468 12682 23480
rect 12989 23477 13001 23480
rect 13035 23508 13047 23511
rect 13722 23508 13728 23520
rect 13035 23480 13728 23508
rect 13035 23477 13047 23480
rect 12989 23471 13047 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 14826 23468 14832 23520
rect 14884 23468 14890 23520
rect 15838 23468 15844 23520
rect 15896 23468 15902 23520
rect 16206 23468 16212 23520
rect 16264 23468 16270 23520
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 18800 23508 18828 23548
rect 19886 23536 19892 23588
rect 19944 23576 19950 23588
rect 20732 23576 20760 23607
rect 20806 23604 20812 23656
rect 20864 23644 20870 23656
rect 21928 23653 21956 23684
rect 23937 23681 23949 23715
rect 23983 23681 23995 23715
rect 23937 23675 23995 23681
rect 24029 23715 24087 23721
rect 24029 23681 24041 23715
rect 24075 23712 24087 23715
rect 24765 23715 24823 23721
rect 24075 23684 24716 23712
rect 24075 23681 24087 23684
rect 24029 23675 24087 23681
rect 21913 23647 21971 23653
rect 20864 23616 21680 23644
rect 20864 23604 20870 23616
rect 19944 23548 21404 23576
rect 19944 23536 19950 23548
rect 21376 23520 21404 23548
rect 20438 23508 20444 23520
rect 18800 23480 20444 23508
rect 20438 23468 20444 23480
rect 20496 23508 20502 23520
rect 20806 23508 20812 23520
rect 20496 23480 20812 23508
rect 20496 23468 20502 23480
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 21358 23468 21364 23520
rect 21416 23468 21422 23520
rect 21652 23508 21680 23616
rect 21913 23613 21925 23647
rect 21959 23644 21971 23647
rect 22097 23647 22155 23653
rect 21959 23616 21993 23644
rect 21959 23613 21971 23616
rect 21913 23607 21971 23613
rect 22097 23613 22109 23647
rect 22143 23613 22155 23647
rect 22649 23647 22707 23653
rect 22649 23644 22661 23647
rect 22097 23607 22155 23613
rect 22572 23616 22661 23644
rect 22002 23536 22008 23588
rect 22060 23576 22066 23588
rect 22112 23576 22140 23607
rect 22572 23585 22600 23616
rect 22649 23613 22661 23616
rect 22695 23613 22707 23647
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 22649 23607 22707 23613
rect 22756 23616 24133 23644
rect 22060 23548 22140 23576
rect 22557 23579 22615 23585
rect 22060 23536 22066 23548
rect 22557 23545 22569 23579
rect 22603 23545 22615 23579
rect 22557 23539 22615 23545
rect 22756 23508 22784 23616
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 24688 23644 24716 23684
rect 24765 23681 24777 23715
rect 24811 23712 24823 23715
rect 24872 23712 24900 23740
rect 24811 23684 24900 23712
rect 24811 23681 24823 23684
rect 24765 23675 24823 23681
rect 24854 23644 24860 23656
rect 24688 23616 24860 23644
rect 24121 23607 24179 23613
rect 24136 23576 24164 23607
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 24964 23653 24992 23752
rect 25314 23740 25320 23752
rect 25372 23740 25378 23792
rect 25866 23740 25872 23792
rect 25924 23740 25930 23792
rect 29730 23740 29736 23792
rect 29788 23780 29794 23792
rect 30374 23780 30380 23792
rect 29788 23752 30380 23780
rect 29788 23740 29794 23752
rect 30374 23740 30380 23752
rect 30432 23780 30438 23792
rect 31205 23783 31263 23789
rect 31205 23780 31217 23783
rect 30432 23752 31217 23780
rect 30432 23740 30438 23752
rect 31205 23749 31217 23752
rect 31251 23780 31263 23783
rect 32048 23780 32076 23820
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 33505 23851 33563 23857
rect 33505 23817 33517 23851
rect 33551 23848 33563 23851
rect 33686 23848 33692 23860
rect 33551 23820 33692 23848
rect 33551 23817 33563 23820
rect 33505 23811 33563 23817
rect 33686 23808 33692 23820
rect 33744 23808 33750 23860
rect 34146 23808 34152 23860
rect 34204 23848 34210 23860
rect 36633 23851 36691 23857
rect 36633 23848 36645 23851
rect 34204 23820 36645 23848
rect 34204 23808 34210 23820
rect 36633 23817 36645 23820
rect 36679 23817 36691 23851
rect 36633 23811 36691 23817
rect 37277 23851 37335 23857
rect 37277 23817 37289 23851
rect 37323 23848 37335 23851
rect 37550 23848 37556 23860
rect 37323 23820 37556 23848
rect 37323 23817 37335 23820
rect 37277 23811 37335 23817
rect 37550 23808 37556 23820
rect 37608 23808 37614 23860
rect 37645 23851 37703 23857
rect 37645 23817 37657 23851
rect 37691 23848 37703 23851
rect 38930 23848 38936 23860
rect 37691 23820 38936 23848
rect 37691 23817 37703 23820
rect 37645 23811 37703 23817
rect 38930 23808 38936 23820
rect 38988 23808 38994 23860
rect 39850 23808 39856 23860
rect 39908 23808 39914 23860
rect 40681 23851 40739 23857
rect 40681 23817 40693 23851
rect 40727 23848 40739 23851
rect 41138 23848 41144 23860
rect 40727 23820 41144 23848
rect 40727 23817 40739 23820
rect 40681 23811 40739 23817
rect 41138 23808 41144 23820
rect 41196 23808 41202 23860
rect 45646 23808 45652 23860
rect 45704 23808 45710 23860
rect 46017 23851 46075 23857
rect 46017 23817 46029 23851
rect 46063 23848 46075 23851
rect 46474 23848 46480 23860
rect 46063 23820 46480 23848
rect 46063 23817 46075 23820
rect 46017 23811 46075 23817
rect 46474 23808 46480 23820
rect 46532 23808 46538 23860
rect 48130 23808 48136 23860
rect 48188 23848 48194 23860
rect 48317 23851 48375 23857
rect 48317 23848 48329 23851
rect 48188 23820 48329 23848
rect 48188 23808 48194 23820
rect 48317 23817 48329 23820
rect 48363 23817 48375 23851
rect 48317 23811 48375 23817
rect 50433 23851 50491 23857
rect 50433 23817 50445 23851
rect 50479 23848 50491 23851
rect 50982 23848 50988 23860
rect 50479 23820 50988 23848
rect 50479 23817 50491 23820
rect 50433 23811 50491 23817
rect 50982 23808 50988 23820
rect 51040 23808 51046 23860
rect 52273 23851 52331 23857
rect 52273 23817 52285 23851
rect 52319 23848 52331 23851
rect 53282 23848 53288 23860
rect 52319 23820 53288 23848
rect 52319 23817 52331 23820
rect 52273 23811 52331 23817
rect 53282 23808 53288 23820
rect 53340 23808 53346 23860
rect 53837 23851 53895 23857
rect 53837 23817 53849 23851
rect 53883 23848 53895 23851
rect 54386 23848 54392 23860
rect 53883 23820 54392 23848
rect 53883 23817 53895 23820
rect 53837 23811 53895 23817
rect 54386 23808 54392 23820
rect 54444 23808 54450 23860
rect 55401 23851 55459 23857
rect 55401 23817 55413 23851
rect 55447 23817 55459 23851
rect 55401 23811 55459 23817
rect 34508 23783 34566 23789
rect 31251 23752 32076 23780
rect 32140 23752 34284 23780
rect 31251 23749 31263 23752
rect 31205 23743 31263 23749
rect 25676 23715 25734 23721
rect 25676 23681 25688 23715
rect 25722 23712 25734 23715
rect 26973 23715 27031 23721
rect 26973 23712 26985 23715
rect 25722 23684 26985 23712
rect 25722 23681 25734 23684
rect 25676 23675 25734 23681
rect 26973 23681 26985 23684
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 32030 23672 32036 23724
rect 32088 23712 32094 23724
rect 32140 23721 32168 23752
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 32088 23684 32137 23712
rect 32088 23672 32094 23684
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 32392 23715 32450 23721
rect 32392 23681 32404 23715
rect 32438 23712 32450 23715
rect 32950 23712 32956 23724
rect 32438 23684 32956 23712
rect 32438 23681 32450 23684
rect 32392 23675 32450 23681
rect 32950 23672 32956 23684
rect 33008 23672 33014 23724
rect 24949 23647 25007 23653
rect 24949 23613 24961 23647
rect 24995 23613 25007 23647
rect 24949 23607 25007 23613
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25409 23647 25467 23653
rect 25409 23644 25421 23647
rect 25096 23616 25421 23644
rect 25096 23604 25102 23616
rect 25409 23613 25421 23616
rect 25455 23613 25467 23647
rect 25409 23607 25467 23613
rect 27617 23647 27675 23653
rect 27617 23613 27629 23647
rect 27663 23644 27675 23647
rect 27706 23644 27712 23656
rect 27663 23616 27712 23644
rect 27663 23613 27675 23616
rect 27617 23607 27675 23613
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 29178 23604 29184 23656
rect 29236 23644 29242 23656
rect 34256 23653 34284 23752
rect 34508 23749 34520 23783
rect 34554 23780 34566 23783
rect 35434 23780 35440 23792
rect 34554 23752 35440 23780
rect 34554 23749 34566 23752
rect 34508 23743 34566 23749
rect 35434 23740 35440 23752
rect 35492 23740 35498 23792
rect 38740 23783 38798 23789
rect 37752 23752 38700 23780
rect 35526 23672 35532 23724
rect 35584 23712 35590 23724
rect 35584 23684 37596 23712
rect 35584 23672 35590 23684
rect 29733 23647 29791 23653
rect 29733 23644 29745 23647
rect 29236 23616 29745 23644
rect 29236 23604 29242 23616
rect 29733 23613 29745 23616
rect 29779 23613 29791 23647
rect 29733 23607 29791 23613
rect 34241 23647 34299 23653
rect 34241 23613 34253 23647
rect 34287 23613 34299 23647
rect 36265 23647 36323 23653
rect 36265 23644 36277 23647
rect 34241 23607 34299 23613
rect 35866 23616 36277 23644
rect 24136 23548 25084 23576
rect 21652 23480 22784 23508
rect 23106 23468 23112 23520
rect 23164 23508 23170 23520
rect 23293 23511 23351 23517
rect 23293 23508 23305 23511
rect 23164 23480 23305 23508
rect 23164 23468 23170 23480
rect 23293 23477 23305 23480
rect 23339 23477 23351 23511
rect 23293 23471 23351 23477
rect 24397 23511 24455 23517
rect 24397 23477 24409 23511
rect 24443 23508 24455 23511
rect 24854 23508 24860 23520
rect 24443 23480 24860 23508
rect 24443 23477 24455 23480
rect 24397 23471 24455 23477
rect 24854 23468 24860 23480
rect 24912 23468 24918 23520
rect 25056 23508 25084 23548
rect 27246 23508 27252 23520
rect 25056 23480 27252 23508
rect 27246 23468 27252 23480
rect 27304 23468 27310 23520
rect 28074 23468 28080 23520
rect 28132 23508 28138 23520
rect 28445 23511 28503 23517
rect 28445 23508 28457 23511
rect 28132 23480 28457 23508
rect 28132 23468 28138 23480
rect 28445 23477 28457 23480
rect 28491 23477 28503 23511
rect 28445 23471 28503 23477
rect 30377 23511 30435 23517
rect 30377 23477 30389 23511
rect 30423 23508 30435 23511
rect 30466 23508 30472 23520
rect 30423 23480 30472 23508
rect 30423 23477 30435 23480
rect 30377 23471 30435 23477
rect 30466 23468 30472 23480
rect 30524 23468 30530 23520
rect 30742 23468 30748 23520
rect 30800 23508 30806 23520
rect 31570 23508 31576 23520
rect 30800 23480 31576 23508
rect 30800 23468 30806 23480
rect 31570 23468 31576 23480
rect 31628 23468 31634 23520
rect 33873 23511 33931 23517
rect 33873 23477 33885 23511
rect 33919 23508 33931 23511
rect 34054 23508 34060 23520
rect 33919 23480 34060 23508
rect 33919 23477 33931 23480
rect 33873 23471 33931 23477
rect 34054 23468 34060 23480
rect 34112 23468 34118 23520
rect 34256 23508 34284 23607
rect 35621 23579 35679 23585
rect 35621 23545 35633 23579
rect 35667 23576 35679 23579
rect 35866 23576 35894 23616
rect 36265 23613 36277 23616
rect 36311 23613 36323 23647
rect 36265 23607 36323 23613
rect 35667 23548 35894 23576
rect 37568 23576 37596 23684
rect 37642 23604 37648 23656
rect 37700 23644 37706 23656
rect 37752 23653 37780 23752
rect 38286 23712 38292 23724
rect 37844 23684 38292 23712
rect 37737 23647 37795 23653
rect 37737 23644 37749 23647
rect 37700 23616 37749 23644
rect 37700 23604 37706 23616
rect 37737 23613 37749 23616
rect 37783 23613 37795 23647
rect 37737 23607 37795 23613
rect 37844 23576 37872 23684
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 38378 23672 38384 23724
rect 38436 23712 38442 23724
rect 38473 23715 38531 23721
rect 38473 23712 38485 23715
rect 38436 23684 38485 23712
rect 38436 23672 38442 23684
rect 38473 23681 38485 23684
rect 38519 23712 38531 23715
rect 38562 23712 38568 23724
rect 38519 23684 38568 23712
rect 38519 23681 38531 23684
rect 38473 23675 38531 23681
rect 38562 23672 38568 23684
rect 38620 23672 38626 23724
rect 38672 23712 38700 23752
rect 38740 23749 38752 23783
rect 38786 23780 38798 23783
rect 39868 23780 39896 23808
rect 38786 23752 39896 23780
rect 42429 23783 42487 23789
rect 38786 23749 38798 23752
rect 38740 23743 38798 23749
rect 42429 23749 42441 23783
rect 42475 23780 42487 23783
rect 42702 23780 42708 23792
rect 42475 23752 42708 23780
rect 42475 23749 42487 23752
rect 42429 23743 42487 23749
rect 42702 23740 42708 23752
rect 42760 23740 42766 23792
rect 42886 23740 42892 23792
rect 42944 23780 42950 23792
rect 44545 23783 44603 23789
rect 44545 23780 44557 23783
rect 42944 23752 44557 23780
rect 42944 23740 42950 23752
rect 44545 23749 44557 23752
rect 44591 23749 44603 23783
rect 45664 23780 45692 23808
rect 47857 23783 47915 23789
rect 45664 23752 46520 23780
rect 44545 23743 44603 23749
rect 40218 23712 40224 23724
rect 38672 23684 40224 23712
rect 40218 23672 40224 23684
rect 40276 23672 40282 23724
rect 40310 23672 40316 23724
rect 40368 23712 40374 23724
rect 40773 23715 40831 23721
rect 40773 23712 40785 23715
rect 40368 23684 40785 23712
rect 40368 23672 40374 23684
rect 40773 23681 40785 23684
rect 40819 23681 40831 23715
rect 40773 23675 40831 23681
rect 41340 23684 44220 23712
rect 37921 23647 37979 23653
rect 37921 23613 37933 23647
rect 37967 23613 37979 23647
rect 37921 23607 37979 23613
rect 37568 23548 37872 23576
rect 35667 23545 35679 23548
rect 35621 23539 35679 23545
rect 34514 23508 34520 23520
rect 34256 23480 34520 23508
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 35710 23468 35716 23520
rect 35768 23468 35774 23520
rect 35894 23468 35900 23520
rect 35952 23508 35958 23520
rect 37093 23511 37151 23517
rect 37093 23508 37105 23511
rect 35952 23480 37105 23508
rect 35952 23468 35958 23480
rect 37093 23477 37105 23480
rect 37139 23508 37151 23511
rect 37936 23508 37964 23607
rect 39666 23604 39672 23656
rect 39724 23644 39730 23656
rect 40037 23647 40095 23653
rect 40037 23644 40049 23647
rect 39724 23616 40049 23644
rect 39724 23604 39730 23616
rect 40037 23613 40049 23616
rect 40083 23644 40095 23647
rect 41340 23644 41368 23684
rect 40083 23616 41368 23644
rect 41417 23647 41475 23653
rect 40083 23613 40095 23616
rect 40037 23607 40095 23613
rect 41417 23613 41429 23647
rect 41463 23644 41475 23647
rect 41598 23644 41604 23656
rect 41463 23616 41604 23644
rect 41463 23613 41475 23616
rect 41417 23607 41475 23613
rect 41598 23604 41604 23616
rect 41656 23604 41662 23656
rect 42061 23647 42119 23653
rect 42061 23613 42073 23647
rect 42107 23613 42119 23647
rect 44192 23644 44220 23684
rect 44266 23672 44272 23724
rect 44324 23712 44330 23724
rect 44634 23712 44640 23724
rect 44324 23684 44640 23712
rect 44324 23672 44330 23684
rect 44634 23672 44640 23684
rect 44692 23672 44698 23724
rect 46492 23721 46520 23752
rect 47857 23749 47869 23783
rect 47903 23780 47915 23783
rect 49050 23780 49056 23792
rect 47903 23752 49056 23780
rect 47903 23749 47915 23752
rect 47857 23743 47915 23749
rect 49050 23740 49056 23752
rect 49108 23740 49114 23792
rect 51905 23783 51963 23789
rect 51905 23780 51917 23783
rect 50816 23752 51917 23780
rect 50816 23724 50844 23752
rect 51905 23749 51917 23752
rect 51951 23749 51963 23783
rect 51905 23743 51963 23749
rect 54205 23783 54263 23789
rect 54205 23749 54217 23783
rect 54251 23780 54263 23783
rect 55214 23780 55220 23792
rect 54251 23752 55220 23780
rect 54251 23749 54263 23752
rect 54205 23743 54263 23749
rect 55214 23740 55220 23752
rect 55272 23740 55278 23792
rect 55416 23780 55444 23811
rect 56594 23789 56600 23792
rect 56588 23780 56600 23789
rect 55416 23752 56180 23780
rect 56555 23752 56600 23780
rect 46385 23715 46443 23721
rect 46385 23681 46397 23715
rect 46431 23681 46443 23715
rect 46385 23675 46443 23681
rect 46477 23715 46535 23721
rect 46477 23681 46489 23715
rect 46523 23712 46535 23715
rect 46566 23712 46572 23724
rect 46523 23684 46572 23712
rect 46523 23681 46535 23684
rect 46477 23675 46535 23681
rect 44453 23647 44511 23653
rect 44453 23644 44465 23647
rect 44192 23616 44465 23644
rect 42061 23607 42119 23613
rect 44453 23613 44465 23616
rect 44499 23644 44511 23647
rect 45278 23644 45284 23656
rect 44499 23616 45284 23644
rect 44499 23613 44511 23616
rect 44453 23607 44511 23613
rect 39853 23579 39911 23585
rect 39853 23545 39865 23579
rect 39899 23576 39911 23579
rect 42076 23576 42104 23607
rect 45278 23604 45284 23616
rect 45336 23604 45342 23656
rect 45649 23647 45707 23653
rect 45649 23613 45661 23647
rect 45695 23613 45707 23647
rect 45649 23607 45707 23613
rect 39899 23548 42104 23576
rect 45005 23579 45063 23585
rect 39899 23545 39911 23548
rect 39853 23539 39911 23545
rect 45005 23545 45017 23579
rect 45051 23576 45063 23579
rect 45664 23576 45692 23607
rect 45051 23548 45692 23576
rect 46400 23576 46428 23675
rect 46566 23672 46572 23684
rect 46624 23712 46630 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 46624 23684 47961 23712
rect 46624 23672 46630 23684
rect 47949 23681 47961 23684
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 50798 23672 50804 23724
rect 50856 23672 50862 23724
rect 50893 23715 50951 23721
rect 50893 23681 50905 23715
rect 50939 23712 50951 23715
rect 50939 23684 51396 23712
rect 50939 23681 50951 23684
rect 50893 23675 50951 23681
rect 51368 23656 51396 23684
rect 51994 23672 52000 23724
rect 52052 23712 52058 23724
rect 52917 23715 52975 23721
rect 52917 23712 52929 23715
rect 52052 23684 52929 23712
rect 52052 23672 52058 23684
rect 52917 23681 52929 23684
rect 52963 23681 52975 23715
rect 52917 23675 52975 23681
rect 54297 23715 54355 23721
rect 54297 23681 54309 23715
rect 54343 23712 54355 23715
rect 54941 23715 54999 23721
rect 54941 23712 54953 23715
rect 54343 23684 54953 23712
rect 54343 23681 54355 23684
rect 54297 23675 54355 23681
rect 54941 23681 54953 23684
rect 54987 23681 54999 23715
rect 54941 23675 54999 23681
rect 55033 23715 55091 23721
rect 55033 23681 55045 23715
rect 55079 23712 55091 23715
rect 55766 23712 55772 23724
rect 55079 23684 55772 23712
rect 55079 23681 55091 23684
rect 55033 23675 55091 23681
rect 46658 23604 46664 23656
rect 46716 23644 46722 23656
rect 47029 23647 47087 23653
rect 47029 23644 47041 23647
rect 46716 23616 47041 23644
rect 46716 23604 46722 23616
rect 47029 23613 47041 23616
rect 47075 23613 47087 23647
rect 47029 23607 47087 23613
rect 47486 23604 47492 23656
rect 47544 23644 47550 23656
rect 47673 23647 47731 23653
rect 47673 23644 47685 23647
rect 47544 23616 47685 23644
rect 47544 23604 47550 23616
rect 47673 23613 47685 23616
rect 47719 23644 47731 23647
rect 47719 23616 48452 23644
rect 47719 23613 47731 23616
rect 47673 23607 47731 23613
rect 48314 23576 48320 23588
rect 46400 23548 48320 23576
rect 45051 23545 45063 23548
rect 45005 23539 45063 23545
rect 48314 23536 48320 23548
rect 48372 23536 48378 23588
rect 48424 23576 48452 23616
rect 48498 23604 48504 23656
rect 48556 23604 48562 23656
rect 50246 23604 50252 23656
rect 50304 23644 50310 23656
rect 50985 23647 51043 23653
rect 50985 23644 50997 23647
rect 50304 23616 50997 23644
rect 50304 23604 50310 23616
rect 50985 23613 50997 23616
rect 51031 23613 51043 23647
rect 50985 23607 51043 23613
rect 51350 23604 51356 23656
rect 51408 23604 51414 23656
rect 51629 23647 51687 23653
rect 51629 23613 51641 23647
rect 51675 23613 51687 23647
rect 51629 23607 51687 23613
rect 51813 23647 51871 23653
rect 51813 23613 51825 23647
rect 51859 23644 51871 23647
rect 52454 23644 52460 23656
rect 51859 23616 52460 23644
rect 51859 23613 51871 23616
rect 51813 23607 51871 23613
rect 49881 23579 49939 23585
rect 49881 23576 49893 23579
rect 48424 23548 49893 23576
rect 49881 23545 49893 23548
rect 49927 23576 49939 23579
rect 51644 23576 51672 23607
rect 52454 23604 52460 23616
rect 52512 23604 52518 23656
rect 53650 23604 53656 23656
rect 53708 23644 53714 23656
rect 54389 23647 54447 23653
rect 54389 23644 54401 23647
rect 53708 23616 54401 23644
rect 53708 23604 53714 23616
rect 54389 23613 54401 23616
rect 54435 23613 54447 23647
rect 54389 23607 54447 23613
rect 54570 23604 54576 23656
rect 54628 23644 54634 23656
rect 54757 23647 54815 23653
rect 54757 23644 54769 23647
rect 54628 23616 54769 23644
rect 54628 23604 54634 23616
rect 54757 23613 54769 23616
rect 54803 23613 54815 23647
rect 54757 23607 54815 23613
rect 49927 23548 51672 23576
rect 54956 23576 54984 23675
rect 55766 23672 55772 23684
rect 55824 23672 55830 23724
rect 56152 23721 56180 23752
rect 56588 23743 56600 23752
rect 56594 23740 56600 23743
rect 56652 23740 56658 23792
rect 56137 23715 56195 23721
rect 56137 23681 56149 23715
rect 56183 23681 56195 23715
rect 56137 23675 56195 23681
rect 56318 23604 56324 23656
rect 56376 23604 56382 23656
rect 57606 23604 57612 23656
rect 57664 23644 57670 23656
rect 58437 23647 58495 23653
rect 58437 23644 58449 23647
rect 57664 23616 58449 23644
rect 57664 23604 57670 23616
rect 58437 23613 58449 23616
rect 58483 23613 58495 23647
rect 58437 23607 58495 23613
rect 57701 23579 57759 23585
rect 54956 23548 55628 23576
rect 49927 23545 49939 23548
rect 49881 23539 49939 23545
rect 41230 23508 41236 23520
rect 37139 23480 41236 23508
rect 37139 23477 37151 23480
rect 37093 23471 37151 23477
rect 41230 23468 41236 23480
rect 41288 23468 41294 23520
rect 41506 23468 41512 23520
rect 41564 23468 41570 23520
rect 42518 23468 42524 23520
rect 42576 23508 42582 23520
rect 43901 23511 43959 23517
rect 43901 23508 43913 23511
rect 42576 23480 43913 23508
rect 42576 23468 42582 23480
rect 43901 23477 43913 23480
rect 43947 23508 43959 23511
rect 44634 23508 44640 23520
rect 43947 23480 44640 23508
rect 43947 23477 43959 23480
rect 43901 23471 43959 23477
rect 44634 23468 44640 23480
rect 44692 23468 44698 23520
rect 45094 23468 45100 23520
rect 45152 23468 45158 23520
rect 45278 23468 45284 23520
rect 45336 23508 45342 23520
rect 48682 23508 48688 23520
rect 45336 23480 48688 23508
rect 45336 23468 45342 23480
rect 48682 23468 48688 23480
rect 48740 23468 48746 23520
rect 50246 23468 50252 23520
rect 50304 23468 50310 23520
rect 53098 23468 53104 23520
rect 53156 23508 53162 23520
rect 53561 23511 53619 23517
rect 53561 23508 53573 23511
rect 53156 23480 53573 23508
rect 53156 23468 53162 23480
rect 53561 23477 53573 23480
rect 53607 23477 53619 23511
rect 53561 23471 53619 23477
rect 55490 23468 55496 23520
rect 55548 23468 55554 23520
rect 55600 23508 55628 23548
rect 57701 23545 57713 23579
rect 57747 23576 57759 23579
rect 58066 23576 58072 23588
rect 57747 23548 58072 23576
rect 57747 23545 57759 23548
rect 57701 23539 57759 23545
rect 58066 23536 58072 23548
rect 58124 23536 58130 23588
rect 57790 23508 57796 23520
rect 55600 23480 57796 23508
rect 57790 23468 57796 23480
rect 57848 23468 57854 23520
rect 57882 23468 57888 23520
rect 57940 23468 57946 23520
rect 1104 23418 58880 23440
rect 1104 23366 8172 23418
rect 8224 23366 8236 23418
rect 8288 23366 8300 23418
rect 8352 23366 8364 23418
rect 8416 23366 8428 23418
rect 8480 23366 22616 23418
rect 22668 23366 22680 23418
rect 22732 23366 22744 23418
rect 22796 23366 22808 23418
rect 22860 23366 22872 23418
rect 22924 23366 37060 23418
rect 37112 23366 37124 23418
rect 37176 23366 37188 23418
rect 37240 23366 37252 23418
rect 37304 23366 37316 23418
rect 37368 23366 51504 23418
rect 51556 23366 51568 23418
rect 51620 23366 51632 23418
rect 51684 23366 51696 23418
rect 51748 23366 51760 23418
rect 51812 23366 58880 23418
rect 1104 23344 58880 23366
rect 4522 23264 4528 23316
rect 4580 23264 4586 23316
rect 5350 23264 5356 23316
rect 5408 23304 5414 23316
rect 5537 23307 5595 23313
rect 5537 23304 5549 23307
rect 5408 23276 5549 23304
rect 5408 23264 5414 23276
rect 5537 23273 5549 23276
rect 5583 23273 5595 23307
rect 5537 23267 5595 23273
rect 12253 23307 12311 23313
rect 12253 23273 12265 23307
rect 12299 23304 12311 23307
rect 12342 23304 12348 23316
rect 12299 23276 12348 23304
rect 12299 23273 12311 23276
rect 12253 23267 12311 23273
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 15933 23307 15991 23313
rect 15933 23273 15945 23307
rect 15979 23304 15991 23307
rect 16390 23304 16396 23316
rect 15979 23276 16396 23304
rect 15979 23273 15991 23276
rect 15933 23267 15991 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 22094 23304 22100 23316
rect 19392 23276 20116 23304
rect 19392 23264 19398 23276
rect 4706 23128 4712 23180
rect 4764 23168 4770 23180
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 4764 23140 5089 23168
rect 4764 23128 4770 23140
rect 5077 23137 5089 23140
rect 5123 23137 5135 23171
rect 5077 23131 5135 23137
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11388 23140 11621 23168
rect 11388 23128 11394 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 17313 23171 17371 23177
rect 17313 23137 17325 23171
rect 17359 23168 17371 23171
rect 18782 23168 18788 23180
rect 17359 23140 18788 23168
rect 17359 23137 17371 23140
rect 17313 23131 17371 23137
rect 13538 23060 13544 23112
rect 13596 23060 13602 23112
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 13780 23072 14473 23100
rect 13780 23060 13786 23072
rect 14461 23069 14473 23072
rect 14507 23100 14519 23103
rect 15102 23100 15108 23112
rect 14507 23072 15108 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 15102 23060 15108 23072
rect 15160 23100 15166 23112
rect 17328 23100 17356 23131
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 19886 23128 19892 23180
rect 19944 23128 19950 23180
rect 20088 23177 20116 23276
rect 20732 23276 22100 23304
rect 20732 23177 20760 23276
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 24210 23264 24216 23316
rect 24268 23264 24274 23316
rect 25133 23307 25191 23313
rect 25133 23273 25145 23307
rect 25179 23304 25191 23307
rect 26786 23304 26792 23316
rect 25179 23276 26792 23304
rect 25179 23273 25191 23276
rect 25133 23267 25191 23273
rect 26786 23264 26792 23276
rect 26844 23264 26850 23316
rect 27065 23307 27123 23313
rect 27065 23273 27077 23307
rect 27111 23304 27123 23307
rect 27706 23304 27712 23316
rect 27111 23276 27712 23304
rect 27111 23273 27123 23276
rect 27065 23267 27123 23273
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 33413 23307 33471 23313
rect 33413 23273 33425 23307
rect 33459 23304 33471 23307
rect 33502 23304 33508 23316
rect 33459 23276 33508 23304
rect 33459 23273 33471 23276
rect 33413 23267 33471 23273
rect 33502 23264 33508 23276
rect 33560 23264 33566 23316
rect 36630 23304 36636 23316
rect 34532 23276 36636 23304
rect 28629 23239 28687 23245
rect 28629 23205 28641 23239
rect 28675 23205 28687 23239
rect 28629 23199 28687 23205
rect 29656 23208 30788 23236
rect 20073 23171 20131 23177
rect 20073 23137 20085 23171
rect 20119 23137 20131 23171
rect 20073 23131 20131 23137
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23137 20775 23171
rect 20717 23131 20775 23137
rect 21174 23128 21180 23180
rect 21232 23128 21238 23180
rect 21266 23128 21272 23180
rect 21324 23168 21330 23180
rect 21570 23171 21628 23177
rect 21570 23168 21582 23171
rect 21324 23140 21582 23168
rect 21324 23128 21330 23140
rect 21570 23137 21582 23140
rect 21616 23137 21628 23171
rect 21570 23131 21628 23137
rect 21744 23140 22416 23168
rect 21744 23112 21772 23140
rect 15160 23072 17356 23100
rect 17957 23103 18015 23109
rect 15160 23060 15166 23072
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 18555 23072 19472 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 12897 23035 12955 23041
rect 12897 23001 12909 23035
rect 12943 23032 12955 23035
rect 14728 23035 14786 23041
rect 12943 23004 13308 23032
rect 12943 23001 12955 23004
rect 12897 22995 12955 23001
rect 13280 22976 13308 23004
rect 14728 23001 14740 23035
rect 14774 23032 14786 23035
rect 14826 23032 14832 23044
rect 14774 23004 14832 23032
rect 14774 23001 14786 23004
rect 14728 22995 14786 23001
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 16850 22992 16856 23044
rect 16908 23032 16914 23044
rect 17046 23035 17104 23041
rect 17046 23032 17058 23035
rect 16908 23004 17058 23032
rect 16908 22992 16914 23004
rect 17046 23001 17058 23004
rect 17092 23001 17104 23035
rect 17972 23032 18000 23063
rect 17046 22995 17104 23001
rect 17328 23004 18000 23032
rect 8570 22924 8576 22976
rect 8628 22964 8634 22976
rect 9125 22967 9183 22973
rect 9125 22964 9137 22967
rect 8628 22936 9137 22964
rect 8628 22924 8634 22936
rect 9125 22933 9137 22936
rect 9171 22933 9183 22967
rect 9125 22927 9183 22933
rect 12986 22924 12992 22976
rect 13044 22924 13050 22976
rect 13262 22924 13268 22976
rect 13320 22924 13326 22976
rect 15841 22967 15899 22973
rect 15841 22933 15853 22967
rect 15887 22964 15899 22967
rect 17328 22964 17356 23004
rect 15887 22936 17356 22964
rect 17405 22967 17463 22973
rect 15887 22933 15899 22936
rect 15841 22927 15899 22933
rect 17405 22933 17417 22967
rect 17451 22964 17463 22967
rect 17586 22964 17592 22976
rect 17451 22936 17592 22964
rect 17451 22933 17463 22936
rect 17405 22927 17463 22933
rect 17586 22924 17592 22936
rect 17644 22924 17650 22976
rect 19058 22924 19064 22976
rect 19116 22924 19122 22976
rect 19444 22973 19472 23072
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20533 23103 20591 23109
rect 20533 23100 20545 23103
rect 20220 23072 20545 23100
rect 20220 23060 20226 23072
rect 20533 23069 20545 23072
rect 20579 23069 20591 23103
rect 20533 23063 20591 23069
rect 21450 23060 21456 23112
rect 21508 23060 21514 23112
rect 21726 23060 21732 23112
rect 21784 23060 21790 23112
rect 22388 23100 22416 23140
rect 22462 23128 22468 23180
rect 22520 23168 22526 23180
rect 22833 23171 22891 23177
rect 22833 23168 22845 23171
rect 22520 23140 22845 23168
rect 22520 23128 22526 23140
rect 22833 23137 22845 23140
rect 22879 23137 22891 23171
rect 22833 23131 22891 23137
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 24949 23171 25007 23177
rect 24949 23168 24961 23171
rect 24912 23140 24961 23168
rect 24912 23128 24918 23140
rect 24949 23137 24961 23140
rect 24995 23137 25007 23171
rect 24949 23131 25007 23137
rect 26050 23128 26056 23180
rect 26108 23128 26114 23180
rect 26326 23128 26332 23180
rect 26384 23128 26390 23180
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 26835 23140 27476 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 22649 23103 22707 23109
rect 22649 23100 22661 23103
rect 22388 23072 22661 23100
rect 22649 23069 22661 23072
rect 22695 23069 22707 23103
rect 22649 23063 22707 23069
rect 23100 23103 23158 23109
rect 23100 23069 23112 23103
rect 23146 23100 23158 23103
rect 23382 23100 23388 23112
rect 23146 23072 23388 23100
rect 23146 23069 23158 23072
rect 23100 23063 23158 23069
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 25774 23060 25780 23112
rect 25832 23060 25838 23112
rect 25866 23060 25872 23112
rect 25924 23109 25930 23112
rect 27448 23109 27476 23140
rect 27522 23128 27528 23180
rect 27580 23168 27586 23180
rect 27617 23171 27675 23177
rect 27617 23168 27629 23171
rect 27580 23140 27629 23168
rect 27580 23128 27586 23140
rect 27617 23137 27629 23140
rect 27663 23137 27675 23171
rect 27617 23131 27675 23137
rect 28074 23128 28080 23180
rect 28132 23128 28138 23180
rect 28537 23171 28595 23177
rect 28537 23137 28549 23171
rect 28583 23168 28595 23171
rect 28644 23168 28672 23199
rect 29656 23180 29684 23208
rect 28583 23140 28672 23168
rect 29181 23171 29239 23177
rect 28583 23137 28595 23140
rect 28537 23131 28595 23137
rect 29181 23137 29193 23171
rect 29227 23137 29239 23171
rect 29181 23131 29239 23137
rect 25924 23103 25973 23109
rect 25924 23069 25927 23103
rect 25961 23069 25973 23103
rect 25924 23063 25973 23069
rect 26973 23103 27031 23109
rect 26973 23069 26985 23103
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 27433 23103 27491 23109
rect 27433 23069 27445 23103
rect 27479 23100 27491 23103
rect 27798 23100 27804 23112
rect 27479 23072 27804 23100
rect 27479 23069 27491 23072
rect 27433 23063 27491 23069
rect 25924 23060 25930 23063
rect 19797 23035 19855 23041
rect 19797 23001 19809 23035
rect 19843 23032 19855 23035
rect 19843 23004 20760 23032
rect 19843 23001 19855 23004
rect 19797 22995 19855 23001
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22933 19487 22967
rect 20732 22964 20760 23004
rect 21450 22964 21456 22976
rect 20732 22936 21456 22964
rect 19429 22927 19487 22933
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 22278 22924 22284 22976
rect 22336 22964 22342 22976
rect 22373 22967 22431 22973
rect 22373 22964 22385 22967
rect 22336 22936 22385 22964
rect 22336 22924 22342 22936
rect 22373 22933 22385 22936
rect 22419 22933 22431 22967
rect 22373 22927 22431 22933
rect 24394 22924 24400 22976
rect 24452 22924 24458 22976
rect 25958 22924 25964 22976
rect 26016 22964 26022 22976
rect 26988 22964 27016 23063
rect 27798 23060 27804 23072
rect 27856 23060 27862 23112
rect 28092 23100 28120 23128
rect 29196 23100 29224 23131
rect 29638 23128 29644 23180
rect 29696 23128 29702 23180
rect 30650 23128 30656 23180
rect 30708 23128 30714 23180
rect 30760 23177 30788 23208
rect 31570 23196 31576 23248
rect 31628 23196 31634 23248
rect 30745 23171 30803 23177
rect 30745 23137 30757 23171
rect 30791 23137 30803 23171
rect 31588 23168 31616 23196
rect 31588 23140 31708 23168
rect 30745 23131 30803 23137
rect 28092 23072 29224 23100
rect 31570 23060 31576 23112
rect 31628 23060 31634 23112
rect 29089 23035 29147 23041
rect 29089 23001 29101 23035
rect 29135 23032 29147 23035
rect 30466 23032 30472 23044
rect 29135 23004 30472 23032
rect 29135 23001 29147 23004
rect 29089 22995 29147 23001
rect 30466 22992 30472 23004
rect 30524 22992 30530 23044
rect 26016 22936 27016 22964
rect 26016 22924 26022 22936
rect 27522 22924 27528 22976
rect 27580 22924 27586 22976
rect 27890 22924 27896 22976
rect 27948 22924 27954 22976
rect 28994 22924 29000 22976
rect 29052 22924 29058 22976
rect 29638 22924 29644 22976
rect 29696 22964 29702 22976
rect 30009 22967 30067 22973
rect 30009 22964 30021 22967
rect 29696 22936 30021 22964
rect 29696 22924 29702 22936
rect 30009 22933 30021 22936
rect 30055 22933 30067 22967
rect 30009 22927 30067 22933
rect 30193 22967 30251 22973
rect 30193 22933 30205 22967
rect 30239 22964 30251 22967
rect 30374 22964 30380 22976
rect 30239 22936 30380 22964
rect 30239 22933 30251 22936
rect 30193 22927 30251 22933
rect 30374 22924 30380 22936
rect 30432 22924 30438 22976
rect 30558 22924 30564 22976
rect 30616 22924 30622 22976
rect 31018 22924 31024 22976
rect 31076 22924 31082 22976
rect 31680 22964 31708 23140
rect 34054 23128 34060 23180
rect 34112 23168 34118 23180
rect 34532 23168 34560 23276
rect 36630 23264 36636 23276
rect 36688 23264 36694 23316
rect 37734 23264 37740 23316
rect 37792 23264 37798 23316
rect 38286 23264 38292 23316
rect 38344 23304 38350 23316
rect 39853 23307 39911 23313
rect 38344 23276 39068 23304
rect 38344 23264 38350 23276
rect 39040 23248 39068 23276
rect 39853 23273 39865 23307
rect 39899 23304 39911 23307
rect 40402 23304 40408 23316
rect 39899 23276 40408 23304
rect 39899 23273 39911 23276
rect 39853 23267 39911 23273
rect 40402 23264 40408 23276
rect 40460 23264 40466 23316
rect 41506 23304 41512 23316
rect 40512 23276 41512 23304
rect 39022 23196 39028 23248
rect 39080 23196 39086 23248
rect 34112 23140 34560 23168
rect 34112 23128 34118 23140
rect 38286 23128 38292 23180
rect 38344 23168 38350 23180
rect 38473 23171 38531 23177
rect 38473 23168 38485 23171
rect 38344 23140 38485 23168
rect 38344 23128 38350 23140
rect 38473 23137 38485 23140
rect 38519 23137 38531 23171
rect 38473 23131 38531 23137
rect 38632 23171 38690 23177
rect 38632 23137 38644 23171
rect 38678 23168 38690 23171
rect 38930 23168 38936 23180
rect 38678 23140 38936 23168
rect 38678 23137 38690 23140
rect 38632 23131 38690 23137
rect 38930 23128 38936 23140
rect 38988 23128 38994 23180
rect 39485 23171 39543 23177
rect 39485 23137 39497 23171
rect 39531 23168 39543 23171
rect 40310 23168 40316 23180
rect 39531 23140 40316 23168
rect 39531 23137 39543 23140
rect 39485 23131 39543 23137
rect 40310 23128 40316 23140
rect 40368 23128 40374 23180
rect 40402 23128 40408 23180
rect 40460 23128 40466 23180
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32030 23100 32036 23112
rect 31987 23072 32036 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32030 23060 32036 23072
rect 32088 23060 32094 23112
rect 33781 23103 33839 23109
rect 33781 23069 33793 23103
rect 33827 23100 33839 23103
rect 34330 23100 34336 23112
rect 33827 23072 34336 23100
rect 33827 23069 33839 23072
rect 33781 23063 33839 23069
rect 34330 23060 34336 23072
rect 34388 23060 34394 23112
rect 34514 23060 34520 23112
rect 34572 23100 34578 23112
rect 34701 23103 34759 23109
rect 34701 23100 34713 23103
rect 34572 23072 34713 23100
rect 34572 23060 34578 23072
rect 34701 23069 34713 23072
rect 34747 23100 34759 23103
rect 36357 23103 36415 23109
rect 36357 23100 36369 23103
rect 34747 23072 36369 23100
rect 34747 23069 34759 23072
rect 34701 23063 34759 23069
rect 36357 23069 36369 23072
rect 36403 23100 36415 23103
rect 36906 23100 36912 23112
rect 36403 23072 36912 23100
rect 36403 23069 36415 23072
rect 36357 23063 36415 23069
rect 36906 23060 36912 23072
rect 36964 23060 36970 23112
rect 38746 23060 38752 23112
rect 38804 23060 38810 23112
rect 39669 23103 39727 23109
rect 39669 23069 39681 23103
rect 39715 23100 39727 23103
rect 40512 23100 40540 23276
rect 41506 23264 41512 23276
rect 41564 23264 41570 23316
rect 44266 23304 44272 23316
rect 42904 23276 44272 23304
rect 42610 23128 42616 23180
rect 42668 23168 42674 23180
rect 42904 23177 42932 23276
rect 44266 23264 44272 23276
rect 44324 23264 44330 23316
rect 45278 23264 45284 23316
rect 45336 23264 45342 23316
rect 46750 23264 46756 23316
rect 46808 23304 46814 23316
rect 46845 23307 46903 23313
rect 46845 23304 46857 23307
rect 46808 23276 46857 23304
rect 46808 23264 46814 23276
rect 46845 23273 46857 23276
rect 46891 23273 46903 23307
rect 46845 23267 46903 23273
rect 48498 23264 48504 23316
rect 48556 23264 48562 23316
rect 51537 23307 51595 23313
rect 51537 23273 51549 23307
rect 51583 23304 51595 23307
rect 51902 23304 51908 23316
rect 51583 23276 51908 23304
rect 51583 23273 51595 23276
rect 51537 23267 51595 23273
rect 51902 23264 51908 23276
rect 51960 23264 51966 23316
rect 52638 23304 52644 23316
rect 52104 23276 52644 23304
rect 51629 23239 51687 23245
rect 51629 23205 51641 23239
rect 51675 23236 51687 23239
rect 52104 23236 52132 23276
rect 52638 23264 52644 23276
rect 52696 23264 52702 23316
rect 54849 23307 54907 23313
rect 54849 23273 54861 23307
rect 54895 23304 54907 23307
rect 55306 23304 55312 23316
rect 54895 23276 55312 23304
rect 54895 23273 54907 23276
rect 54849 23267 54907 23273
rect 55306 23264 55312 23276
rect 55364 23264 55370 23316
rect 55766 23264 55772 23316
rect 55824 23304 55830 23316
rect 55824 23276 56447 23304
rect 55824 23264 55830 23276
rect 51675 23208 52132 23236
rect 51675 23205 51687 23208
rect 51629 23199 51687 23205
rect 42705 23171 42763 23177
rect 42705 23168 42717 23171
rect 42668 23140 42717 23168
rect 42668 23128 42674 23140
rect 42705 23137 42717 23140
rect 42751 23137 42763 23171
rect 42705 23131 42763 23137
rect 42889 23171 42947 23177
rect 42889 23137 42901 23171
rect 42935 23137 42947 23171
rect 42889 23131 42947 23137
rect 43349 23171 43407 23177
rect 43349 23137 43361 23171
rect 43395 23168 43407 23171
rect 43438 23168 43444 23180
rect 43395 23140 43444 23168
rect 43395 23137 43407 23140
rect 43349 23131 43407 23137
rect 43438 23128 43444 23140
rect 43496 23128 43502 23180
rect 43901 23171 43959 23177
rect 43901 23137 43913 23171
rect 43947 23168 43959 23171
rect 43947 23140 45048 23168
rect 43947 23137 43959 23140
rect 43901 23131 43959 23137
rect 45020 23112 45048 23140
rect 56042 23128 56048 23180
rect 56100 23177 56106 23180
rect 56100 23171 56149 23177
rect 56100 23137 56103 23171
rect 56137 23137 56149 23171
rect 56100 23131 56149 23137
rect 56229 23171 56287 23177
rect 56229 23137 56241 23171
rect 56275 23168 56287 23171
rect 56419 23168 56447 23276
rect 57238 23264 57244 23316
rect 57296 23264 57302 23316
rect 58253 23239 58311 23245
rect 58253 23236 58265 23239
rect 57808 23208 58265 23236
rect 56275 23140 56447 23168
rect 56275 23137 56287 23140
rect 56229 23131 56287 23137
rect 56100 23128 56106 23131
rect 56502 23128 56508 23180
rect 56560 23128 56566 23180
rect 57808 23177 57836 23208
rect 58253 23205 58265 23208
rect 58299 23205 58311 23239
rect 58253 23199 58311 23205
rect 57793 23171 57851 23177
rect 57793 23168 57805 23171
rect 57072 23140 57805 23168
rect 39715 23072 40540 23100
rect 39715 23069 39727 23072
rect 39669 23063 39727 23069
rect 32208 23035 32266 23041
rect 32208 23001 32220 23035
rect 32254 23032 32266 23035
rect 32306 23032 32312 23044
rect 32254 23004 32312 23032
rect 32254 23001 32266 23004
rect 32208 22995 32266 23001
rect 32306 22992 32312 23004
rect 32364 22992 32370 23044
rect 34606 23032 34612 23044
rect 33060 23004 34612 23032
rect 33060 22964 33088 23004
rect 34606 22992 34612 23004
rect 34664 23032 34670 23044
rect 34968 23035 35026 23041
rect 34664 23004 34928 23032
rect 34664 22992 34670 23004
rect 31680 22936 33088 22964
rect 33318 22924 33324 22976
rect 33376 22924 33382 22976
rect 33873 22967 33931 22973
rect 33873 22933 33885 22967
rect 33919 22964 33931 22967
rect 34790 22964 34796 22976
rect 33919 22936 34796 22964
rect 33919 22933 33931 22936
rect 33873 22927 33931 22933
rect 34790 22924 34796 22936
rect 34848 22924 34854 22976
rect 34900 22964 34928 23004
rect 34968 23001 34980 23035
rect 35014 23032 35026 23035
rect 36170 23032 36176 23044
rect 35014 23004 36176 23032
rect 35014 23001 35026 23004
rect 34968 22995 35026 23001
rect 36170 22992 36176 23004
rect 36228 22992 36234 23044
rect 36624 23035 36682 23041
rect 36624 23001 36636 23035
rect 36670 23032 36682 23035
rect 36814 23032 36820 23044
rect 36670 23004 36820 23032
rect 36670 23001 36682 23004
rect 36624 22995 36682 23001
rect 36814 22992 36820 23004
rect 36872 22992 36878 23044
rect 40218 22992 40224 23044
rect 40276 22992 40282 23044
rect 40313 23035 40371 23041
rect 40313 23001 40325 23035
rect 40359 23032 40371 23035
rect 40512 23032 40540 23072
rect 41233 23103 41291 23109
rect 41233 23069 41245 23103
rect 41279 23100 41291 23103
rect 41279 23072 41368 23100
rect 41279 23069 41291 23072
rect 41233 23063 41291 23069
rect 41340 23044 41368 23072
rect 43622 23060 43628 23112
rect 43680 23060 43686 23112
rect 43714 23060 43720 23112
rect 43772 23109 43778 23112
rect 43772 23103 43800 23109
rect 43788 23069 43800 23103
rect 43772 23063 43800 23069
rect 43772 23060 43778 23063
rect 45002 23060 45008 23112
rect 45060 23060 45066 23112
rect 45462 23060 45468 23112
rect 45520 23100 45526 23112
rect 47394 23109 47400 23112
rect 47121 23103 47179 23109
rect 47121 23100 47133 23103
rect 45520 23072 47133 23100
rect 45520 23060 45526 23072
rect 47121 23069 47133 23072
rect 47167 23069 47179 23103
rect 47388 23100 47400 23109
rect 47355 23072 47400 23100
rect 47121 23063 47179 23069
rect 47388 23063 47400 23072
rect 47394 23060 47400 23063
rect 47452 23060 47458 23112
rect 50157 23103 50215 23109
rect 50157 23069 50169 23103
rect 50203 23100 50215 23103
rect 51258 23100 51264 23112
rect 50203 23072 51264 23100
rect 50203 23069 50215 23072
rect 50157 23063 50215 23069
rect 51258 23060 51264 23072
rect 51316 23100 51322 23112
rect 53009 23103 53067 23109
rect 53009 23100 53021 23103
rect 51316 23072 53021 23100
rect 51316 23060 51322 23072
rect 53009 23069 53021 23072
rect 53055 23100 53067 23103
rect 53469 23103 53527 23109
rect 53469 23100 53481 23103
rect 53055 23072 53481 23100
rect 53055 23069 53067 23072
rect 53009 23063 53067 23069
rect 53469 23069 53481 23072
rect 53515 23100 53527 23103
rect 53515 23072 53604 23100
rect 53515 23069 53527 23072
rect 53469 23063 53527 23069
rect 40359 23004 40540 23032
rect 40359 23001 40371 23004
rect 40313 22995 40371 23001
rect 41322 22992 41328 23044
rect 41380 22992 41386 23044
rect 41506 23041 41512 23044
rect 41500 22995 41512 23041
rect 41506 22992 41512 22995
rect 41564 22992 41570 23044
rect 45554 23032 45560 23044
rect 44376 23004 45560 23032
rect 35526 22964 35532 22976
rect 34900 22936 35532 22964
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 36078 22924 36084 22976
rect 36136 22924 36142 22976
rect 37829 22967 37887 22973
rect 37829 22933 37841 22967
rect 37875 22964 37887 22967
rect 40034 22964 40040 22976
rect 37875 22936 40040 22964
rect 37875 22933 37887 22936
rect 37829 22927 37887 22933
rect 40034 22924 40040 22936
rect 40092 22924 40098 22976
rect 40402 22924 40408 22976
rect 40460 22964 40466 22976
rect 40954 22964 40960 22976
rect 40460 22936 40960 22964
rect 40460 22924 40466 22936
rect 40954 22924 40960 22936
rect 41012 22964 41018 22976
rect 42242 22964 42248 22976
rect 41012 22936 42248 22964
rect 41012 22924 41018 22936
rect 42242 22924 42248 22936
rect 42300 22924 42306 22976
rect 42613 22967 42671 22973
rect 42613 22933 42625 22967
rect 42659 22964 42671 22967
rect 43070 22964 43076 22976
rect 42659 22936 43076 22964
rect 42659 22933 42671 22936
rect 42613 22927 42671 22933
rect 43070 22924 43076 22936
rect 43128 22924 43134 22976
rect 43438 22924 43444 22976
rect 43496 22964 43502 22976
rect 44376 22964 44404 23004
rect 45554 22992 45560 23004
rect 45612 22992 45618 23044
rect 45732 23035 45790 23041
rect 45732 23001 45744 23035
rect 45778 23032 45790 23035
rect 45922 23032 45928 23044
rect 45778 23004 45928 23032
rect 45778 23001 45790 23004
rect 45732 22995 45790 23001
rect 45922 22992 45928 23004
rect 45980 22992 45986 23044
rect 46842 22992 46848 23044
rect 46900 23032 46906 23044
rect 50246 23032 50252 23044
rect 46900 23004 50252 23032
rect 46900 22992 46906 23004
rect 50246 22992 50252 23004
rect 50304 22992 50310 23044
rect 50430 23041 50436 23044
rect 50424 23032 50436 23041
rect 50391 23004 50436 23032
rect 50424 22995 50436 23004
rect 50430 22992 50436 22995
rect 50488 22992 50494 23044
rect 52730 22992 52736 23044
rect 52788 23041 52794 23044
rect 52788 23032 52800 23041
rect 52788 23004 52833 23032
rect 52788 22995 52800 23004
rect 52788 22992 52794 22995
rect 53576 22976 53604 23072
rect 55950 23060 55956 23112
rect 56008 23060 56014 23112
rect 56962 23060 56968 23112
rect 57020 23060 57026 23112
rect 53736 23035 53794 23041
rect 53736 23001 53748 23035
rect 53782 23032 53794 23035
rect 53834 23032 53840 23044
rect 53782 23004 53840 23032
rect 53782 23001 53794 23004
rect 53736 22995 53794 23001
rect 53834 22992 53840 23004
rect 53892 22992 53898 23044
rect 57072 22976 57100 23140
rect 57793 23137 57805 23140
rect 57839 23137 57851 23171
rect 57793 23131 57851 23137
rect 57882 23128 57888 23180
rect 57940 23128 57946 23180
rect 57149 23103 57207 23109
rect 57149 23069 57161 23103
rect 57195 23100 57207 23103
rect 57701 23103 57759 23109
rect 57701 23100 57713 23103
rect 57195 23072 57713 23100
rect 57195 23069 57207 23072
rect 57149 23063 57207 23069
rect 57701 23069 57713 23072
rect 57747 23100 57759 23103
rect 57900 23100 57928 23128
rect 57747 23072 57928 23100
rect 57747 23069 57759 23072
rect 57701 23063 57759 23069
rect 43496 22936 44404 22964
rect 44545 22967 44603 22973
rect 43496 22924 43502 22936
rect 44545 22933 44557 22967
rect 44591 22964 44603 22967
rect 44726 22964 44732 22976
rect 44591 22936 44732 22964
rect 44591 22933 44603 22936
rect 44545 22927 44603 22933
rect 44726 22924 44732 22936
rect 44784 22924 44790 22976
rect 50614 22924 50620 22976
rect 50672 22964 50678 22976
rect 51810 22964 51816 22976
rect 50672 22936 51816 22964
rect 50672 22924 50678 22936
rect 51810 22924 51816 22936
rect 51868 22924 51874 22976
rect 53558 22924 53564 22976
rect 53616 22924 53622 22976
rect 55309 22967 55367 22973
rect 55309 22933 55321 22967
rect 55355 22964 55367 22967
rect 56686 22964 56692 22976
rect 55355 22936 56692 22964
rect 55355 22933 55367 22936
rect 55309 22927 55367 22933
rect 56686 22924 56692 22936
rect 56744 22924 56750 22976
rect 57054 22924 57060 22976
rect 57112 22924 57118 22976
rect 57609 22967 57667 22973
rect 57609 22933 57621 22967
rect 57655 22964 57667 22967
rect 57790 22964 57796 22976
rect 57655 22936 57796 22964
rect 57655 22933 57667 22936
rect 57609 22927 57667 22933
rect 57790 22924 57796 22936
rect 57848 22924 57854 22976
rect 1104 22874 59040 22896
rect 1104 22822 15394 22874
rect 15446 22822 15458 22874
rect 15510 22822 15522 22874
rect 15574 22822 15586 22874
rect 15638 22822 15650 22874
rect 15702 22822 29838 22874
rect 29890 22822 29902 22874
rect 29954 22822 29966 22874
rect 30018 22822 30030 22874
rect 30082 22822 30094 22874
rect 30146 22822 44282 22874
rect 44334 22822 44346 22874
rect 44398 22822 44410 22874
rect 44462 22822 44474 22874
rect 44526 22822 44538 22874
rect 44590 22822 58726 22874
rect 58778 22822 58790 22874
rect 58842 22822 58854 22874
rect 58906 22822 58918 22874
rect 58970 22822 58982 22874
rect 59034 22822 59040 22874
rect 1104 22800 59040 22822
rect 7558 22720 7564 22772
rect 7616 22760 7622 22772
rect 8297 22763 8355 22769
rect 8297 22760 8309 22763
rect 7616 22732 8309 22760
rect 7616 22720 7622 22732
rect 8297 22729 8309 22732
rect 8343 22729 8355 22763
rect 8297 22723 8355 22729
rect 13173 22763 13231 22769
rect 13173 22729 13185 22763
rect 13219 22760 13231 22763
rect 13538 22760 13544 22772
rect 13219 22732 13544 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 13630 22720 13636 22772
rect 13688 22720 13694 22772
rect 14921 22763 14979 22769
rect 14921 22729 14933 22763
rect 14967 22760 14979 22763
rect 15194 22760 15200 22772
rect 14967 22732 15200 22760
rect 14967 22729 14979 22732
rect 14921 22723 14979 22729
rect 15194 22720 15200 22732
rect 15252 22720 15258 22772
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 16025 22763 16083 22769
rect 16025 22760 16037 22763
rect 15896 22732 16037 22760
rect 15896 22720 15902 22732
rect 16025 22729 16037 22732
rect 16071 22729 16083 22763
rect 16025 22723 16083 22729
rect 16114 22720 16120 22772
rect 16172 22720 16178 22772
rect 16485 22763 16543 22769
rect 16485 22729 16497 22763
rect 16531 22760 16543 22763
rect 17402 22760 17408 22772
rect 16531 22732 17408 22760
rect 16531 22729 16543 22732
rect 16485 22723 16543 22729
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 17494 22720 17500 22772
rect 17552 22760 17558 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 17552 22732 17693 22760
rect 17552 22720 17558 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 17681 22723 17739 22729
rect 20165 22763 20223 22769
rect 20165 22729 20177 22763
rect 20211 22760 20223 22763
rect 20898 22760 20904 22772
rect 20211 22732 20904 22760
rect 20211 22729 20223 22732
rect 20165 22723 20223 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21821 22763 21879 22769
rect 21821 22729 21833 22763
rect 21867 22760 21879 22763
rect 22186 22760 22192 22772
rect 21867 22732 22192 22760
rect 21867 22729 21879 22732
rect 21821 22723 21879 22729
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 24912 22732 25360 22760
rect 24912 22720 24918 22732
rect 7742 22652 7748 22704
rect 7800 22692 7806 22704
rect 11701 22695 11759 22701
rect 11701 22692 11713 22695
rect 7800 22664 11713 22692
rect 7800 22652 7806 22664
rect 11701 22661 11713 22664
rect 11747 22692 11759 22695
rect 12250 22692 12256 22704
rect 11747 22664 12256 22692
rect 11747 22661 11759 22664
rect 11701 22655 11759 22661
rect 12250 22652 12256 22664
rect 12308 22652 12314 22704
rect 13648 22692 13676 22720
rect 19058 22701 19064 22704
rect 13556 22664 13676 22692
rect 15381 22695 15439 22701
rect 7650 22584 7656 22636
rect 7708 22624 7714 22636
rect 13556 22633 13584 22664
rect 15381 22661 15393 22695
rect 15427 22692 15439 22695
rect 19052 22692 19064 22701
rect 15427 22664 17540 22692
rect 19019 22664 19064 22692
rect 15427 22661 15439 22664
rect 15381 22655 15439 22661
rect 17512 22636 17540 22664
rect 19052 22655 19064 22664
rect 19058 22652 19064 22655
rect 19116 22652 19122 22704
rect 20714 22652 20720 22704
rect 20772 22692 20778 22704
rect 21726 22692 21732 22704
rect 20772 22664 21732 22692
rect 20772 22652 20778 22664
rect 21726 22652 21732 22664
rect 21784 22652 21790 22704
rect 22002 22652 22008 22704
rect 22060 22652 22066 22704
rect 25038 22692 25044 22704
rect 22480 22664 23244 22692
rect 8389 22627 8447 22633
rect 8389 22624 8401 22627
rect 7708 22596 8401 22624
rect 7708 22584 7714 22596
rect 8389 22593 8401 22596
rect 8435 22593 8447 22627
rect 8389 22587 8447 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22593 13599 22627
rect 13541 22587 13599 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22624 13691 22627
rect 14001 22627 14059 22633
rect 14001 22624 14013 22627
rect 13679 22596 14013 22624
rect 13679 22593 13691 22596
rect 13633 22587 13691 22593
rect 14001 22593 14013 22596
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 16114 22624 16120 22636
rect 15335 22596 16120 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 17494 22584 17500 22636
rect 17552 22584 17558 22636
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 17635 22596 18061 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 18782 22584 18788 22636
rect 18840 22584 18846 22636
rect 20162 22584 20168 22636
rect 20220 22624 20226 22636
rect 21177 22627 21235 22633
rect 21177 22624 21189 22627
rect 20220 22596 21189 22624
rect 20220 22584 20226 22596
rect 21177 22593 21189 22596
rect 21223 22593 21235 22627
rect 21177 22587 21235 22593
rect 21266 22584 21272 22636
rect 21324 22624 21330 22636
rect 22020 22624 22048 22652
rect 22480 22636 22508 22664
rect 21324 22596 22048 22624
rect 21324 22584 21330 22596
rect 22462 22584 22468 22636
rect 22520 22584 22526 22636
rect 22945 22627 23003 22633
rect 22945 22593 22957 22627
rect 22991 22624 23003 22627
rect 23106 22624 23112 22636
rect 22991 22596 23112 22624
rect 22991 22593 23003 22596
rect 22945 22587 23003 22593
rect 23106 22584 23112 22596
rect 23164 22584 23170 22636
rect 23216 22633 23244 22664
rect 23676 22664 25044 22692
rect 23676 22633 23704 22664
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 25332 22692 25360 22732
rect 25590 22720 25596 22772
rect 25648 22760 25654 22772
rect 25958 22760 25964 22772
rect 25648 22732 25964 22760
rect 25648 22720 25654 22732
rect 25958 22720 25964 22732
rect 26016 22720 26022 22772
rect 27249 22763 27307 22769
rect 27249 22729 27261 22763
rect 27295 22760 27307 22763
rect 27430 22760 27436 22772
rect 27295 22732 27436 22760
rect 27295 22729 27307 22732
rect 27249 22723 27307 22729
rect 27430 22720 27436 22732
rect 27488 22720 27494 22772
rect 27890 22720 27896 22772
rect 27948 22720 27954 22772
rect 29178 22720 29184 22772
rect 29236 22720 29242 22772
rect 29273 22763 29331 22769
rect 29273 22729 29285 22763
rect 29319 22760 29331 22763
rect 30558 22760 30564 22772
rect 29319 22732 30564 22760
rect 29319 22729 29331 22732
rect 29273 22723 29331 22729
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 31205 22763 31263 22769
rect 31205 22729 31217 22763
rect 31251 22760 31263 22763
rect 31570 22760 31576 22772
rect 31251 22732 31576 22760
rect 31251 22729 31263 22732
rect 31205 22723 31263 22729
rect 31570 22720 31576 22732
rect 31628 22720 31634 22772
rect 32861 22763 32919 22769
rect 32861 22729 32873 22763
rect 32907 22760 32919 22763
rect 34790 22760 34796 22772
rect 32907 22732 34796 22760
rect 32907 22729 32919 22732
rect 32861 22723 32919 22729
rect 34790 22720 34796 22732
rect 34848 22720 34854 22772
rect 35710 22760 35716 22772
rect 35084 22732 35716 22760
rect 26053 22695 26111 22701
rect 26053 22692 26065 22695
rect 25332 22664 26065 22692
rect 26053 22661 26065 22664
rect 26099 22661 26111 22695
rect 27908 22692 27936 22720
rect 28046 22695 28104 22701
rect 28046 22692 28058 22695
rect 27908 22664 28058 22692
rect 26053 22655 26111 22661
rect 28046 22661 28058 22664
rect 28092 22661 28104 22695
rect 28046 22655 28104 22661
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22624 23259 22627
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 23247 22596 23673 22624
rect 23247 22593 23259 22596
rect 23201 22587 23259 22593
rect 23661 22593 23673 22596
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 23928 22627 23986 22633
rect 23928 22593 23940 22627
rect 23974 22624 23986 22627
rect 24394 22624 24400 22636
rect 23974 22596 24400 22624
rect 23974 22593 23986 22596
rect 23928 22587 23986 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 26068 22624 26096 22655
rect 33134 22652 33140 22704
rect 33192 22692 33198 22704
rect 33192 22664 33548 22692
rect 33192 22652 33198 22664
rect 26418 22624 26424 22636
rect 26068 22596 26424 22624
rect 26418 22584 26424 22596
rect 26476 22624 26482 22636
rect 27522 22624 27528 22636
rect 26476 22596 27528 22624
rect 26476 22584 26482 22596
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27672 22596 27813 22624
rect 27672 22584 27678 22596
rect 27801 22593 27813 22596
rect 27847 22593 27859 22627
rect 31573 22627 31631 22633
rect 31573 22624 31585 22627
rect 27801 22587 27859 22593
rect 30760 22596 31585 22624
rect 5902 22516 5908 22568
rect 5960 22516 5966 22568
rect 8205 22559 8263 22565
rect 8205 22525 8217 22559
rect 8251 22556 8263 22559
rect 8570 22556 8576 22568
rect 8251 22528 8576 22556
rect 8251 22525 8263 22528
rect 8205 22519 8263 22525
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 9398 22516 9404 22568
rect 9456 22516 9462 22568
rect 10594 22516 10600 22568
rect 10652 22516 10658 22568
rect 11330 22516 11336 22568
rect 11388 22516 11394 22568
rect 11882 22516 11888 22568
rect 11940 22516 11946 22568
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22525 13783 22559
rect 13725 22519 13783 22525
rect 5261 22491 5319 22497
rect 5261 22457 5273 22491
rect 5307 22488 5319 22491
rect 5442 22488 5448 22500
rect 5307 22460 5448 22488
rect 5307 22457 5319 22460
rect 5261 22451 5319 22457
rect 5442 22448 5448 22460
rect 5500 22488 5506 22500
rect 7558 22488 7564 22500
rect 5500 22460 7564 22488
rect 5500 22448 5506 22460
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8757 22491 8815 22497
rect 8757 22457 8769 22491
rect 8803 22488 8815 22491
rect 9122 22488 9128 22500
rect 8803 22460 9128 22488
rect 8803 22457 8815 22460
rect 8757 22451 8815 22457
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 10612 22488 10640 22516
rect 13538 22488 13544 22500
rect 10612 22460 13544 22488
rect 13538 22448 13544 22460
rect 13596 22488 13602 22500
rect 13740 22488 13768 22519
rect 13906 22516 13912 22568
rect 13964 22556 13970 22568
rect 14553 22559 14611 22565
rect 14553 22556 14565 22559
rect 13964 22528 14565 22556
rect 13964 22516 13970 22528
rect 14553 22525 14565 22528
rect 14599 22525 14611 22559
rect 14553 22519 14611 22525
rect 14734 22516 14740 22568
rect 14792 22516 14798 22568
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22525 15531 22559
rect 15473 22519 15531 22525
rect 13596 22460 13768 22488
rect 14752 22488 14780 22516
rect 15488 22488 15516 22519
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 15620 22528 15853 22556
rect 15620 22516 15626 22528
rect 15841 22525 15853 22528
rect 15887 22525 15899 22559
rect 15841 22519 15899 22525
rect 17773 22559 17831 22565
rect 17773 22525 17785 22559
rect 17819 22525 17831 22559
rect 17773 22519 17831 22525
rect 14752 22460 15516 22488
rect 13596 22448 13602 22460
rect 17126 22448 17132 22500
rect 17184 22488 17190 22500
rect 17788 22488 17816 22519
rect 18598 22516 18604 22568
rect 18656 22516 18662 22568
rect 20806 22516 20812 22568
rect 20864 22556 20870 22568
rect 20993 22559 21051 22565
rect 20993 22556 21005 22559
rect 20864 22528 21005 22556
rect 20864 22516 20870 22528
rect 20993 22525 21005 22528
rect 21039 22525 21051 22559
rect 25774 22556 25780 22568
rect 20993 22519 21051 22525
rect 25516 22528 25780 22556
rect 17184 22460 17816 22488
rect 17184 22448 17190 22460
rect 5350 22380 5356 22432
rect 5408 22380 5414 22432
rect 6641 22423 6699 22429
rect 6641 22389 6653 22423
rect 6687 22420 6699 22423
rect 6914 22420 6920 22432
rect 6687 22392 6920 22420
rect 6687 22389 6699 22392
rect 6641 22383 6699 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 8846 22380 8852 22432
rect 8904 22380 8910 22432
rect 10686 22380 10692 22432
rect 10744 22380 10750 22432
rect 12526 22380 12532 22432
rect 12584 22380 12590 22432
rect 17221 22423 17279 22429
rect 17221 22389 17233 22423
rect 17267 22420 17279 22423
rect 17402 22420 17408 22432
rect 17267 22392 17408 22420
rect 17267 22389 17279 22392
rect 17221 22383 17279 22389
rect 17402 22380 17408 22392
rect 17460 22380 17466 22432
rect 21008 22420 21036 22519
rect 21637 22491 21695 22497
rect 21637 22457 21649 22491
rect 21683 22488 21695 22491
rect 22186 22488 22192 22500
rect 21683 22460 22192 22488
rect 21683 22457 21695 22460
rect 21637 22451 21695 22457
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 25516 22497 25544 22528
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 29730 22516 29736 22568
rect 29788 22556 29794 22568
rect 30098 22565 30104 22568
rect 29917 22559 29975 22565
rect 29917 22556 29929 22559
rect 29788 22528 29929 22556
rect 29788 22516 29794 22528
rect 29917 22525 29929 22528
rect 29963 22525 29975 22559
rect 29917 22519 29975 22525
rect 30076 22559 30104 22565
rect 30076 22525 30088 22559
rect 30076 22519 30104 22525
rect 30098 22516 30104 22519
rect 30156 22516 30162 22568
rect 30193 22559 30251 22565
rect 30193 22525 30205 22559
rect 30239 22556 30251 22559
rect 30558 22556 30564 22568
rect 30239 22528 30564 22556
rect 30239 22525 30251 22528
rect 30193 22519 30251 22525
rect 30558 22516 30564 22528
rect 30616 22516 30622 22568
rect 25501 22491 25559 22497
rect 25501 22488 25513 22491
rect 24596 22460 25513 22488
rect 24596 22420 24624 22460
rect 25501 22457 25513 22460
rect 25547 22457 25559 22491
rect 25501 22451 25559 22457
rect 26421 22491 26479 22497
rect 26421 22457 26433 22491
rect 26467 22488 26479 22491
rect 26467 22460 27292 22488
rect 26467 22457 26479 22460
rect 26421 22451 26479 22457
rect 21008 22392 24624 22420
rect 24946 22380 24952 22432
rect 25004 22420 25010 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 25004 22392 25053 22420
rect 25004 22380 25010 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 27264 22420 27292 22460
rect 29086 22448 29092 22500
rect 29144 22448 29150 22500
rect 30469 22491 30527 22497
rect 30469 22457 30481 22491
rect 30515 22488 30527 22491
rect 30650 22488 30656 22500
rect 30515 22460 30656 22488
rect 30515 22457 30527 22460
rect 30469 22451 30527 22457
rect 30650 22448 30656 22460
rect 30708 22448 30714 22500
rect 27982 22420 27988 22432
rect 27264 22392 27988 22420
rect 25041 22383 25099 22389
rect 27982 22380 27988 22392
rect 28040 22380 28046 22432
rect 29104 22420 29132 22448
rect 30760 22420 30788 22596
rect 31573 22593 31585 22596
rect 31619 22593 31631 22627
rect 31573 22587 31631 22593
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22624 31723 22627
rect 32769 22627 32827 22633
rect 31711 22596 32168 22624
rect 31711 22593 31723 22596
rect 31665 22587 31723 22593
rect 30926 22516 30932 22568
rect 30984 22516 30990 22568
rect 31113 22559 31171 22565
rect 31113 22525 31125 22559
rect 31159 22556 31171 22559
rect 31680 22556 31708 22587
rect 32140 22568 32168 22596
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 33410 22624 33416 22636
rect 32815 22596 33416 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 31159 22528 31708 22556
rect 31757 22559 31815 22565
rect 31159 22525 31171 22528
rect 31113 22519 31171 22525
rect 31757 22525 31769 22559
rect 31803 22525 31815 22559
rect 31757 22519 31815 22525
rect 31386 22448 31392 22500
rect 31444 22488 31450 22500
rect 31772 22488 31800 22519
rect 32122 22516 32128 22568
rect 32180 22516 32186 22568
rect 33042 22516 33048 22568
rect 33100 22516 33106 22568
rect 33520 22556 33548 22664
rect 34330 22584 34336 22636
rect 34388 22584 34394 22636
rect 35084 22633 35112 22732
rect 35710 22720 35716 22732
rect 35768 22720 35774 22772
rect 36170 22720 36176 22772
rect 36228 22720 36234 22772
rect 40221 22763 40279 22769
rect 40221 22729 40233 22763
rect 40267 22760 40279 22763
rect 41598 22760 41604 22772
rect 40267 22732 41604 22760
rect 40267 22729 40279 22732
rect 40221 22723 40279 22729
rect 41598 22720 41604 22732
rect 41656 22720 41662 22772
rect 42334 22720 42340 22772
rect 42392 22760 42398 22772
rect 42429 22763 42487 22769
rect 42429 22760 42441 22763
rect 42392 22732 42441 22760
rect 42392 22720 42398 22732
rect 42429 22729 42441 22732
rect 42475 22729 42487 22763
rect 42429 22723 42487 22729
rect 42886 22720 42892 22772
rect 42944 22720 42950 22772
rect 43257 22763 43315 22769
rect 43257 22729 43269 22763
rect 43303 22760 43315 22763
rect 43990 22760 43996 22772
rect 43303 22732 43996 22760
rect 43303 22729 43315 22732
rect 43257 22723 43315 22729
rect 43990 22720 43996 22732
rect 44048 22720 44054 22772
rect 48774 22760 48780 22772
rect 47044 22732 48780 22760
rect 35802 22652 35808 22704
rect 35860 22692 35866 22704
rect 41414 22692 41420 22704
rect 35860 22664 35940 22692
rect 35860 22652 35866 22664
rect 35069 22627 35127 22633
rect 35069 22593 35081 22627
rect 35115 22593 35127 22627
rect 35069 22587 35127 22593
rect 35176 22596 35480 22624
rect 34054 22556 34060 22568
rect 33520 22528 34060 22556
rect 34054 22516 34060 22528
rect 34112 22516 34118 22568
rect 34146 22516 34152 22568
rect 34204 22565 34210 22568
rect 34204 22559 34253 22565
rect 34204 22525 34207 22559
rect 34241 22525 34253 22559
rect 34204 22519 34253 22525
rect 34204 22516 34210 22519
rect 34606 22516 34612 22568
rect 34664 22516 34670 22568
rect 35176 22556 35204 22596
rect 34808 22528 35204 22556
rect 34808 22500 34836 22528
rect 35250 22516 35256 22568
rect 35308 22516 35314 22568
rect 35452 22556 35480 22596
rect 35912 22565 35940 22664
rect 38856 22664 41420 22692
rect 37544 22627 37602 22633
rect 37544 22593 37556 22627
rect 37590 22624 37602 22627
rect 38010 22624 38016 22636
rect 37590 22596 38016 22624
rect 37590 22593 37602 22596
rect 37544 22587 37602 22593
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 38654 22584 38660 22636
rect 38712 22624 38718 22636
rect 38856 22633 38884 22664
rect 38841 22627 38899 22633
rect 38841 22624 38853 22627
rect 38712 22596 38853 22624
rect 38712 22584 38718 22596
rect 38841 22593 38853 22596
rect 38887 22593 38899 22627
rect 38841 22587 38899 22593
rect 39108 22627 39166 22633
rect 39108 22593 39120 22627
rect 39154 22624 39166 22627
rect 40586 22624 40592 22636
rect 39154 22596 40592 22624
rect 39154 22593 39166 22596
rect 39108 22587 39166 22593
rect 40586 22584 40592 22596
rect 40644 22584 40650 22636
rect 40880 22633 40908 22664
rect 41414 22652 41420 22664
rect 41472 22692 41478 22704
rect 42518 22692 42524 22704
rect 41472 22664 42524 22692
rect 41472 22652 41478 22664
rect 42518 22652 42524 22664
rect 42576 22652 42582 22704
rect 42797 22695 42855 22701
rect 42797 22661 42809 22695
rect 42843 22692 42855 22695
rect 43714 22692 43720 22704
rect 42843 22664 43720 22692
rect 42843 22661 42855 22664
rect 42797 22655 42855 22661
rect 43714 22652 43720 22664
rect 43772 22652 43778 22704
rect 44174 22652 44180 22704
rect 44232 22652 44238 22704
rect 44392 22695 44450 22701
rect 44392 22661 44404 22695
rect 44438 22692 44450 22695
rect 45094 22692 45100 22704
rect 44438 22664 45100 22692
rect 44438 22661 44450 22664
rect 44392 22655 44450 22661
rect 45094 22652 45100 22664
rect 45152 22652 45158 22704
rect 45373 22695 45431 22701
rect 45373 22661 45385 22695
rect 45419 22692 45431 22695
rect 45554 22692 45560 22704
rect 45419 22664 45560 22692
rect 45419 22661 45431 22664
rect 45373 22655 45431 22661
rect 45554 22652 45560 22664
rect 45612 22692 45618 22704
rect 45833 22695 45891 22701
rect 45833 22692 45845 22695
rect 45612 22664 45845 22692
rect 45612 22652 45618 22664
rect 45833 22661 45845 22664
rect 45879 22692 45891 22695
rect 47044 22692 47072 22732
rect 48774 22720 48780 22732
rect 48832 22720 48838 22772
rect 50433 22763 50491 22769
rect 50433 22729 50445 22763
rect 50479 22760 50491 22763
rect 50614 22760 50620 22772
rect 50479 22732 50620 22760
rect 50479 22729 50491 22732
rect 50433 22723 50491 22729
rect 50614 22720 50620 22732
rect 50672 22720 50678 22772
rect 50709 22763 50767 22769
rect 50709 22729 50721 22763
rect 50755 22760 50767 22763
rect 51994 22760 52000 22772
rect 50755 22732 52000 22760
rect 50755 22729 50767 22732
rect 50709 22723 50767 22729
rect 51994 22720 52000 22732
rect 52052 22720 52058 22772
rect 53098 22720 53104 22772
rect 53156 22720 53162 22772
rect 53190 22720 53196 22772
rect 53248 22720 53254 22772
rect 55766 22720 55772 22772
rect 55824 22720 55830 22772
rect 57606 22720 57612 22772
rect 57664 22720 57670 22772
rect 45879 22664 47072 22692
rect 45879 22661 45891 22664
rect 45833 22655 45891 22661
rect 53558 22652 53564 22704
rect 53616 22692 53622 22704
rect 56496 22695 56554 22701
rect 53616 22664 56272 22692
rect 53616 22652 53622 22664
rect 40865 22627 40923 22633
rect 40865 22593 40877 22627
rect 40911 22593 40923 22627
rect 40865 22587 40923 22593
rect 41132 22627 41190 22633
rect 41132 22593 41144 22627
rect 41178 22624 41190 22627
rect 41690 22624 41696 22636
rect 41178 22596 41696 22624
rect 41178 22593 41190 22596
rect 41132 22587 41190 22593
rect 41690 22584 41696 22596
rect 41748 22584 41754 22636
rect 44192 22624 44220 22652
rect 43180 22596 44220 22624
rect 43180 22568 43208 22596
rect 44634 22584 44640 22636
rect 44692 22624 44698 22636
rect 45462 22624 45468 22636
rect 44692 22596 45468 22624
rect 44692 22584 44698 22596
rect 45462 22584 45468 22596
rect 45520 22624 45526 22636
rect 46198 22633 46204 22636
rect 45925 22627 45983 22633
rect 45925 22624 45937 22627
rect 45520 22596 45937 22624
rect 45520 22584 45526 22596
rect 45925 22593 45937 22596
rect 45971 22593 45983 22627
rect 45925 22587 45983 22593
rect 46192 22587 46204 22633
rect 46198 22584 46204 22587
rect 46256 22584 46262 22636
rect 46934 22584 46940 22636
rect 46992 22584 46998 22636
rect 48314 22584 48320 22636
rect 48372 22633 48378 22636
rect 48372 22627 48421 22633
rect 48372 22593 48375 22627
rect 48409 22593 48421 22627
rect 48372 22587 48421 22593
rect 48372 22584 48378 22587
rect 49050 22584 49056 22636
rect 49108 22624 49114 22636
rect 49421 22627 49479 22633
rect 49421 22624 49433 22627
rect 49108 22596 49433 22624
rect 49108 22584 49114 22596
rect 49421 22593 49433 22596
rect 49467 22593 49479 22627
rect 49421 22587 49479 22593
rect 51353 22627 51411 22633
rect 51353 22593 51365 22627
rect 51399 22593 51411 22627
rect 51353 22587 51411 22593
rect 35805 22559 35863 22565
rect 35805 22556 35817 22559
rect 35452 22528 35817 22556
rect 35805 22525 35817 22528
rect 35851 22525 35863 22559
rect 35805 22519 35863 22525
rect 35897 22559 35955 22565
rect 35897 22525 35909 22559
rect 35943 22525 35955 22559
rect 35897 22519 35955 22525
rect 36722 22516 36728 22568
rect 36780 22516 36786 22568
rect 36906 22516 36912 22568
rect 36964 22556 36970 22568
rect 37277 22559 37335 22565
rect 37277 22556 37289 22559
rect 36964 22528 37289 22556
rect 36964 22516 36970 22528
rect 37277 22525 37289 22528
rect 37323 22525 37335 22559
rect 37277 22519 37335 22525
rect 43073 22559 43131 22565
rect 43073 22525 43085 22559
rect 43119 22556 43131 22559
rect 43162 22556 43168 22568
rect 43119 22528 43168 22556
rect 43119 22525 43131 22528
rect 43073 22519 43131 22525
rect 43162 22516 43168 22528
rect 43220 22516 43226 22568
rect 44910 22516 44916 22568
rect 44968 22516 44974 22568
rect 46952 22556 46980 22584
rect 48225 22559 48283 22565
rect 48225 22556 48237 22559
rect 46952 22528 48237 22556
rect 31444 22460 31800 22488
rect 31444 22448 31450 22460
rect 34790 22448 34796 22500
rect 34848 22448 34854 22500
rect 35345 22491 35403 22497
rect 35345 22457 35357 22491
rect 35391 22488 35403 22491
rect 35986 22488 35992 22500
rect 35391 22460 35992 22488
rect 35391 22457 35403 22460
rect 35345 22451 35403 22457
rect 35986 22448 35992 22460
rect 36044 22448 36050 22500
rect 29104 22392 30788 22420
rect 32398 22380 32404 22432
rect 32456 22380 32462 22432
rect 33413 22423 33471 22429
rect 33413 22389 33425 22423
rect 33459 22420 33471 22423
rect 35526 22420 35532 22432
rect 33459 22392 35532 22420
rect 33459 22389 33471 22392
rect 33413 22383 33471 22389
rect 35526 22380 35532 22392
rect 35584 22380 35590 22432
rect 38654 22380 38660 22432
rect 38712 22380 38718 22432
rect 42242 22380 42248 22432
rect 42300 22380 42306 22432
rect 42610 22380 42616 22432
rect 42668 22420 42674 22432
rect 44928 22420 44956 22516
rect 42668 22392 44956 22420
rect 42668 22380 42674 22392
rect 45002 22380 45008 22432
rect 45060 22420 45066 22432
rect 46952 22420 46980 22528
rect 48225 22525 48237 22528
rect 48271 22525 48283 22559
rect 48225 22519 48283 22525
rect 48501 22559 48559 22565
rect 48501 22525 48513 22559
rect 48547 22556 48559 22559
rect 48547 22528 48728 22556
rect 48547 22525 48559 22528
rect 48501 22519 48559 22525
rect 45060 22392 46980 22420
rect 45060 22380 45066 22392
rect 47302 22380 47308 22432
rect 47360 22380 47366 22432
rect 47578 22380 47584 22432
rect 47636 22380 47642 22432
rect 48222 22380 48228 22432
rect 48280 22420 48286 22432
rect 48700 22420 48728 22528
rect 49234 22516 49240 22568
rect 49292 22516 49298 22568
rect 51166 22516 51172 22568
rect 51224 22556 51230 22568
rect 51368 22556 51396 22587
rect 51626 22584 51632 22636
rect 51684 22584 51690 22636
rect 52454 22584 52460 22636
rect 52512 22624 52518 22636
rect 53668 22633 53696 22664
rect 52549 22627 52607 22633
rect 52549 22624 52561 22627
rect 52512 22596 52561 22624
rect 52512 22584 52518 22596
rect 52549 22593 52561 22596
rect 52595 22593 52607 22627
rect 52549 22587 52607 22593
rect 53653 22627 53711 22633
rect 53653 22593 53665 22627
rect 53699 22593 53711 22627
rect 53653 22587 53711 22593
rect 53920 22627 53978 22633
rect 53920 22593 53932 22627
rect 53966 22624 53978 22627
rect 55490 22624 55496 22636
rect 53966 22596 55496 22624
rect 53966 22593 53978 22596
rect 53920 22587 53978 22593
rect 55490 22584 55496 22596
rect 55548 22584 55554 22636
rect 56244 22633 56272 22664
rect 56496 22661 56508 22695
rect 56542 22692 56554 22695
rect 57330 22692 57336 22704
rect 56542 22664 57336 22692
rect 56542 22661 56554 22664
rect 56496 22655 56554 22661
rect 57330 22652 57336 22664
rect 57388 22652 57394 22704
rect 56229 22627 56287 22633
rect 56229 22593 56241 22627
rect 56275 22624 56287 22627
rect 56318 22624 56324 22636
rect 56275 22596 56324 22624
rect 56275 22593 56287 22596
rect 56229 22587 56287 22593
rect 56318 22584 56324 22596
rect 56376 22584 56382 22636
rect 58066 22584 58072 22636
rect 58124 22624 58130 22636
rect 58437 22627 58495 22633
rect 58437 22624 58449 22627
rect 58124 22596 58449 22624
rect 58124 22584 58130 22596
rect 58437 22593 58449 22596
rect 58483 22593 58495 22627
rect 58437 22587 58495 22593
rect 51224 22528 51396 22556
rect 51224 22516 51230 22528
rect 51442 22516 51448 22568
rect 51500 22565 51506 22568
rect 51500 22559 51549 22565
rect 51500 22525 51503 22559
rect 51537 22525 51549 22559
rect 51500 22519 51549 22525
rect 51500 22516 51506 22519
rect 52362 22516 52368 22568
rect 52420 22516 52426 22568
rect 52638 22516 52644 22568
rect 52696 22556 52702 22568
rect 53285 22559 53343 22565
rect 53285 22556 53297 22559
rect 52696 22528 53297 22556
rect 52696 22516 52702 22528
rect 53285 22525 53297 22528
rect 53331 22525 53343 22559
rect 53285 22519 53343 22525
rect 55125 22559 55183 22565
rect 55125 22525 55137 22559
rect 55171 22525 55183 22559
rect 55125 22519 55183 22525
rect 48774 22448 48780 22500
rect 48832 22488 48838 22500
rect 49602 22488 49608 22500
rect 48832 22460 49608 22488
rect 48832 22448 48838 22460
rect 49602 22448 49608 22460
rect 49660 22448 49666 22500
rect 51810 22448 51816 22500
rect 51868 22488 51874 22500
rect 51905 22491 51963 22497
rect 51905 22488 51917 22491
rect 51868 22460 51917 22488
rect 51868 22448 51874 22460
rect 51905 22457 51917 22460
rect 51951 22457 51963 22491
rect 51905 22451 51963 22457
rect 55033 22491 55091 22497
rect 55033 22457 55045 22491
rect 55079 22488 55091 22491
rect 55140 22488 55168 22519
rect 55079 22460 55168 22488
rect 55079 22457 55091 22460
rect 55033 22451 55091 22457
rect 48280 22392 48728 22420
rect 49789 22423 49847 22429
rect 48280 22380 48286 22392
rect 49789 22389 49801 22423
rect 49835 22420 49847 22423
rect 51166 22420 51172 22432
rect 49835 22392 51172 22420
rect 49835 22389 49847 22392
rect 49789 22383 49847 22389
rect 51166 22380 51172 22392
rect 51224 22380 51230 22432
rect 52730 22380 52736 22432
rect 52788 22380 52794 22432
rect 56962 22380 56968 22432
rect 57020 22420 57026 22432
rect 57885 22423 57943 22429
rect 57885 22420 57897 22423
rect 57020 22392 57897 22420
rect 57020 22380 57026 22392
rect 57885 22389 57897 22392
rect 57931 22389 57943 22423
rect 57885 22383 57943 22389
rect 1104 22330 58880 22352
rect 1104 22278 8172 22330
rect 8224 22278 8236 22330
rect 8288 22278 8300 22330
rect 8352 22278 8364 22330
rect 8416 22278 8428 22330
rect 8480 22278 22616 22330
rect 22668 22278 22680 22330
rect 22732 22278 22744 22330
rect 22796 22278 22808 22330
rect 22860 22278 22872 22330
rect 22924 22278 37060 22330
rect 37112 22278 37124 22330
rect 37176 22278 37188 22330
rect 37240 22278 37252 22330
rect 37304 22278 37316 22330
rect 37368 22278 51504 22330
rect 51556 22278 51568 22330
rect 51620 22278 51632 22330
rect 51684 22278 51696 22330
rect 51748 22278 51760 22330
rect 51812 22278 58880 22330
rect 1104 22256 58880 22278
rect 5442 22176 5448 22228
rect 5500 22176 5506 22228
rect 5629 22219 5687 22225
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5902 22216 5908 22228
rect 5675 22188 5908 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5902 22176 5908 22188
rect 5960 22176 5966 22228
rect 8941 22219 8999 22225
rect 8941 22185 8953 22219
rect 8987 22216 8999 22219
rect 9398 22216 9404 22228
rect 8987 22188 9404 22216
rect 8987 22185 8999 22188
rect 8941 22179 8999 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 11330 22176 11336 22228
rect 11388 22176 11394 22228
rect 11609 22219 11667 22225
rect 11609 22185 11621 22219
rect 11655 22216 11667 22219
rect 11882 22216 11888 22228
rect 11655 22188 11888 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 12250 22176 12256 22228
rect 12308 22216 12314 22228
rect 12308 22188 13492 22216
rect 12308 22176 12314 22188
rect 5460 22089 5488 22176
rect 6914 22148 6920 22160
rect 6288 22120 6920 22148
rect 5445 22083 5503 22089
rect 5445 22049 5457 22083
rect 5491 22049 5503 22083
rect 5445 22043 5503 22049
rect 6181 22083 6239 22089
rect 6181 22049 6193 22083
rect 6227 22080 6239 22083
rect 6288 22080 6316 22120
rect 6914 22108 6920 22120
rect 6972 22148 6978 22160
rect 7742 22148 7748 22160
rect 6972 22120 7748 22148
rect 6972 22108 6978 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 11348 22148 11376 22176
rect 11701 22151 11759 22157
rect 11701 22148 11713 22151
rect 9508 22120 10088 22148
rect 11348 22120 11713 22148
rect 8846 22080 8852 22092
rect 6227 22052 6316 22080
rect 8680 22052 8852 22080
rect 6227 22049 6239 22052
rect 6181 22043 6239 22049
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 8501 22015 8559 22021
rect 8501 21981 8513 22015
rect 8547 22012 8559 22015
rect 8680 22012 8708 22052
rect 8846 22040 8852 22052
rect 8904 22040 8910 22092
rect 8547 21984 8708 22012
rect 8757 22015 8815 22021
rect 8547 21981 8559 21984
rect 8501 21975 8559 21981
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 9508 22012 9536 22120
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 9631 22052 9996 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 9674 22012 9680 22024
rect 8803 21984 9680 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 5166 21904 5172 21956
rect 5224 21944 5230 21956
rect 7190 21944 7196 21956
rect 5224 21916 7196 21944
rect 5224 21904 5230 21916
rect 7190 21904 7196 21916
rect 7248 21904 7254 21956
rect 7466 21904 7472 21956
rect 7524 21944 7530 21956
rect 9309 21947 9367 21953
rect 9309 21944 9321 21947
rect 7524 21916 9321 21944
rect 7524 21904 7530 21916
rect 9309 21913 9321 21916
rect 9355 21913 9367 21947
rect 9968 21944 9996 22052
rect 10060 22012 10088 22120
rect 11701 22117 11713 22120
rect 11747 22117 11759 22151
rect 11701 22111 11759 22117
rect 12268 22089 12296 22176
rect 13464 22148 13492 22188
rect 13906 22176 13912 22228
rect 13964 22176 13970 22228
rect 14734 22176 14740 22228
rect 14792 22216 14798 22228
rect 16390 22216 16396 22228
rect 14792 22188 16396 22216
rect 14792 22176 14798 22188
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 17126 22176 17132 22228
rect 17184 22216 17190 22228
rect 17586 22216 17592 22228
rect 17184 22188 17592 22216
rect 17184 22176 17190 22188
rect 17586 22176 17592 22188
rect 17644 22176 17650 22228
rect 18049 22219 18107 22225
rect 18049 22185 18061 22219
rect 18095 22216 18107 22219
rect 18598 22216 18604 22228
rect 18095 22188 18604 22216
rect 18095 22185 18107 22188
rect 18049 22179 18107 22185
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 20162 22176 20168 22228
rect 20220 22176 20226 22228
rect 21174 22216 21180 22228
rect 20732 22188 21180 22216
rect 13464 22120 14412 22148
rect 12253 22083 12311 22089
rect 12253 22049 12265 22083
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 13630 22040 13636 22092
rect 13688 22080 13694 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 13688 22052 14289 22080
rect 13688 22040 13694 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14384 22080 14412 22120
rect 14734 22080 14740 22092
rect 14384 22052 14740 22080
rect 14277 22043 14335 22049
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10060 21984 10241 22012
rect 10229 21981 10241 21984
rect 10275 22012 10287 22015
rect 10318 22012 10324 22024
rect 10275 21984 10324 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10318 21972 10324 21984
rect 10376 22012 10382 22024
rect 12434 22012 12440 22024
rect 10376 21984 12440 22012
rect 10376 21972 10382 21984
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 12802 22021 12808 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12492 21984 12541 22012
rect 12492 21972 12498 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 12796 21975 12808 22021
rect 12802 21972 12808 21975
rect 12860 21972 12866 22024
rect 14292 22012 14320 22043
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 15838 22040 15844 22092
rect 15896 22080 15902 22092
rect 16209 22083 16267 22089
rect 16209 22080 16221 22083
rect 15896 22052 16221 22080
rect 15896 22040 15902 22052
rect 16209 22049 16221 22052
rect 16255 22049 16267 22083
rect 16209 22043 16267 22049
rect 16316 22080 16712 22094
rect 16853 22083 16911 22089
rect 16853 22080 16865 22083
rect 16316 22066 16865 22080
rect 15562 22012 15568 22024
rect 14292 21984 15568 22012
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 10496 21947 10554 21953
rect 9968 21916 10088 21944
rect 9309 21907 9367 21913
rect 4798 21836 4804 21888
rect 4856 21836 4862 21888
rect 5261 21879 5319 21885
rect 5261 21845 5273 21879
rect 5307 21876 5319 21879
rect 5534 21876 5540 21888
rect 5307 21848 5540 21876
rect 5307 21845 5319 21848
rect 5261 21839 5319 21845
rect 5534 21836 5540 21848
rect 5592 21876 5598 21888
rect 5994 21876 6000 21888
rect 5592 21848 6000 21876
rect 5592 21836 5598 21848
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6089 21879 6147 21885
rect 6089 21845 6101 21879
rect 6135 21876 6147 21879
rect 7101 21879 7159 21885
rect 7101 21876 7113 21879
rect 6135 21848 7113 21876
rect 6135 21845 6147 21848
rect 6089 21839 6147 21845
rect 7101 21845 7113 21848
rect 7147 21876 7159 21879
rect 7282 21876 7288 21888
rect 7147 21848 7288 21876
rect 7147 21845 7159 21848
rect 7101 21839 7159 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 7377 21879 7435 21885
rect 7377 21845 7389 21879
rect 7423 21876 7435 21879
rect 8294 21876 8300 21888
rect 7423 21848 8300 21876
rect 7423 21845 7435 21848
rect 7377 21839 7435 21845
rect 8294 21836 8300 21848
rect 8352 21836 8358 21888
rect 9398 21836 9404 21888
rect 9456 21836 9462 21888
rect 10060 21885 10088 21916
rect 10496 21913 10508 21947
rect 10542 21944 10554 21947
rect 10686 21944 10692 21956
rect 10542 21916 10692 21944
rect 10542 21913 10554 21916
rect 10496 21907 10554 21913
rect 10686 21904 10692 21916
rect 10744 21904 10750 21956
rect 13722 21944 13728 21956
rect 12084 21916 13728 21944
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 10594 21876 10600 21888
rect 10091 21848 10600 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 12084 21885 12112 21916
rect 13722 21904 13728 21916
rect 13780 21904 13786 21956
rect 16316 21888 16344 22066
rect 16684 22052 16865 22066
rect 16853 22049 16865 22052
rect 16899 22049 16911 22083
rect 16853 22043 16911 22049
rect 17126 22040 17132 22092
rect 17184 22040 17190 22092
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22080 17463 22083
rect 17451 22052 18460 22080
rect 17451 22049 17463 22052
rect 17405 22043 17463 22049
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 16574 22012 16580 22024
rect 16439 21984 16580 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17218 21972 17224 22024
rect 17276 22021 17282 22024
rect 17276 22015 17304 22021
rect 17292 21981 17304 22015
rect 17276 21975 17304 21981
rect 17276 21972 17282 21975
rect 12069 21879 12127 21885
rect 12069 21876 12081 21879
rect 11112 21848 12081 21876
rect 11112 21836 11118 21848
rect 12069 21845 12081 21848
rect 12115 21845 12127 21879
rect 12069 21839 12127 21845
rect 12161 21879 12219 21885
rect 12161 21845 12173 21879
rect 12207 21876 12219 21879
rect 12526 21876 12532 21888
rect 12207 21848 12532 21876
rect 12207 21845 12219 21848
rect 12161 21839 12219 21845
rect 12526 21836 12532 21848
rect 12584 21876 12590 21888
rect 12986 21876 12992 21888
rect 12584 21848 12992 21876
rect 12584 21836 12590 21848
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 16298 21876 16304 21888
rect 16163 21848 16304 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 18432 21885 18460 22052
rect 20622 21944 20628 21956
rect 19812 21916 20628 21944
rect 19812 21888 19840 21916
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 18417 21879 18475 21885
rect 18417 21876 18429 21879
rect 17368 21848 18429 21876
rect 17368 21836 17374 21848
rect 18417 21845 18429 21848
rect 18463 21876 18475 21879
rect 19794 21876 19800 21888
rect 18463 21848 19800 21876
rect 18463 21845 18475 21848
rect 18417 21839 18475 21845
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 19944 21848 20085 21876
rect 19944 21836 19950 21848
rect 20073 21845 20085 21848
rect 20119 21876 20131 21879
rect 20438 21876 20444 21888
rect 20119 21848 20444 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20438 21836 20444 21848
rect 20496 21876 20502 21888
rect 20732 21876 20760 22188
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 25774 22176 25780 22228
rect 25832 22216 25838 22228
rect 57054 22216 57060 22228
rect 25832 22188 57060 22216
rect 25832 22176 25838 22188
rect 57054 22176 57060 22188
rect 57112 22176 57118 22228
rect 26326 22148 26332 22160
rect 26206 22120 26332 22148
rect 22281 22083 22339 22089
rect 22281 22049 22293 22083
rect 22327 22080 22339 22083
rect 22462 22080 22468 22092
rect 22327 22052 22468 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 22925 22083 22983 22089
rect 22925 22049 22937 22083
rect 22971 22049 22983 22083
rect 26206 22080 26234 22120
rect 26326 22108 26332 22120
rect 26384 22148 26390 22160
rect 26970 22148 26976 22160
rect 26384 22120 26976 22148
rect 26384 22108 26390 22120
rect 26970 22108 26976 22120
rect 27028 22108 27034 22160
rect 31205 22151 31263 22157
rect 31205 22117 31217 22151
rect 31251 22117 31263 22151
rect 31205 22111 31263 22117
rect 22925 22043 22983 22049
rect 25332 22052 26234 22080
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 20496 21848 20760 21876
rect 20824 21876 20852 21975
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22940 22012 22968 22043
rect 22244 21984 22968 22012
rect 22244 21972 22250 21984
rect 22036 21947 22094 21953
rect 22036 21913 22048 21947
rect 22082 21944 22094 21947
rect 22373 21947 22431 21953
rect 22373 21944 22385 21947
rect 22082 21916 22385 21944
rect 22082 21913 22094 21916
rect 22036 21907 22094 21913
rect 22373 21913 22385 21916
rect 22419 21913 22431 21947
rect 22373 21907 22431 21913
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20824 21848 20913 21876
rect 20496 21836 20502 21848
rect 20901 21845 20913 21848
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24912 21848 24961 21876
rect 24912 21836 24918 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25332 21885 25360 22052
rect 27798 22040 27804 22092
rect 27856 22040 27862 22092
rect 28902 22040 28908 22092
rect 28960 22080 28966 22092
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 28960 22052 29837 22080
rect 28960 22040 28966 22052
rect 29825 22049 29837 22052
rect 29871 22049 29883 22083
rect 31220 22080 31248 22111
rect 32122 22108 32128 22160
rect 32180 22108 32186 22160
rect 32306 22108 32312 22160
rect 32364 22108 32370 22160
rect 33410 22108 33416 22160
rect 33468 22148 33474 22160
rect 33781 22151 33839 22157
rect 33781 22148 33793 22151
rect 33468 22120 33793 22148
rect 33468 22108 33474 22120
rect 33781 22117 33793 22120
rect 33827 22148 33839 22151
rect 34146 22148 34152 22160
rect 33827 22120 34152 22148
rect 33827 22117 33839 22120
rect 33781 22111 33839 22117
rect 34146 22108 34152 22120
rect 34204 22108 34210 22160
rect 35250 22148 35256 22160
rect 34716 22120 34928 22148
rect 31481 22083 31539 22089
rect 31481 22080 31493 22083
rect 31220 22052 31493 22080
rect 29825 22043 29883 22049
rect 31481 22049 31493 22052
rect 31527 22049 31539 22083
rect 31481 22043 31539 22049
rect 32398 22040 32404 22092
rect 32456 22080 32462 22092
rect 32861 22083 32919 22089
rect 32861 22080 32873 22083
rect 32456 22052 32873 22080
rect 32456 22040 32462 22052
rect 32861 22049 32873 22052
rect 32907 22049 32919 22083
rect 32861 22043 32919 22049
rect 33042 22040 33048 22092
rect 33100 22040 33106 22092
rect 33229 22083 33287 22089
rect 33229 22049 33241 22083
rect 33275 22080 33287 22083
rect 33318 22080 33324 22092
rect 33275 22052 33324 22080
rect 33275 22049 33287 22052
rect 33229 22043 33287 22049
rect 33318 22040 33324 22052
rect 33376 22040 33382 22092
rect 34716 22080 34744 22120
rect 34440 22052 34744 22080
rect 34793 22083 34851 22089
rect 30092 22015 30150 22021
rect 30092 21981 30104 22015
rect 30138 22012 30150 22015
rect 31018 22012 31024 22024
rect 30138 21984 31024 22012
rect 30138 21981 30150 21984
rect 30092 21975 30150 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 33060 22012 33088 22040
rect 34440 22012 34468 22052
rect 34793 22049 34805 22083
rect 34839 22049 34851 22083
rect 34793 22043 34851 22049
rect 34808 22012 34836 22043
rect 33060 21984 34468 22012
rect 34532 21984 34836 22012
rect 34900 22012 34928 22120
rect 34992 22120 35256 22148
rect 34992 22089 35020 22120
rect 35250 22108 35256 22120
rect 35308 22148 35314 22160
rect 35529 22151 35587 22157
rect 35529 22148 35541 22151
rect 35308 22120 35541 22148
rect 35308 22108 35314 22120
rect 35529 22117 35541 22120
rect 35575 22117 35587 22151
rect 35529 22111 35587 22117
rect 36630 22108 36636 22160
rect 36688 22108 36694 22160
rect 38010 22108 38016 22160
rect 38068 22108 38074 22160
rect 38746 22148 38752 22160
rect 38580 22120 38752 22148
rect 34977 22083 35035 22089
rect 34977 22049 34989 22083
rect 35023 22080 35035 22083
rect 35023 22052 35057 22080
rect 35023 22049 35035 22052
rect 34977 22043 35035 22049
rect 36078 22040 36084 22092
rect 36136 22040 36142 22092
rect 36648 22080 36676 22108
rect 37001 22083 37059 22089
rect 37001 22080 37013 22083
rect 36648 22052 37013 22080
rect 37001 22049 37013 22052
rect 37047 22080 37059 22083
rect 37277 22083 37335 22089
rect 37277 22080 37289 22083
rect 37047 22052 37289 22080
rect 37047 22049 37059 22052
rect 37001 22043 37059 22049
rect 37277 22049 37289 22052
rect 37323 22049 37335 22083
rect 38580 22080 38608 22120
rect 38746 22108 38752 22120
rect 38804 22108 38810 22160
rect 41506 22108 41512 22160
rect 41564 22108 41570 22160
rect 42610 22108 42616 22160
rect 42668 22148 42674 22160
rect 42668 22120 42840 22148
rect 42668 22108 42674 22120
rect 37277 22043 37335 22049
rect 37568 22052 38608 22080
rect 35802 22012 35808 22024
rect 34900 21984 35808 22012
rect 28068 21947 28126 21953
rect 28068 21913 28080 21947
rect 28114 21944 28126 21947
rect 28258 21944 28264 21956
rect 28114 21916 28264 21944
rect 28114 21913 28126 21916
rect 28068 21907 28126 21913
rect 28258 21904 28264 21916
rect 28316 21904 28322 21956
rect 30834 21904 30840 21956
rect 30892 21944 30898 21956
rect 31294 21944 31300 21956
rect 30892 21916 31300 21944
rect 30892 21904 30898 21916
rect 31294 21904 31300 21916
rect 31352 21944 31358 21956
rect 34532 21953 34560 21984
rect 35802 21972 35808 21984
rect 35860 21972 35866 22024
rect 37568 22021 37596 22052
rect 38654 22040 38660 22092
rect 38712 22080 38718 22092
rect 39301 22083 39359 22089
rect 39301 22080 39313 22083
rect 38712 22052 39313 22080
rect 38712 22040 38718 22052
rect 39301 22049 39313 22052
rect 39347 22049 39359 22083
rect 39301 22043 39359 22049
rect 41322 22040 41328 22092
rect 41380 22080 41386 22092
rect 42812 22089 42840 22120
rect 43622 22108 43628 22160
rect 43680 22148 43686 22160
rect 43717 22151 43775 22157
rect 43717 22148 43729 22151
rect 43680 22120 43729 22148
rect 43680 22108 43686 22120
rect 43717 22117 43729 22120
rect 43763 22117 43775 22151
rect 55585 22151 55643 22157
rect 43717 22111 43775 22117
rect 47872 22120 48314 22148
rect 41417 22083 41475 22089
rect 41417 22080 41429 22083
rect 41380 22052 41429 22080
rect 41380 22040 41386 22052
rect 41417 22049 41429 22052
rect 41463 22080 41475 22083
rect 42797 22083 42855 22089
rect 41463 22052 42564 22080
rect 41463 22049 41475 22052
rect 41417 22043 41475 22049
rect 37553 22015 37611 22021
rect 37553 21981 37565 22015
rect 37599 21981 37611 22015
rect 37553 21975 37611 21981
rect 38565 22015 38623 22021
rect 38565 21981 38577 22015
rect 38611 21981 38623 22015
rect 38565 21975 38623 21981
rect 42153 22015 42211 22021
rect 42153 21981 42165 22015
rect 42199 22012 42211 22015
rect 42199 21984 42288 22012
rect 42199 21981 42211 21984
rect 42153 21975 42211 21981
rect 34517 21947 34575 21953
rect 34517 21944 34529 21947
rect 31352 21916 34529 21944
rect 31352 21904 31358 21916
rect 34517 21913 34529 21916
rect 34563 21913 34575 21947
rect 34517 21907 34575 21913
rect 25317 21879 25375 21885
rect 25317 21876 25329 21879
rect 25096 21848 25329 21876
rect 25096 21836 25102 21848
rect 25317 21845 25329 21848
rect 25363 21845 25375 21879
rect 25317 21839 25375 21845
rect 29181 21879 29239 21885
rect 29181 21845 29193 21879
rect 29227 21876 29239 21879
rect 29270 21876 29276 21888
rect 29227 21848 29276 21876
rect 29227 21845 29239 21848
rect 29181 21839 29239 21845
rect 29270 21836 29276 21848
rect 29328 21836 29334 21888
rect 34054 21836 34060 21888
rect 34112 21836 34118 21888
rect 34882 21836 34888 21888
rect 34940 21876 34946 21888
rect 35069 21879 35127 21885
rect 35069 21876 35081 21879
rect 34940 21848 35081 21876
rect 34940 21836 34946 21848
rect 35069 21845 35081 21848
rect 35115 21845 35127 21879
rect 35069 21839 35127 21845
rect 35437 21879 35495 21885
rect 35437 21845 35449 21879
rect 35483 21876 35495 21879
rect 36722 21876 36728 21888
rect 35483 21848 36728 21876
rect 35483 21845 35495 21848
rect 35437 21839 35495 21845
rect 36722 21836 36728 21848
rect 36780 21836 36786 21888
rect 37461 21879 37519 21885
rect 37461 21845 37473 21879
rect 37507 21876 37519 21879
rect 37642 21876 37648 21888
rect 37507 21848 37648 21876
rect 37507 21845 37519 21848
rect 37461 21839 37519 21845
rect 37642 21836 37648 21848
rect 37700 21836 37706 21888
rect 37921 21879 37979 21885
rect 37921 21845 37933 21879
rect 37967 21876 37979 21879
rect 38580 21876 38608 21975
rect 42260 21885 42288 21984
rect 42536 21944 42564 22052
rect 42797 22049 42809 22083
rect 42843 22080 42855 22083
rect 42843 22052 42877 22080
rect 42843 22049 42855 22052
rect 42797 22043 42855 22049
rect 43070 22040 43076 22092
rect 43128 22040 43134 22092
rect 42613 22015 42671 22021
rect 42613 21981 42625 22015
rect 42659 22012 42671 22015
rect 43640 22012 43668 22108
rect 46382 22040 46388 22092
rect 46440 22080 46446 22092
rect 46842 22080 46848 22092
rect 46440 22052 46848 22080
rect 46440 22040 46446 22052
rect 46842 22040 46848 22052
rect 46900 22080 46906 22092
rect 47872 22089 47900 22120
rect 47029 22083 47087 22089
rect 47029 22080 47041 22083
rect 46900 22052 47041 22080
rect 46900 22040 46906 22052
rect 47029 22049 47041 22052
rect 47075 22049 47087 22083
rect 47857 22083 47915 22089
rect 47857 22080 47869 22083
rect 47029 22043 47087 22049
rect 47504 22052 47869 22080
rect 42659 21984 43668 22012
rect 42659 21981 42671 21984
rect 42613 21975 42671 21981
rect 46934 21972 46940 22024
rect 46992 21972 46998 22024
rect 47504 21944 47532 22052
rect 47857 22049 47869 22052
rect 47903 22049 47915 22083
rect 47857 22043 47915 22049
rect 48038 22040 48044 22092
rect 48096 22040 48102 22092
rect 48286 22080 48314 22120
rect 55585 22117 55597 22151
rect 55631 22148 55643 22151
rect 55950 22148 55956 22160
rect 55631 22120 55956 22148
rect 55631 22117 55643 22120
rect 55585 22111 55643 22117
rect 55950 22108 55956 22120
rect 56008 22108 56014 22160
rect 56502 22148 56508 22160
rect 56060 22120 56508 22148
rect 56060 22092 56088 22120
rect 56502 22108 56508 22120
rect 56560 22108 56566 22160
rect 48286 22052 50292 22080
rect 47578 21972 47584 22024
rect 47636 22012 47642 22024
rect 48133 22015 48191 22021
rect 48133 22012 48145 22015
rect 47636 21984 48145 22012
rect 47636 21972 47642 21984
rect 48133 21981 48145 21984
rect 48179 21981 48191 22015
rect 48133 21975 48191 21981
rect 50154 21972 50160 22024
rect 50212 21972 50218 22024
rect 50264 22012 50292 22052
rect 51350 22040 51356 22092
rect 51408 22080 51414 22092
rect 51721 22083 51779 22089
rect 51721 22080 51733 22083
rect 51408 22052 51733 22080
rect 51408 22040 51414 22052
rect 51721 22049 51733 22052
rect 51767 22049 51779 22083
rect 52638 22080 52644 22092
rect 51721 22043 51779 22049
rect 52196 22052 52644 22080
rect 52196 22012 52224 22052
rect 52638 22040 52644 22052
rect 52696 22040 52702 22092
rect 56042 22080 56048 22092
rect 55232 22052 56048 22080
rect 50264 21984 52224 22012
rect 52365 22015 52423 22021
rect 52365 21981 52377 22015
rect 52411 21981 52423 22015
rect 52365 21975 52423 21981
rect 47673 21947 47731 21953
rect 47673 21944 47685 21947
rect 42536 21916 43208 21944
rect 43180 21888 43208 21916
rect 44652 21916 47685 21944
rect 44652 21888 44680 21916
rect 47673 21913 47685 21916
rect 47719 21913 47731 21947
rect 47673 21907 47731 21913
rect 50424 21947 50482 21953
rect 50424 21913 50436 21947
rect 50470 21944 50482 21947
rect 50982 21944 50988 21956
rect 50470 21916 50988 21944
rect 50470 21913 50482 21916
rect 50424 21907 50482 21913
rect 50982 21904 50988 21916
rect 51040 21904 51046 21956
rect 37967 21848 38608 21876
rect 42245 21879 42303 21885
rect 37967 21845 37979 21848
rect 37921 21839 37979 21845
rect 42245 21845 42257 21879
rect 42291 21845 42303 21879
rect 42245 21839 42303 21845
rect 42705 21879 42763 21885
rect 42705 21845 42717 21879
rect 42751 21876 42763 21879
rect 42886 21876 42892 21888
rect 42751 21848 42892 21876
rect 42751 21845 42763 21848
rect 42705 21839 42763 21845
rect 42886 21836 42892 21848
rect 42944 21836 42950 21888
rect 43162 21836 43168 21888
rect 43220 21836 43226 21888
rect 44634 21836 44640 21888
rect 44692 21836 44698 21888
rect 46474 21836 46480 21888
rect 46532 21836 46538 21888
rect 46658 21836 46664 21888
rect 46716 21876 46722 21888
rect 46845 21879 46903 21885
rect 46845 21876 46857 21879
rect 46716 21848 46857 21876
rect 46716 21836 46722 21848
rect 46845 21845 46857 21848
rect 46891 21876 46903 21879
rect 48314 21876 48320 21888
rect 46891 21848 48320 21876
rect 46891 21845 46903 21848
rect 46845 21839 46903 21845
rect 48314 21836 48320 21848
rect 48372 21836 48378 21888
rect 48501 21879 48559 21885
rect 48501 21845 48513 21879
rect 48547 21876 48559 21879
rect 48958 21876 48964 21888
rect 48547 21848 48964 21876
rect 48547 21845 48559 21848
rect 48501 21839 48559 21845
rect 48958 21836 48964 21848
rect 49016 21836 49022 21888
rect 49973 21879 50031 21885
rect 49973 21845 49985 21879
rect 50019 21876 50031 21879
rect 50062 21876 50068 21888
rect 50019 21848 50068 21876
rect 50019 21845 50031 21848
rect 49973 21839 50031 21845
rect 50062 21836 50068 21848
rect 50120 21876 50126 21888
rect 51074 21876 51080 21888
rect 50120 21848 51080 21876
rect 50120 21836 50126 21848
rect 51074 21836 51080 21848
rect 51132 21836 51138 21888
rect 51537 21879 51595 21885
rect 51537 21845 51549 21879
rect 51583 21876 51595 21879
rect 52380 21876 52408 21975
rect 55232 21888 55260 22052
rect 56042 22040 56048 22052
rect 56100 22040 56106 22092
rect 57149 22083 57207 22089
rect 57149 22080 57161 22083
rect 56428 22052 57161 22080
rect 51583 21848 52408 21876
rect 55033 21879 55091 21885
rect 51583 21845 51595 21848
rect 51537 21839 51595 21845
rect 55033 21845 55045 21879
rect 55079 21876 55091 21879
rect 55214 21876 55220 21888
rect 55079 21848 55220 21876
rect 55079 21845 55091 21848
rect 55033 21839 55091 21845
rect 55214 21836 55220 21848
rect 55272 21836 55278 21888
rect 55858 21836 55864 21888
rect 55916 21876 55922 21888
rect 56428 21885 56456 22052
rect 57149 22049 57161 22052
rect 57195 22049 57207 22083
rect 57149 22043 57207 22049
rect 56962 21972 56968 22024
rect 57020 21972 57026 22024
rect 57057 22015 57115 22021
rect 57057 21981 57069 22015
rect 57103 22012 57115 22015
rect 57790 22012 57796 22024
rect 57103 21984 57796 22012
rect 57103 21981 57115 21984
rect 57057 21975 57115 21981
rect 57790 21972 57796 21984
rect 57848 21972 57854 22024
rect 57974 21972 57980 22024
rect 58032 21972 58038 22024
rect 56413 21879 56471 21885
rect 56413 21876 56425 21879
rect 55916 21848 56425 21876
rect 55916 21836 55922 21848
rect 56413 21845 56425 21848
rect 56459 21845 56471 21879
rect 56413 21839 56471 21845
rect 56597 21879 56655 21885
rect 56597 21845 56609 21879
rect 56643 21876 56655 21879
rect 56870 21876 56876 21888
rect 56643 21848 56876 21876
rect 56643 21845 56655 21848
rect 56597 21839 56655 21845
rect 56870 21836 56876 21848
rect 56928 21836 56934 21888
rect 57422 21836 57428 21888
rect 57480 21836 57486 21888
rect 1104 21786 59040 21808
rect 1104 21734 15394 21786
rect 15446 21734 15458 21786
rect 15510 21734 15522 21786
rect 15574 21734 15586 21786
rect 15638 21734 15650 21786
rect 15702 21734 29838 21786
rect 29890 21734 29902 21786
rect 29954 21734 29966 21786
rect 30018 21734 30030 21786
rect 30082 21734 30094 21786
rect 30146 21734 44282 21786
rect 44334 21734 44346 21786
rect 44398 21734 44410 21786
rect 44462 21734 44474 21786
rect 44526 21734 44538 21786
rect 44590 21734 58726 21786
rect 58778 21734 58790 21786
rect 58842 21734 58854 21786
rect 58906 21734 58918 21786
rect 58970 21734 58982 21786
rect 59034 21734 59040 21786
rect 1104 21712 59040 21734
rect 4709 21675 4767 21681
rect 4709 21641 4721 21675
rect 4755 21672 4767 21675
rect 5166 21672 5172 21684
rect 4755 21644 5172 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 6181 21675 6239 21681
rect 6181 21641 6193 21675
rect 6227 21672 6239 21675
rect 6454 21672 6460 21684
rect 6227 21644 6460 21672
rect 6227 21641 6239 21644
rect 6181 21635 6239 21641
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 7650 21672 7656 21684
rect 6564 21644 7656 21672
rect 5068 21607 5126 21613
rect 5068 21573 5080 21607
rect 5114 21604 5126 21607
rect 5350 21604 5356 21616
rect 5114 21576 5356 21604
rect 5114 21573 5126 21576
rect 5068 21567 5126 21573
rect 5350 21564 5356 21576
rect 5408 21564 5414 21616
rect 6365 21607 6423 21613
rect 6365 21573 6377 21607
rect 6411 21604 6423 21607
rect 6564 21604 6592 21644
rect 7650 21632 7656 21644
rect 7708 21632 7714 21684
rect 8941 21675 8999 21681
rect 8941 21641 8953 21675
rect 8987 21672 8999 21675
rect 9398 21672 9404 21684
rect 8987 21644 9404 21672
rect 8987 21641 8999 21644
rect 8941 21635 8999 21641
rect 8956 21604 8984 21635
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 11054 21632 11060 21684
rect 11112 21632 11118 21684
rect 12069 21675 12127 21681
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 14369 21675 14427 21681
rect 14369 21672 14381 21675
rect 12115 21644 14381 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 14369 21641 14381 21644
rect 14415 21641 14427 21675
rect 14369 21635 14427 21641
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 25682 21672 25688 21684
rect 24912 21644 25688 21672
rect 24912 21632 24918 21644
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 28813 21675 28871 21681
rect 28813 21641 28825 21675
rect 28859 21672 28871 21675
rect 29917 21675 29975 21681
rect 29917 21672 29929 21675
rect 28859 21644 29929 21672
rect 28859 21641 28871 21644
rect 28813 21635 28871 21641
rect 29917 21641 29929 21644
rect 29963 21672 29975 21675
rect 30190 21672 30196 21684
rect 29963 21644 30196 21672
rect 29963 21641 29975 21644
rect 29917 21635 29975 21641
rect 30190 21632 30196 21644
rect 30248 21632 30254 21684
rect 30650 21632 30656 21684
rect 30708 21672 30714 21684
rect 31386 21672 31392 21684
rect 30708 21644 31392 21672
rect 30708 21632 30714 21644
rect 31386 21632 31392 21644
rect 31444 21632 31450 21684
rect 32401 21675 32459 21681
rect 32401 21641 32413 21675
rect 32447 21672 32459 21675
rect 33042 21672 33048 21684
rect 32447 21644 33048 21672
rect 32447 21641 32459 21644
rect 32401 21635 32459 21641
rect 33042 21632 33048 21644
rect 33100 21632 33106 21684
rect 35253 21675 35311 21681
rect 35253 21641 35265 21675
rect 35299 21672 35311 21675
rect 35434 21672 35440 21684
rect 35299 21644 35440 21672
rect 35299 21641 35311 21644
rect 35253 21635 35311 21641
rect 35434 21632 35440 21644
rect 35492 21672 35498 21684
rect 35710 21672 35716 21684
rect 35492 21644 35716 21672
rect 35492 21632 35498 21644
rect 35710 21632 35716 21644
rect 35768 21632 35774 21684
rect 43257 21675 43315 21681
rect 43257 21641 43269 21675
rect 43303 21672 43315 21675
rect 43714 21672 43720 21684
rect 43303 21644 43720 21672
rect 43303 21641 43315 21644
rect 43257 21635 43315 21641
rect 43714 21632 43720 21644
rect 43772 21632 43778 21684
rect 46198 21632 46204 21684
rect 46256 21672 46262 21684
rect 46385 21675 46443 21681
rect 46385 21672 46397 21675
rect 46256 21644 46397 21672
rect 46256 21632 46262 21644
rect 46385 21641 46397 21644
rect 46431 21641 46443 21675
rect 46385 21635 46443 21641
rect 46934 21632 46940 21684
rect 46992 21672 46998 21684
rect 48222 21672 48228 21684
rect 46992 21644 48228 21672
rect 46992 21632 46998 21644
rect 48222 21632 48228 21644
rect 48280 21632 48286 21684
rect 50982 21632 50988 21684
rect 51040 21632 51046 21684
rect 51166 21632 51172 21684
rect 51224 21672 51230 21684
rect 54757 21675 54815 21681
rect 54757 21672 54769 21675
rect 51224 21644 54769 21672
rect 51224 21632 51230 21644
rect 54757 21641 54769 21644
rect 54803 21672 54815 21675
rect 55398 21672 55404 21684
rect 54803 21644 55404 21672
rect 54803 21641 54815 21644
rect 54757 21635 54815 21641
rect 55398 21632 55404 21644
rect 55456 21672 55462 21684
rect 55950 21672 55956 21684
rect 55456 21644 55956 21672
rect 55456 21632 55462 21644
rect 55950 21632 55956 21644
rect 56008 21632 56014 21684
rect 56686 21632 56692 21684
rect 56744 21632 56750 21684
rect 57149 21675 57207 21681
rect 57149 21641 57161 21675
rect 57195 21672 57207 21675
rect 57974 21672 57980 21684
rect 57195 21644 57980 21672
rect 57195 21641 57207 21644
rect 57149 21635 57207 21641
rect 57974 21632 57980 21644
rect 58032 21632 58038 21684
rect 6411 21576 6592 21604
rect 8220 21576 8984 21604
rect 6411 21573 6423 21576
rect 6365 21567 6423 21573
rect 7190 21545 7196 21548
rect 7168 21539 7196 21545
rect 7168 21505 7180 21539
rect 7168 21499 7196 21505
rect 7190 21496 7196 21499
rect 7248 21496 7254 21548
rect 7282 21496 7288 21548
rect 7340 21496 7346 21548
rect 8220 21545 8248 21576
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 14461 21607 14519 21613
rect 14461 21604 14473 21607
rect 13872 21576 14473 21604
rect 13872 21564 13878 21576
rect 14461 21573 14473 21576
rect 14507 21573 14519 21607
rect 14461 21567 14519 21573
rect 28905 21607 28963 21613
rect 28905 21573 28917 21607
rect 28951 21604 28963 21607
rect 28994 21604 29000 21616
rect 28951 21576 29000 21604
rect 28951 21573 28963 21576
rect 28905 21567 28963 21573
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 50525 21607 50583 21613
rect 50525 21573 50537 21607
rect 50571 21604 50583 21607
rect 51350 21604 51356 21616
rect 50571 21576 51356 21604
rect 50571 21573 50583 21576
rect 50525 21567 50583 21573
rect 51350 21564 51356 21576
rect 51408 21564 51414 21616
rect 52822 21564 52828 21616
rect 52880 21604 52886 21616
rect 54389 21607 54447 21613
rect 54389 21604 54401 21607
rect 52880 21576 54401 21604
rect 52880 21564 52886 21576
rect 54389 21573 54401 21576
rect 54435 21604 54447 21607
rect 55214 21604 55220 21616
rect 54435 21576 55220 21604
rect 54435 21573 54447 21576
rect 54389 21567 54447 21573
rect 55214 21564 55220 21576
rect 55272 21564 55278 21616
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 8294 21496 8300 21548
rect 8352 21496 8358 21548
rect 9122 21496 9128 21548
rect 9180 21496 9186 21548
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11011 21508 11928 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 4801 21471 4859 21477
rect 4801 21437 4813 21471
rect 4847 21437 4859 21471
rect 4801 21431 4859 21437
rect 4816 21332 4844 21431
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 7064 21440 7696 21468
rect 7064 21428 7070 21440
rect 7561 21403 7619 21409
rect 7561 21369 7573 21403
rect 7607 21369 7619 21403
rect 7561 21363 7619 21369
rect 5902 21332 5908 21344
rect 4816 21304 5908 21332
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 7282 21292 7288 21344
rect 7340 21332 7346 21344
rect 7576 21332 7604 21363
rect 7340 21304 7604 21332
rect 7668 21332 7696 21440
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 8021 21471 8079 21477
rect 8021 21468 8033 21471
rect 7984 21440 8033 21468
rect 7984 21428 7990 21440
rect 8021 21437 8033 21440
rect 8067 21437 8079 21471
rect 8021 21431 8079 21437
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 9953 21431 10011 21437
rect 10704 21440 11161 21468
rect 9968 21400 9996 21431
rect 10597 21403 10655 21409
rect 10597 21400 10609 21403
rect 9968 21372 10609 21400
rect 10597 21369 10609 21372
rect 10643 21369 10655 21403
rect 10597 21363 10655 21369
rect 10704 21344 10732 21440
rect 11149 21437 11161 21440
rect 11195 21437 11207 21471
rect 11900 21468 11928 21508
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 12986 21496 12992 21548
rect 13044 21496 13050 21548
rect 13906 21496 13912 21548
rect 13964 21496 13970 21548
rect 29270 21496 29276 21548
rect 29328 21496 29334 21548
rect 30374 21496 30380 21548
rect 30432 21496 30438 21548
rect 42242 21496 42248 21548
rect 42300 21536 42306 21548
rect 42613 21539 42671 21545
rect 42613 21536 42625 21539
rect 42300 21508 42625 21536
rect 42300 21496 42306 21508
rect 42613 21505 42625 21508
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 46474 21496 46480 21548
rect 46532 21536 46538 21548
rect 46937 21539 46995 21545
rect 46937 21536 46949 21539
rect 46532 21508 46949 21536
rect 46532 21496 46538 21508
rect 46937 21505 46949 21508
rect 46983 21505 46995 21539
rect 46937 21499 46995 21505
rect 47302 21496 47308 21548
rect 47360 21536 47366 21548
rect 47581 21539 47639 21545
rect 47581 21536 47593 21539
rect 47360 21508 47593 21536
rect 47360 21496 47366 21508
rect 47581 21505 47593 21508
rect 47627 21505 47639 21539
rect 47581 21499 47639 21505
rect 48958 21496 48964 21548
rect 49016 21496 49022 21548
rect 52365 21539 52423 21545
rect 49252 21508 52316 21536
rect 12342 21468 12348 21480
rect 11900 21440 12348 21468
rect 11149 21431 11207 21437
rect 12342 21428 12348 21440
rect 12400 21468 12406 21480
rect 12851 21471 12909 21477
rect 12851 21468 12863 21471
rect 12400 21440 12863 21468
rect 12400 21428 12406 21440
rect 12851 21437 12863 21440
rect 12897 21437 12909 21471
rect 12851 21431 12909 21437
rect 13725 21471 13783 21477
rect 13725 21437 13737 21471
rect 13771 21468 13783 21471
rect 14458 21468 14464 21480
rect 13771 21440 14464 21468
rect 13771 21437 13783 21440
rect 13725 21431 13783 21437
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21437 14611 21471
rect 14553 21431 14611 21437
rect 13170 21360 13176 21412
rect 13228 21400 13234 21412
rect 13265 21403 13323 21409
rect 13265 21400 13277 21403
rect 13228 21372 13277 21400
rect 13228 21360 13234 21372
rect 13265 21369 13277 21372
rect 13311 21369 13323 21403
rect 14568 21400 14596 21431
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 19058 21428 19064 21480
rect 19116 21428 19122 21480
rect 28997 21471 29055 21477
rect 28997 21468 29009 21471
rect 28368 21440 29009 21468
rect 17034 21400 17040 21412
rect 13265 21363 13323 21369
rect 13924 21372 17040 21400
rect 13924 21344 13952 21372
rect 17034 21360 17040 21372
rect 17092 21360 17098 21412
rect 28368 21344 28396 21440
rect 28997 21437 29009 21440
rect 29043 21437 29055 21471
rect 28997 21431 29055 21437
rect 36722 21428 36728 21480
rect 36780 21468 36786 21480
rect 37093 21471 37151 21477
rect 37093 21468 37105 21471
rect 36780 21440 37105 21468
rect 36780 21428 36786 21440
rect 37093 21437 37105 21440
rect 37139 21468 37151 21471
rect 42518 21468 42524 21480
rect 37139 21440 42524 21468
rect 37139 21437 37151 21440
rect 37093 21431 37151 21437
rect 42518 21428 42524 21440
rect 42576 21428 42582 21480
rect 48590 21428 48596 21480
rect 48648 21468 48654 21480
rect 49145 21471 49203 21477
rect 49145 21468 49157 21471
rect 48648 21440 49157 21468
rect 48648 21428 48654 21440
rect 49145 21437 49157 21440
rect 49191 21437 49203 21471
rect 49145 21431 49203 21437
rect 29638 21360 29644 21412
rect 29696 21400 29702 21412
rect 49252 21400 49280 21508
rect 50246 21428 50252 21480
rect 50304 21428 50310 21480
rect 50433 21471 50491 21477
rect 50433 21437 50445 21471
rect 50479 21468 50491 21471
rect 50798 21468 50804 21480
rect 50479 21440 50804 21468
rect 50479 21437 50491 21440
rect 50433 21431 50491 21437
rect 50798 21428 50804 21440
rect 50856 21468 50862 21480
rect 51258 21468 51264 21480
rect 50856 21440 51264 21468
rect 50856 21428 50862 21440
rect 51258 21428 51264 21440
rect 51316 21428 51322 21480
rect 51537 21471 51595 21477
rect 51537 21437 51549 21471
rect 51583 21437 51595 21471
rect 52288 21468 52316 21508
rect 52365 21505 52377 21539
rect 52411 21536 52423 21539
rect 52730 21536 52736 21548
rect 52411 21508 52736 21536
rect 52411 21505 52423 21508
rect 52365 21499 52423 21505
rect 52730 21496 52736 21508
rect 52788 21496 52794 21548
rect 55766 21496 55772 21548
rect 55824 21536 55830 21548
rect 56781 21539 56839 21545
rect 56781 21536 56793 21539
rect 55824 21508 56793 21536
rect 55824 21496 55830 21508
rect 56781 21505 56793 21508
rect 56827 21505 56839 21539
rect 56781 21499 56839 21505
rect 56229 21471 56287 21477
rect 56229 21468 56241 21471
rect 52288 21440 56241 21468
rect 51537 21431 51595 21437
rect 56229 21437 56241 21440
rect 56275 21468 56287 21471
rect 56505 21471 56563 21477
rect 56505 21468 56517 21471
rect 56275 21440 56517 21468
rect 56275 21437 56287 21440
rect 56229 21431 56287 21437
rect 56505 21437 56517 21440
rect 56551 21437 56563 21471
rect 56505 21431 56563 21437
rect 29696 21372 49280 21400
rect 50893 21403 50951 21409
rect 29696 21360 29702 21372
rect 50893 21369 50905 21403
rect 50939 21400 50951 21403
rect 51552 21400 51580 21431
rect 57606 21428 57612 21480
rect 57664 21468 57670 21480
rect 58437 21471 58495 21477
rect 58437 21468 58449 21471
rect 57664 21440 58449 21468
rect 57664 21428 57670 21440
rect 58437 21437 58449 21440
rect 58483 21437 58495 21471
rect 58437 21431 58495 21437
rect 50939 21372 51580 21400
rect 50939 21369 50951 21372
rect 50893 21363 50951 21369
rect 8018 21332 8024 21344
rect 7668 21304 8024 21332
rect 7340 21292 7346 21304
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 8754 21332 8760 21344
rect 8536 21304 8760 21332
rect 8536 21292 8542 21304
rect 8754 21292 8760 21304
rect 8812 21292 8818 21344
rect 9766 21292 9772 21344
rect 9824 21292 9830 21344
rect 10502 21292 10508 21344
rect 10560 21292 10566 21344
rect 10686 21292 10692 21344
rect 10744 21292 10750 21344
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12710 21332 12716 21344
rect 12032 21304 12716 21332
rect 12032 21292 12038 21304
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15344 21304 15577 21332
rect 15344 21292 15350 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 15565 21295 15623 21301
rect 19610 21292 19616 21344
rect 19668 21292 19674 21344
rect 25317 21335 25375 21341
rect 25317 21301 25329 21335
rect 25363 21332 25375 21335
rect 25958 21332 25964 21344
rect 25363 21304 25964 21332
rect 25363 21301 25375 21304
rect 25317 21295 25375 21301
rect 25958 21292 25964 21304
rect 26016 21332 26022 21344
rect 28350 21332 28356 21344
rect 26016 21304 28356 21332
rect 26016 21292 26022 21304
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 28442 21292 28448 21344
rect 28500 21292 28506 21344
rect 31018 21292 31024 21344
rect 31076 21292 31082 21344
rect 35618 21292 35624 21344
rect 35676 21292 35682 21344
rect 37553 21335 37611 21341
rect 37553 21301 37565 21335
rect 37599 21332 37611 21335
rect 37826 21332 37832 21344
rect 37599 21304 37832 21332
rect 37599 21301 37611 21304
rect 37553 21295 37611 21301
rect 37826 21292 37832 21304
rect 37884 21292 37890 21344
rect 42150 21292 42156 21344
rect 42208 21332 42214 21344
rect 42610 21332 42616 21344
rect 42208 21304 42616 21332
rect 42208 21292 42214 21304
rect 42610 21292 42616 21304
rect 42668 21292 42674 21344
rect 48406 21292 48412 21344
rect 48464 21292 48470 21344
rect 49050 21292 49056 21344
rect 49108 21332 49114 21344
rect 49789 21335 49847 21341
rect 49789 21332 49801 21335
rect 49108 21304 49801 21332
rect 49108 21292 49114 21304
rect 49789 21301 49801 21304
rect 49835 21301 49847 21335
rect 49789 21295 49847 21301
rect 51350 21292 51356 21344
rect 51408 21332 51414 21344
rect 51721 21335 51779 21341
rect 51721 21332 51733 21335
rect 51408 21304 51733 21332
rect 51408 21292 51414 21304
rect 51721 21301 51733 21304
rect 51767 21301 51779 21335
rect 51721 21295 51779 21301
rect 56778 21292 56784 21344
rect 56836 21332 56842 21344
rect 57425 21335 57483 21341
rect 57425 21332 57437 21335
rect 56836 21304 57437 21332
rect 56836 21292 56842 21304
rect 57425 21301 57437 21304
rect 57471 21301 57483 21335
rect 57425 21295 57483 21301
rect 57882 21292 57888 21344
rect 57940 21292 57946 21344
rect 1104 21242 58880 21264
rect 1104 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 22616 21242
rect 22668 21190 22680 21242
rect 22732 21190 22744 21242
rect 22796 21190 22808 21242
rect 22860 21190 22872 21242
rect 22924 21190 37060 21242
rect 37112 21190 37124 21242
rect 37176 21190 37188 21242
rect 37240 21190 37252 21242
rect 37304 21190 37316 21242
rect 37368 21190 51504 21242
rect 51556 21190 51568 21242
rect 51620 21190 51632 21242
rect 51684 21190 51696 21242
rect 51748 21190 51760 21242
rect 51812 21190 58880 21242
rect 1104 21168 58880 21190
rect 4154 21088 4160 21140
rect 4212 21128 4218 21140
rect 4525 21131 4583 21137
rect 4525 21128 4537 21131
rect 4212 21100 4537 21128
rect 4212 21088 4218 21100
rect 4525 21097 4537 21100
rect 4571 21097 4583 21131
rect 4525 21091 4583 21097
rect 7282 21088 7288 21140
rect 7340 21088 7346 21140
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 10229 21131 10287 21137
rect 10229 21128 10241 21131
rect 7616 21100 10241 21128
rect 7616 21088 7622 21100
rect 10229 21097 10241 21100
rect 10275 21128 10287 21131
rect 10686 21128 10692 21140
rect 10275 21100 10692 21128
rect 10275 21097 10287 21100
rect 10229 21091 10287 21097
rect 10686 21088 10692 21100
rect 10744 21128 10750 21140
rect 10744 21100 12296 21128
rect 10744 21088 10750 21100
rect 7300 21060 7328 21088
rect 9125 21063 9183 21069
rect 9125 21060 9137 21063
rect 7300 21032 9137 21060
rect 9125 21029 9137 21032
rect 9171 21029 9183 21063
rect 9125 21023 9183 21029
rect 11793 21063 11851 21069
rect 11793 21029 11805 21063
rect 11839 21060 11851 21063
rect 11839 21032 11928 21060
rect 11839 21029 11851 21032
rect 11793 21023 11851 21029
rect 9674 20992 9680 21004
rect 7392 20964 9680 20992
rect 5902 20884 5908 20936
rect 5960 20924 5966 20936
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 5960 20896 6377 20924
rect 5960 20884 5966 20896
rect 6365 20893 6377 20896
rect 6411 20924 6423 20927
rect 7392 20924 7420 20964
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 11900 21001 11928 21032
rect 11974 21020 11980 21072
rect 12032 21020 12038 21072
rect 12268 21060 12296 21100
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 12529 21131 12587 21137
rect 12529 21128 12541 21131
rect 12400 21100 12541 21128
rect 12400 21088 12406 21100
rect 12529 21097 12541 21100
rect 12575 21097 12587 21131
rect 12529 21091 12587 21097
rect 15749 21131 15807 21137
rect 15749 21097 15761 21131
rect 15795 21128 15807 21131
rect 16114 21128 16120 21140
rect 15795 21100 16120 21128
rect 15795 21097 15807 21100
rect 15749 21091 15807 21097
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 17218 21088 17224 21140
rect 17276 21088 17282 21140
rect 28258 21088 28264 21140
rect 28316 21088 28322 21140
rect 28442 21088 28448 21140
rect 28500 21088 28506 21140
rect 33318 21088 33324 21140
rect 33376 21128 33382 21140
rect 34054 21128 34060 21140
rect 33376 21100 34060 21128
rect 33376 21088 33382 21100
rect 34054 21088 34060 21100
rect 34112 21128 34118 21140
rect 34885 21131 34943 21137
rect 34885 21128 34897 21131
rect 34112 21100 34897 21128
rect 34112 21088 34118 21100
rect 34885 21097 34897 21100
rect 34931 21128 34943 21131
rect 42153 21131 42211 21137
rect 34931 21100 38332 21128
rect 34931 21097 34943 21100
rect 34885 21091 34943 21097
rect 17236 21060 17264 21088
rect 12268 21032 15700 21060
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 10376 20964 10425 20992
rect 10376 20952 10382 20964
rect 10413 20961 10425 20964
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20961 11943 20995
rect 11885 20955 11943 20961
rect 7837 20927 7895 20933
rect 7837 20924 7849 20927
rect 6411 20896 7420 20924
rect 7760 20896 7849 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 5534 20816 5540 20868
rect 5592 20856 5598 20868
rect 5638 20859 5696 20865
rect 5638 20856 5650 20859
rect 5592 20828 5650 20856
rect 5592 20816 5598 20828
rect 5638 20825 5650 20828
rect 5684 20825 5696 20859
rect 5638 20819 5696 20825
rect 6632 20859 6690 20865
rect 6632 20825 6644 20859
rect 6678 20856 6690 20859
rect 7190 20856 7196 20868
rect 6678 20828 7196 20856
rect 6678 20825 6690 20828
rect 6632 20819 6690 20825
rect 7190 20816 7196 20828
rect 7248 20816 7254 20868
rect 5994 20748 6000 20800
rect 6052 20788 6058 20800
rect 7466 20788 7472 20800
rect 6052 20760 7472 20788
rect 6052 20748 6058 20760
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 7760 20797 7788 20896
rect 7837 20893 7849 20896
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 10669 20927 10727 20933
rect 10669 20924 10681 20927
rect 10560 20896 10681 20924
rect 10560 20884 10566 20896
rect 10669 20893 10681 20896
rect 10715 20893 10727 20927
rect 10669 20887 10727 20893
rect 8018 20816 8024 20868
rect 8076 20856 8082 20868
rect 9585 20859 9643 20865
rect 9585 20856 9597 20859
rect 8076 20828 9597 20856
rect 8076 20816 8082 20828
rect 9585 20825 9597 20828
rect 9631 20856 9643 20859
rect 11992 20856 12020 21020
rect 13446 20884 13452 20936
rect 13504 20884 13510 20936
rect 15672 20865 15700 21032
rect 16132 21032 17264 21060
rect 16132 20933 16160 21032
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20992 16451 20995
rect 18598 20992 18604 21004
rect 16439 20964 18604 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 9631 20828 12020 20856
rect 15657 20859 15715 20865
rect 9631 20825 9643 20828
rect 9585 20819 9643 20825
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16408 20856 16436 20955
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 28460 20992 28488 21088
rect 38304 21072 38332 21100
rect 42153 21097 42165 21131
rect 42199 21128 42211 21131
rect 46382 21128 46388 21140
rect 42199 21100 46388 21128
rect 42199 21097 42211 21100
rect 42153 21091 42211 21097
rect 38286 21020 38292 21072
rect 38344 21020 38350 21072
rect 28813 20995 28871 21001
rect 28813 20992 28825 20995
rect 28460 20964 28825 20992
rect 28813 20961 28825 20964
rect 28859 20961 28871 20995
rect 28813 20955 28871 20961
rect 36722 20952 36728 21004
rect 36780 20952 36786 21004
rect 37826 20952 37832 21004
rect 37884 20992 37890 21004
rect 42444 21001 42472 21100
rect 46382 21088 46388 21100
rect 46440 21088 46446 21140
rect 46750 21088 46756 21140
rect 46808 21128 46814 21140
rect 50246 21128 50252 21140
rect 46808 21100 50252 21128
rect 46808 21088 46814 21100
rect 50246 21088 50252 21100
rect 50304 21128 50310 21140
rect 50341 21131 50399 21137
rect 50341 21128 50353 21131
rect 50304 21100 50353 21128
rect 50304 21088 50310 21100
rect 50341 21097 50353 21100
rect 50387 21128 50399 21131
rect 51629 21131 51687 21137
rect 50387 21100 51074 21128
rect 50387 21097 50399 21100
rect 50341 21091 50399 21097
rect 42981 21063 43039 21069
rect 42981 21029 42993 21063
rect 43027 21029 43039 21063
rect 42981 21023 43039 21029
rect 42429 20995 42487 21001
rect 42429 20992 42441 20995
rect 37884 20964 42441 20992
rect 37884 20952 37890 20964
rect 42429 20961 42441 20964
rect 42475 20961 42487 20995
rect 42996 20992 43024 21023
rect 44818 21020 44824 21072
rect 44876 21060 44882 21072
rect 45189 21063 45247 21069
rect 45189 21060 45201 21063
rect 44876 21032 45201 21060
rect 44876 21020 44882 21032
rect 45189 21029 45201 21032
rect 45235 21029 45247 21063
rect 45189 21023 45247 21029
rect 43625 20995 43683 21001
rect 43625 20992 43637 20995
rect 42996 20964 43637 20992
rect 42429 20955 42487 20961
rect 43625 20961 43637 20964
rect 43671 20961 43683 20995
rect 43625 20955 43683 20961
rect 16574 20884 16580 20936
rect 16632 20884 16638 20936
rect 19334 20884 19340 20936
rect 19392 20884 19398 20936
rect 22925 20927 22983 20933
rect 22925 20893 22937 20927
rect 22971 20924 22983 20927
rect 23014 20924 23020 20936
rect 22971 20896 23020 20924
rect 22971 20893 22983 20896
rect 22925 20887 22983 20893
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 25222 20884 25228 20936
rect 25280 20884 25286 20936
rect 25314 20884 25320 20936
rect 25372 20884 25378 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 25832 20896 26065 20924
rect 25832 20884 25838 20896
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 27522 20884 27528 20936
rect 27580 20884 27586 20936
rect 29730 20884 29736 20936
rect 29788 20884 29794 20936
rect 34146 20884 34152 20936
rect 34204 20884 34210 20936
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20924 35219 20927
rect 36740 20924 36768 20952
rect 35207 20896 36768 20924
rect 35207 20893 35219 20896
rect 35161 20887 35219 20893
rect 37550 20884 37556 20936
rect 37608 20884 37614 20936
rect 37734 20884 37740 20936
rect 37792 20884 37798 20936
rect 38930 20884 38936 20936
rect 38988 20884 38994 20936
rect 40494 20884 40500 20936
rect 40552 20924 40558 20936
rect 40773 20927 40831 20933
rect 40773 20924 40785 20927
rect 40552 20896 40785 20924
rect 40552 20884 40558 20896
rect 40773 20893 40785 20896
rect 40819 20893 40831 20927
rect 40773 20887 40831 20893
rect 42334 20884 42340 20936
rect 42392 20924 42398 20936
rect 43162 20924 43168 20936
rect 42392 20896 43168 20924
rect 42392 20884 42398 20896
rect 43162 20884 43168 20896
rect 43220 20884 43226 20936
rect 44174 20884 44180 20936
rect 44232 20924 44238 20936
rect 44361 20927 44419 20933
rect 44361 20924 44373 20927
rect 44232 20896 44373 20924
rect 44232 20884 44238 20896
rect 44361 20893 44373 20896
rect 44407 20893 44419 20927
rect 44361 20887 44419 20893
rect 15703 20828 16436 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 36722 20816 36728 20868
rect 36780 20856 36786 20868
rect 37001 20859 37059 20865
rect 37001 20856 37013 20859
rect 36780 20828 37013 20856
rect 36780 20816 36786 20828
rect 37001 20825 37013 20828
rect 37047 20825 37059 20859
rect 37001 20819 37059 20825
rect 40129 20859 40187 20865
rect 40129 20825 40141 20859
rect 40175 20856 40187 20859
rect 42521 20859 42579 20865
rect 40175 20828 40448 20856
rect 40175 20825 40187 20828
rect 40129 20819 40187 20825
rect 40420 20800 40448 20828
rect 42521 20825 42533 20859
rect 42567 20856 42579 20859
rect 43809 20859 43867 20865
rect 43809 20856 43821 20859
rect 42567 20828 43821 20856
rect 42567 20825 42579 20828
rect 42521 20819 42579 20825
rect 43809 20825 43821 20828
rect 43855 20856 43867 20859
rect 43898 20856 43904 20868
rect 43855 20828 43904 20856
rect 43855 20825 43867 20828
rect 43809 20819 43867 20825
rect 43898 20816 43904 20828
rect 43956 20816 43962 20868
rect 51046 20856 51074 21100
rect 51629 21097 51641 21131
rect 51675 21128 51687 21131
rect 52086 21128 52092 21140
rect 51675 21100 52092 21128
rect 51675 21097 51687 21100
rect 51629 21091 51687 21097
rect 52086 21088 52092 21100
rect 52144 21128 52150 21140
rect 52362 21128 52368 21140
rect 52144 21100 52368 21128
rect 52144 21088 52150 21100
rect 52362 21088 52368 21100
rect 52420 21088 52426 21140
rect 57606 21088 57612 21140
rect 57664 21088 57670 21140
rect 57882 21088 57888 21140
rect 57940 21088 57946 21140
rect 52178 20884 52184 20936
rect 52236 20884 52242 20936
rect 53558 20884 53564 20936
rect 53616 20924 53622 20936
rect 53929 20927 53987 20933
rect 53929 20924 53941 20927
rect 53616 20896 53941 20924
rect 53616 20884 53622 20896
rect 53929 20893 53941 20896
rect 53975 20893 53987 20927
rect 53929 20887 53987 20893
rect 54294 20884 54300 20936
rect 54352 20884 54358 20936
rect 55674 20884 55680 20936
rect 55732 20924 55738 20936
rect 56137 20927 56195 20933
rect 56137 20924 56149 20927
rect 55732 20896 56149 20924
rect 55732 20884 55738 20896
rect 56137 20893 56149 20896
rect 56183 20893 56195 20927
rect 56137 20887 56195 20893
rect 56404 20927 56462 20933
rect 56404 20893 56416 20927
rect 56450 20924 56462 20927
rect 57900 20924 57928 21088
rect 58161 20995 58219 21001
rect 58161 20961 58173 20995
rect 58207 20961 58219 20995
rect 58161 20955 58219 20961
rect 56450 20896 57928 20924
rect 56450 20893 56462 20896
rect 56404 20887 56462 20893
rect 53834 20856 53840 20868
rect 51046 20828 53840 20856
rect 53834 20816 53840 20828
rect 53892 20816 53898 20868
rect 56778 20816 56784 20868
rect 56836 20856 56842 20868
rect 58176 20856 58204 20955
rect 56836 20828 58204 20856
rect 56836 20816 56842 20828
rect 7745 20791 7803 20797
rect 7745 20757 7757 20791
rect 7791 20757 7803 20791
rect 7745 20751 7803 20757
rect 7926 20748 7932 20800
rect 7984 20788 7990 20800
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 7984 20760 8493 20788
rect 7984 20748 7990 20760
rect 8481 20757 8493 20760
rect 8527 20757 8539 20791
rect 8481 20751 8539 20757
rect 12802 20748 12808 20800
rect 12860 20748 12866 20800
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 15838 20748 15844 20800
rect 15896 20788 15902 20800
rect 16209 20791 16267 20797
rect 16209 20788 16221 20791
rect 15896 20760 16221 20788
rect 15896 20748 15902 20760
rect 16209 20757 16221 20760
rect 16255 20757 16267 20791
rect 16209 20751 16267 20757
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 19576 20760 19993 20788
rect 19576 20748 19582 20760
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 19981 20751 20039 20757
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22002 20788 22008 20800
rect 21867 20760 22008 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 22281 20791 22339 20797
rect 22281 20757 22293 20791
rect 22327 20788 22339 20791
rect 22370 20788 22376 20800
rect 22327 20760 22376 20788
rect 22327 20757 22339 20760
rect 22281 20751 22339 20757
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 22462 20748 22468 20800
rect 22520 20788 22526 20800
rect 23017 20791 23075 20797
rect 23017 20788 23029 20791
rect 22520 20760 23029 20788
rect 22520 20748 22526 20760
rect 23017 20757 23029 20760
rect 23063 20757 23075 20791
rect 23017 20751 23075 20757
rect 24578 20748 24584 20800
rect 24636 20748 24642 20800
rect 25961 20791 26019 20797
rect 25961 20757 25973 20791
rect 26007 20788 26019 20791
rect 26050 20788 26056 20800
rect 26007 20760 26056 20788
rect 26007 20757 26019 20760
rect 25961 20751 26019 20757
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 26510 20748 26516 20800
rect 26568 20788 26574 20800
rect 26697 20791 26755 20797
rect 26697 20788 26709 20791
rect 26568 20760 26709 20788
rect 26568 20748 26574 20760
rect 26697 20757 26709 20760
rect 26743 20757 26755 20791
rect 26697 20751 26755 20757
rect 26878 20748 26884 20800
rect 26936 20788 26942 20800
rect 26973 20791 27031 20797
rect 26973 20788 26985 20791
rect 26936 20760 26985 20788
rect 26936 20748 26942 20760
rect 26973 20757 26985 20760
rect 27019 20757 27031 20791
rect 26973 20751 27031 20757
rect 30374 20748 30380 20800
rect 30432 20748 30438 20800
rect 32033 20791 32091 20797
rect 32033 20757 32045 20791
rect 32079 20788 32091 20791
rect 32674 20788 32680 20800
rect 32079 20760 32680 20788
rect 32079 20757 32091 20760
rect 32033 20751 32091 20757
rect 32674 20748 32680 20760
rect 32732 20748 32738 20800
rect 33594 20748 33600 20800
rect 33652 20748 33658 20800
rect 36633 20791 36691 20797
rect 36633 20757 36645 20791
rect 36679 20788 36691 20791
rect 36906 20788 36912 20800
rect 36679 20760 36912 20788
rect 36679 20757 36691 20760
rect 36633 20751 36691 20757
rect 36906 20748 36912 20760
rect 36964 20748 36970 20800
rect 38378 20748 38384 20800
rect 38436 20748 38442 20800
rect 38746 20748 38752 20800
rect 38804 20748 38810 20800
rect 39574 20748 39580 20800
rect 39632 20748 39638 20800
rect 40218 20748 40224 20800
rect 40276 20748 40282 20800
rect 40402 20748 40408 20800
rect 40460 20748 40466 20800
rect 42613 20791 42671 20797
rect 42613 20757 42625 20791
rect 42659 20788 42671 20791
rect 42886 20788 42892 20800
rect 42659 20760 42892 20788
rect 42659 20757 42671 20760
rect 42613 20751 42671 20757
rect 42886 20748 42892 20760
rect 42944 20748 42950 20800
rect 43070 20748 43076 20800
rect 43128 20748 43134 20800
rect 44634 20748 44640 20800
rect 44692 20788 44698 20800
rect 44729 20791 44787 20797
rect 44729 20788 44741 20791
rect 44692 20760 44741 20788
rect 44692 20748 44698 20760
rect 44729 20757 44741 20760
rect 44775 20757 44787 20791
rect 44729 20751 44787 20757
rect 45554 20748 45560 20800
rect 45612 20748 45618 20800
rect 53190 20748 53196 20800
rect 53248 20788 53254 20800
rect 53377 20791 53435 20797
rect 53377 20788 53389 20791
rect 53248 20760 53389 20788
rect 53248 20748 53254 20760
rect 53377 20757 53389 20760
rect 53423 20757 53435 20791
rect 53377 20751 53435 20757
rect 54018 20748 54024 20800
rect 54076 20788 54082 20800
rect 54846 20788 54852 20800
rect 54076 20760 54852 20788
rect 54076 20748 54082 20760
rect 54846 20748 54852 20760
rect 54904 20748 54910 20800
rect 56045 20791 56103 20797
rect 56045 20757 56057 20791
rect 56091 20788 56103 20791
rect 56318 20788 56324 20800
rect 56091 20760 56324 20788
rect 56091 20757 56103 20760
rect 56045 20751 56103 20757
rect 56318 20748 56324 20760
rect 56376 20748 56382 20800
rect 57514 20748 57520 20800
rect 57572 20748 57578 20800
rect 57974 20748 57980 20800
rect 58032 20748 58038 20800
rect 58066 20748 58072 20800
rect 58124 20748 58130 20800
rect 1104 20698 59040 20720
rect 1104 20646 15394 20698
rect 15446 20646 15458 20698
rect 15510 20646 15522 20698
rect 15574 20646 15586 20698
rect 15638 20646 15650 20698
rect 15702 20646 29838 20698
rect 29890 20646 29902 20698
rect 29954 20646 29966 20698
rect 30018 20646 30030 20698
rect 30082 20646 30094 20698
rect 30146 20646 44282 20698
rect 44334 20646 44346 20698
rect 44398 20646 44410 20698
rect 44462 20646 44474 20698
rect 44526 20646 44538 20698
rect 44590 20646 58726 20698
rect 58778 20646 58790 20698
rect 58842 20646 58854 20698
rect 58906 20646 58918 20698
rect 58970 20646 58982 20698
rect 59034 20646 59040 20698
rect 1104 20624 59040 20646
rect 5445 20587 5503 20593
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 5534 20584 5540 20596
rect 5491 20556 5540 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 7190 20544 7196 20596
rect 7248 20584 7254 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7248 20556 7757 20584
rect 7248 20544 7254 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 7745 20547 7803 20553
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13504 20556 13645 20584
rect 13504 20544 13510 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 13998 20544 14004 20596
rect 14056 20544 14062 20596
rect 15286 20584 15292 20596
rect 15273 20544 15292 20584
rect 15344 20544 15350 20596
rect 16485 20587 16543 20593
rect 16485 20553 16497 20587
rect 16531 20584 16543 20587
rect 16574 20584 16580 20596
rect 16531 20556 16580 20584
rect 16531 20553 16543 20556
rect 16485 20547 16543 20553
rect 16574 20544 16580 20556
rect 16632 20544 16638 20596
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 17310 20584 17316 20596
rect 16724 20556 17316 20584
rect 16724 20544 16730 20556
rect 17310 20544 17316 20556
rect 17368 20584 17374 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17368 20556 17601 20584
rect 17368 20544 17374 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 18509 20587 18567 20593
rect 18509 20553 18521 20587
rect 18555 20584 18567 20587
rect 19334 20584 19340 20596
rect 18555 20556 19340 20584
rect 18555 20553 18567 20556
rect 18509 20547 18567 20553
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 22281 20587 22339 20593
rect 22281 20553 22293 20587
rect 22327 20584 22339 20587
rect 22462 20584 22468 20596
rect 22327 20556 22468 20584
rect 22327 20553 22339 20556
rect 22281 20547 22339 20553
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 24854 20584 24860 20596
rect 24136 20556 24860 20584
rect 7285 20519 7343 20525
rect 7285 20485 7297 20519
rect 7331 20516 7343 20519
rect 7926 20516 7932 20528
rect 7331 20488 7932 20516
rect 7331 20485 7343 20488
rect 7285 20479 7343 20485
rect 7926 20476 7932 20488
rect 7984 20476 7990 20528
rect 13265 20519 13323 20525
rect 8680 20488 9996 20516
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 8680 20457 8708 20488
rect 9674 20457 9680 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 7116 20420 8677 20448
rect 2222 20340 2228 20392
rect 2280 20340 2286 20392
rect 7116 20389 7144 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 9668 20411 9680 20457
rect 9674 20408 9680 20411
rect 9732 20408 9738 20460
rect 9968 20448 9996 20488
rect 13265 20485 13277 20519
rect 13311 20516 13323 20519
rect 14016 20516 14044 20544
rect 13311 20488 14044 20516
rect 13311 20485 13323 20488
rect 13265 20479 13323 20485
rect 10410 20448 10416 20460
rect 9968 20420 10416 20448
rect 10410 20408 10416 20420
rect 10468 20448 10474 20460
rect 14642 20448 14648 20460
rect 10468 20420 14648 20448
rect 10468 20408 10474 20420
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15102 20408 15108 20460
rect 15160 20408 15166 20460
rect 15273 20448 15301 20544
rect 16390 20476 16396 20528
rect 16448 20516 16454 20528
rect 18046 20516 18052 20528
rect 16448 20488 18052 20516
rect 16448 20476 16454 20488
rect 18046 20476 18052 20488
rect 18104 20476 18110 20528
rect 19610 20476 19616 20528
rect 19668 20525 19674 20528
rect 19668 20516 19680 20525
rect 19668 20488 19713 20516
rect 19668 20479 19680 20488
rect 19668 20476 19674 20479
rect 21174 20476 21180 20528
rect 21232 20516 21238 20528
rect 24136 20516 24164 20556
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 25869 20587 25927 20593
rect 25869 20553 25881 20587
rect 25915 20584 25927 20587
rect 26326 20584 26332 20596
rect 25915 20556 26332 20584
rect 25915 20553 25927 20556
rect 25869 20547 25927 20553
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 26694 20544 26700 20596
rect 26752 20584 26758 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 26752 20556 27261 20584
rect 26752 20544 26758 20556
rect 27249 20553 27261 20556
rect 27295 20553 27307 20587
rect 27249 20547 27307 20553
rect 29641 20587 29699 20593
rect 29641 20553 29653 20587
rect 29687 20584 29699 20587
rect 29730 20584 29736 20596
rect 29687 20556 29736 20584
rect 29687 20553 29699 20556
rect 29641 20547 29699 20553
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 30009 20587 30067 20593
rect 30009 20553 30021 20587
rect 30055 20584 30067 20587
rect 30561 20587 30619 20593
rect 30561 20584 30573 20587
rect 30055 20556 30573 20584
rect 30055 20553 30067 20556
rect 30009 20547 30067 20553
rect 30561 20553 30573 20556
rect 30607 20584 30619 20587
rect 30926 20584 30932 20596
rect 30607 20556 30932 20584
rect 30607 20553 30619 20556
rect 30561 20547 30619 20553
rect 30926 20544 30932 20556
rect 30984 20544 30990 20596
rect 38102 20544 38108 20596
rect 38160 20584 38166 20596
rect 38746 20584 38752 20596
rect 38160 20556 38752 20584
rect 38160 20544 38166 20556
rect 38746 20544 38752 20556
rect 38804 20544 38810 20596
rect 38841 20587 38899 20593
rect 38841 20553 38853 20587
rect 38887 20584 38899 20587
rect 38930 20584 38936 20596
rect 38887 20556 38936 20584
rect 38887 20553 38899 20556
rect 38841 20547 38899 20553
rect 38930 20544 38936 20556
rect 38988 20544 38994 20596
rect 42886 20544 42892 20596
rect 42944 20584 42950 20596
rect 43714 20584 43720 20596
rect 42944 20556 43720 20584
rect 42944 20544 42950 20556
rect 43714 20544 43720 20556
rect 43772 20544 43778 20596
rect 44726 20544 44732 20596
rect 44784 20544 44790 20596
rect 48133 20587 48191 20593
rect 48133 20553 48145 20587
rect 48179 20584 48191 20587
rect 48406 20584 48412 20596
rect 48179 20556 48412 20584
rect 48179 20553 48191 20556
rect 48133 20547 48191 20553
rect 48406 20544 48412 20556
rect 48464 20544 48470 20596
rect 51169 20587 51227 20593
rect 51169 20553 51181 20587
rect 51215 20584 51227 20587
rect 52178 20584 52184 20596
rect 51215 20556 52184 20584
rect 51215 20553 51227 20556
rect 51169 20547 51227 20553
rect 52178 20544 52184 20556
rect 52236 20544 52242 20596
rect 53558 20544 53564 20596
rect 53616 20544 53622 20596
rect 54018 20544 54024 20596
rect 54076 20544 54082 20596
rect 54757 20587 54815 20593
rect 54757 20553 54769 20587
rect 54803 20584 54815 20587
rect 55766 20584 55772 20596
rect 54803 20556 55772 20584
rect 54803 20553 54815 20556
rect 54757 20547 54815 20553
rect 55766 20544 55772 20556
rect 55824 20544 55830 20596
rect 57057 20587 57115 20593
rect 57057 20553 57069 20587
rect 57103 20584 57115 20587
rect 57422 20584 57428 20596
rect 57103 20556 57428 20584
rect 57103 20553 57115 20556
rect 57057 20547 57115 20553
rect 57422 20544 57428 20556
rect 57480 20544 57486 20596
rect 21232 20488 24164 20516
rect 24204 20519 24262 20525
rect 21232 20476 21238 20488
rect 24204 20485 24216 20519
rect 24250 20516 24262 20519
rect 24578 20516 24584 20528
rect 24250 20488 24584 20516
rect 24250 20485 24262 20488
rect 24204 20479 24262 20485
rect 24578 20476 24584 20488
rect 24636 20476 24642 20528
rect 25406 20476 25412 20528
rect 25464 20516 25470 20528
rect 28074 20516 28080 20528
rect 25464 20488 28080 20516
rect 25464 20476 25470 20488
rect 28074 20476 28080 20488
rect 28132 20476 28138 20528
rect 37553 20519 37611 20525
rect 37553 20485 37565 20519
rect 37599 20516 37611 20519
rect 38654 20516 38660 20528
rect 37599 20488 38660 20516
rect 37599 20485 37611 20488
rect 37553 20479 37611 20485
rect 38654 20476 38660 20488
rect 38712 20476 38718 20528
rect 39200 20519 39258 20525
rect 39200 20485 39212 20519
rect 39246 20516 39258 20519
rect 40218 20516 40224 20528
rect 39246 20488 40224 20516
rect 39246 20485 39258 20488
rect 39200 20479 39258 20485
rect 40218 20476 40224 20488
rect 40276 20476 40282 20528
rect 42978 20476 42984 20528
rect 43036 20516 43042 20528
rect 44821 20519 44879 20525
rect 44821 20516 44833 20519
rect 43036 20488 44833 20516
rect 43036 20476 43042 20488
rect 44821 20485 44833 20488
rect 44867 20485 44879 20519
rect 44821 20479 44879 20485
rect 48225 20519 48283 20525
rect 48225 20485 48237 20519
rect 48271 20516 48283 20519
rect 49418 20516 49424 20528
rect 48271 20488 49424 20516
rect 48271 20485 48283 20488
rect 48225 20479 48283 20485
rect 49418 20476 49424 20488
rect 49476 20476 49482 20528
rect 50154 20476 50160 20528
rect 50212 20516 50218 20528
rect 58066 20516 58072 20528
rect 50212 20488 52592 20516
rect 50212 20476 50218 20488
rect 15361 20451 15419 20457
rect 15361 20448 15373 20451
rect 15273 20420 15373 20448
rect 15361 20417 15373 20420
rect 15407 20417 15419 20451
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 15361 20411 15419 20417
rect 17880 20420 19901 20448
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20380 7251 20383
rect 7466 20380 7472 20392
rect 7239 20352 7472 20380
rect 7239 20349 7251 20352
rect 7193 20343 7251 20349
rect 7466 20340 7472 20352
rect 7524 20340 7530 20392
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 7653 20315 7711 20321
rect 7653 20281 7665 20315
rect 7699 20312 7711 20315
rect 8312 20312 8340 20343
rect 9030 20340 9036 20392
rect 9088 20380 9094 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 9088 20352 9413 20380
rect 9088 20340 9094 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 10928 20352 12817 20380
rect 10928 20340 10934 20352
rect 12805 20349 12817 20352
rect 12851 20380 12863 20383
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12851 20352 13093 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13219 20352 13737 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14550 20380 14556 20392
rect 14415 20352 14556 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 7699 20284 8340 20312
rect 13096 20312 13124 20343
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 16942 20340 16948 20392
rect 17000 20340 17006 20392
rect 13096 20284 14780 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 2866 20204 2872 20256
rect 2924 20204 2930 20256
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 13170 20244 13176 20256
rect 11756 20216 13176 20244
rect 11756 20204 11762 20216
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 14752 20244 14780 20284
rect 17880 20256 17908 20420
rect 19889 20417 19901 20420
rect 19935 20448 19947 20451
rect 20530 20448 20536 20460
rect 19935 20420 20536 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 21266 20408 21272 20460
rect 21324 20448 21330 20460
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21324 20420 22201 20448
rect 21324 20408 21330 20420
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20448 25835 20451
rect 26050 20448 26056 20460
rect 25823 20420 26056 20448
rect 25823 20417 25835 20420
rect 25777 20411 25835 20417
rect 26050 20408 26056 20420
rect 26108 20408 26114 20460
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 27341 20451 27399 20457
rect 27341 20448 27353 20451
rect 26476 20420 27353 20448
rect 26476 20408 26482 20420
rect 27341 20417 27353 20420
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 32493 20451 32551 20457
rect 32493 20417 32505 20451
rect 32539 20448 32551 20451
rect 33502 20448 33508 20460
rect 32539 20420 33508 20448
rect 32539 20417 32551 20420
rect 32493 20411 32551 20417
rect 33502 20408 33508 20420
rect 33560 20448 33566 20460
rect 33597 20451 33655 20457
rect 33597 20448 33609 20451
rect 33560 20420 33609 20448
rect 33560 20408 33566 20420
rect 33597 20417 33609 20420
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 33781 20451 33839 20457
rect 33781 20417 33793 20451
rect 33827 20448 33839 20451
rect 33870 20448 33876 20460
rect 33827 20420 33876 20448
rect 33827 20417 33839 20420
rect 33781 20411 33839 20417
rect 33870 20408 33876 20420
rect 33928 20408 33934 20460
rect 34048 20451 34106 20457
rect 34048 20417 34060 20451
rect 34094 20448 34106 20451
rect 35253 20451 35311 20457
rect 35253 20448 35265 20451
rect 34094 20420 35265 20448
rect 34094 20417 34106 20420
rect 34048 20411 34106 20417
rect 35253 20417 35265 20420
rect 35299 20417 35311 20451
rect 35253 20411 35311 20417
rect 37642 20408 37648 20460
rect 37700 20448 37706 20460
rect 38473 20451 38531 20457
rect 38473 20448 38485 20451
rect 37700 20420 38485 20448
rect 37700 20408 37706 20420
rect 38473 20417 38485 20420
rect 38519 20448 38531 20451
rect 38562 20448 38568 20460
rect 38519 20420 38568 20448
rect 38519 20417 38531 20420
rect 38473 20411 38531 20417
rect 38562 20408 38568 20420
rect 38620 20448 38626 20460
rect 40862 20448 40868 20460
rect 38620 20420 40868 20448
rect 38620 20408 38626 20420
rect 40862 20408 40868 20420
rect 40920 20408 40926 20460
rect 42797 20451 42855 20457
rect 41432 20420 42748 20448
rect 18230 20340 18236 20392
rect 18288 20340 18294 20392
rect 19978 20340 19984 20392
rect 20036 20340 20042 20392
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 22097 20383 22155 20389
rect 22097 20380 22109 20383
rect 22060 20352 22109 20380
rect 22060 20340 22066 20352
rect 22097 20349 22109 20352
rect 22143 20349 22155 20383
rect 22097 20343 22155 20349
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 23937 20383 23995 20389
rect 23937 20349 23949 20383
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 20438 20272 20444 20324
rect 20496 20312 20502 20324
rect 21450 20312 21456 20324
rect 20496 20284 21456 20312
rect 20496 20272 20502 20284
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 22649 20315 22707 20321
rect 22649 20281 22661 20315
rect 22695 20312 22707 20315
rect 23768 20312 23796 20343
rect 22695 20284 23796 20312
rect 22695 20281 22707 20284
rect 22649 20275 22707 20281
rect 23952 20256 23980 20343
rect 25222 20340 25228 20392
rect 25280 20340 25286 20392
rect 25958 20340 25964 20392
rect 26016 20340 26022 20392
rect 26602 20340 26608 20392
rect 26660 20380 26666 20392
rect 26789 20383 26847 20389
rect 26789 20380 26801 20383
rect 26660 20352 26801 20380
rect 26660 20340 26666 20352
rect 26789 20349 26801 20352
rect 26835 20380 26847 20383
rect 27065 20383 27123 20389
rect 27065 20380 27077 20383
rect 26835 20352 27077 20380
rect 26835 20349 26847 20352
rect 26789 20343 26847 20349
rect 27065 20349 27077 20352
rect 27111 20349 27123 20383
rect 27065 20343 27123 20349
rect 27246 20340 27252 20392
rect 27304 20380 27310 20392
rect 27801 20383 27859 20389
rect 27801 20380 27813 20383
rect 27304 20352 27813 20380
rect 27304 20340 27310 20352
rect 27801 20349 27813 20352
rect 27847 20349 27859 20383
rect 27801 20343 27859 20349
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 30101 20383 30159 20389
rect 30101 20380 30113 20383
rect 29052 20352 30113 20380
rect 29052 20340 29058 20352
rect 30101 20349 30113 20352
rect 30147 20349 30159 20383
rect 30101 20343 30159 20349
rect 30193 20383 30251 20389
rect 30193 20349 30205 20383
rect 30239 20349 30251 20383
rect 30193 20343 30251 20349
rect 25240 20312 25268 20340
rect 25409 20315 25467 20321
rect 25409 20312 25421 20315
rect 25240 20284 25421 20312
rect 25409 20281 25421 20284
rect 25455 20281 25467 20315
rect 30208 20312 30236 20343
rect 31110 20340 31116 20392
rect 31168 20340 31174 20392
rect 31941 20383 31999 20389
rect 31941 20349 31953 20383
rect 31987 20349 31999 20383
rect 31941 20343 31999 20349
rect 25409 20275 25467 20281
rect 29472 20284 30236 20312
rect 31956 20312 31984 20343
rect 32582 20340 32588 20392
rect 32640 20340 32646 20392
rect 32674 20340 32680 20392
rect 32732 20340 32738 20392
rect 32950 20340 32956 20392
rect 33008 20340 33014 20392
rect 35802 20340 35808 20392
rect 35860 20340 35866 20392
rect 36541 20383 36599 20389
rect 36541 20349 36553 20383
rect 36587 20349 36599 20383
rect 36541 20343 36599 20349
rect 32125 20315 32183 20321
rect 32125 20312 32137 20315
rect 31956 20284 32137 20312
rect 29472 20256 29500 20284
rect 32125 20281 32137 20284
rect 32171 20281 32183 20315
rect 32125 20275 32183 20281
rect 15286 20244 15292 20256
rect 14752 20216 15292 20244
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 17586 20204 17592 20256
rect 17644 20244 17650 20256
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17644 20216 17693 20244
rect 17644 20204 17650 20216
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 17862 20204 17868 20256
rect 17920 20204 17926 20256
rect 19702 20204 19708 20256
rect 19760 20244 19766 20256
rect 20625 20247 20683 20253
rect 20625 20244 20637 20247
rect 19760 20216 20637 20244
rect 19760 20204 19766 20216
rect 20625 20213 20637 20216
rect 20671 20244 20683 20247
rect 21542 20244 21548 20256
rect 20671 20216 21548 20244
rect 20671 20213 20683 20216
rect 20625 20207 20683 20213
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 21637 20247 21695 20253
rect 21637 20213 21649 20247
rect 21683 20244 21695 20247
rect 21818 20244 21824 20256
rect 21683 20216 21824 20244
rect 21683 20213 21695 20216
rect 21637 20207 21695 20213
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 23198 20204 23204 20256
rect 23256 20204 23262 20256
rect 23934 20204 23940 20256
rect 23992 20204 23998 20256
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 26142 20244 26148 20256
rect 24912 20216 26148 20244
rect 24912 20204 24918 20216
rect 26142 20204 26148 20216
rect 26200 20204 26206 20256
rect 27338 20204 27344 20256
rect 27396 20244 27402 20256
rect 27709 20247 27767 20253
rect 27709 20244 27721 20247
rect 27396 20216 27721 20244
rect 27396 20204 27402 20216
rect 27709 20213 27721 20216
rect 27755 20213 27767 20247
rect 27709 20207 27767 20213
rect 28442 20204 28448 20256
rect 28500 20204 28506 20256
rect 29454 20204 29460 20256
rect 29512 20204 29518 20256
rect 31297 20247 31355 20253
rect 31297 20213 31309 20247
rect 31343 20244 31355 20247
rect 31386 20244 31392 20256
rect 31343 20216 31392 20244
rect 31343 20213 31355 20216
rect 31297 20207 31355 20213
rect 31386 20204 31392 20216
rect 31444 20204 31450 20256
rect 32692 20244 32720 20340
rect 35161 20315 35219 20321
rect 35161 20281 35173 20315
rect 35207 20312 35219 20315
rect 36556 20312 36584 20343
rect 37458 20340 37464 20392
rect 37516 20380 37522 20392
rect 37826 20380 37832 20392
rect 37516 20352 37832 20380
rect 37516 20340 37522 20352
rect 37826 20340 37832 20352
rect 37884 20340 37890 20392
rect 38102 20340 38108 20392
rect 38160 20380 38166 20392
rect 38197 20383 38255 20389
rect 38197 20380 38209 20383
rect 38160 20352 38209 20380
rect 38160 20340 38166 20352
rect 38197 20349 38209 20352
rect 38243 20349 38255 20383
rect 38197 20343 38255 20349
rect 38381 20383 38439 20389
rect 38381 20349 38393 20383
rect 38427 20380 38439 20383
rect 38838 20380 38844 20392
rect 38427 20352 38844 20380
rect 38427 20349 38439 20352
rect 38381 20343 38439 20349
rect 38838 20340 38844 20352
rect 38896 20340 38902 20392
rect 38933 20383 38991 20389
rect 38933 20349 38945 20383
rect 38979 20349 38991 20383
rect 40405 20383 40463 20389
rect 40405 20380 40417 20383
rect 38933 20343 38991 20349
rect 40328 20352 40417 20380
rect 35207 20284 36584 20312
rect 35207 20281 35219 20284
rect 35161 20275 35219 20281
rect 36906 20272 36912 20324
rect 36964 20312 36970 20324
rect 38948 20312 38976 20343
rect 40328 20321 40356 20352
rect 40405 20349 40417 20352
rect 40451 20349 40463 20383
rect 40405 20343 40463 20349
rect 36964 20284 38976 20312
rect 36964 20272 36970 20284
rect 35710 20244 35716 20256
rect 32692 20216 35716 20244
rect 35710 20204 35716 20216
rect 35768 20204 35774 20256
rect 35986 20204 35992 20256
rect 36044 20204 36050 20256
rect 37093 20247 37151 20253
rect 37093 20213 37105 20247
rect 37139 20244 37151 20247
rect 37826 20244 37832 20256
rect 37139 20216 37832 20244
rect 37139 20213 37151 20216
rect 37093 20207 37151 20213
rect 37826 20204 37832 20216
rect 37884 20204 37890 20256
rect 38010 20204 38016 20256
rect 38068 20204 38074 20256
rect 38948 20244 38976 20284
rect 40313 20315 40371 20321
rect 40313 20281 40325 20315
rect 40359 20281 40371 20315
rect 40313 20275 40371 20281
rect 41432 20256 41460 20420
rect 42245 20383 42303 20389
rect 42245 20349 42257 20383
rect 42291 20349 42303 20383
rect 42720 20380 42748 20420
rect 42797 20417 42809 20451
rect 42843 20448 42855 20451
rect 43806 20448 43812 20460
rect 42843 20420 43812 20448
rect 42843 20417 42855 20420
rect 42797 20411 42855 20417
rect 43806 20408 43812 20420
rect 43864 20448 43870 20460
rect 43901 20451 43959 20457
rect 43901 20448 43913 20451
rect 43864 20420 43913 20448
rect 43864 20408 43870 20420
rect 43901 20417 43913 20420
rect 43947 20417 43959 20451
rect 46750 20448 46756 20460
rect 43901 20411 43959 20417
rect 44376 20420 46756 20448
rect 42981 20383 43039 20389
rect 42981 20380 42993 20383
rect 42720 20352 42993 20380
rect 42245 20343 42303 20349
rect 42981 20349 42993 20352
rect 43027 20349 43039 20383
rect 42981 20343 43039 20349
rect 42260 20312 42288 20343
rect 42429 20315 42487 20321
rect 42429 20312 42441 20315
rect 42260 20284 42441 20312
rect 42429 20281 42441 20284
rect 42475 20281 42487 20315
rect 42996 20312 43024 20343
rect 43254 20340 43260 20392
rect 43312 20340 43318 20392
rect 44376 20380 44404 20420
rect 46750 20408 46756 20420
rect 46808 20408 46814 20460
rect 52564 20457 52592 20488
rect 56612 20488 58072 20516
rect 52293 20451 52351 20457
rect 52293 20417 52305 20451
rect 52339 20448 52351 20451
rect 52549 20451 52607 20457
rect 52339 20420 52500 20448
rect 52339 20417 52351 20420
rect 52293 20411 52351 20417
rect 43548 20352 44404 20380
rect 43548 20312 43576 20352
rect 44450 20340 44456 20392
rect 44508 20380 44514 20392
rect 44545 20383 44603 20389
rect 44545 20380 44557 20383
rect 44508 20352 44557 20380
rect 44508 20340 44514 20352
rect 44545 20349 44557 20352
rect 44591 20380 44603 20383
rect 44634 20380 44640 20392
rect 44591 20352 44640 20380
rect 44591 20349 44603 20352
rect 44545 20343 44603 20349
rect 44634 20340 44640 20352
rect 44692 20340 44698 20392
rect 45278 20340 45284 20392
rect 45336 20340 45342 20392
rect 46017 20383 46075 20389
rect 46017 20349 46029 20383
rect 46063 20349 46075 20383
rect 48317 20383 48375 20389
rect 48317 20380 48329 20383
rect 46017 20343 46075 20349
rect 47320 20352 48329 20380
rect 42996 20284 43576 20312
rect 42429 20275 42487 20281
rect 43622 20272 43628 20324
rect 43680 20312 43686 20324
rect 43990 20312 43996 20324
rect 43680 20284 43996 20312
rect 43680 20272 43686 20284
rect 43990 20272 43996 20284
rect 44048 20312 44054 20324
rect 44818 20312 44824 20324
rect 44048 20284 44824 20312
rect 44048 20272 44054 20284
rect 44818 20272 44824 20284
rect 44876 20272 44882 20324
rect 45189 20315 45247 20321
rect 45189 20281 45201 20315
rect 45235 20312 45247 20315
rect 46032 20312 46060 20343
rect 45235 20284 46060 20312
rect 45235 20281 45247 20284
rect 45189 20275 45247 20281
rect 47320 20256 47348 20352
rect 48317 20349 48329 20352
rect 48363 20349 48375 20383
rect 48317 20343 48375 20349
rect 49142 20340 49148 20392
rect 49200 20340 49206 20392
rect 52472 20380 52500 20420
rect 52549 20417 52561 20451
rect 52595 20448 52607 20451
rect 52730 20448 52736 20460
rect 52595 20420 52736 20448
rect 52595 20417 52607 20420
rect 52549 20411 52607 20417
rect 52730 20408 52736 20420
rect 52788 20408 52794 20460
rect 53929 20451 53987 20457
rect 53929 20417 53941 20451
rect 53975 20417 53987 20451
rect 53929 20411 53987 20417
rect 53285 20383 53343 20389
rect 52472 20352 52776 20380
rect 47486 20272 47492 20324
rect 47544 20312 47550 20324
rect 52748 20321 52776 20352
rect 53285 20349 53297 20383
rect 53331 20349 53343 20383
rect 53285 20343 53343 20349
rect 48593 20315 48651 20321
rect 48593 20312 48605 20315
rect 47544 20284 48605 20312
rect 47544 20272 47550 20284
rect 48593 20281 48605 20284
rect 48639 20281 48651 20315
rect 48593 20275 48651 20281
rect 52733 20315 52791 20321
rect 52733 20281 52745 20315
rect 52779 20281 52791 20315
rect 52733 20275 52791 20281
rect 39114 20244 39120 20256
rect 38948 20216 39120 20244
rect 39114 20204 39120 20216
rect 39172 20204 39178 20256
rect 41046 20204 41052 20256
rect 41104 20204 41110 20256
rect 41414 20204 41420 20256
rect 41472 20204 41478 20256
rect 41601 20247 41659 20253
rect 41601 20213 41613 20247
rect 41647 20244 41659 20247
rect 41690 20244 41696 20256
rect 41647 20216 41696 20244
rect 41647 20213 41659 20216
rect 41601 20207 41659 20213
rect 41690 20204 41696 20216
rect 41748 20204 41754 20256
rect 44361 20247 44419 20253
rect 44361 20213 44373 20247
rect 44407 20244 44419 20247
rect 45094 20244 45100 20256
rect 44407 20216 45100 20244
rect 44407 20213 44419 20216
rect 44361 20207 44419 20213
rect 45094 20204 45100 20216
rect 45152 20204 45158 20256
rect 45922 20204 45928 20256
rect 45980 20204 45986 20256
rect 46658 20204 46664 20256
rect 46716 20204 46722 20256
rect 47302 20204 47308 20256
rect 47360 20204 47366 20256
rect 47765 20247 47823 20253
rect 47765 20213 47777 20247
rect 47811 20244 47823 20247
rect 47854 20244 47860 20256
rect 47811 20216 47860 20244
rect 47811 20213 47823 20216
rect 47765 20207 47823 20213
rect 47854 20204 47860 20216
rect 47912 20204 47918 20256
rect 52362 20204 52368 20256
rect 52420 20244 52426 20256
rect 53300 20244 53328 20343
rect 52420 20216 53328 20244
rect 53944 20244 53972 20411
rect 55398 20408 55404 20460
rect 55456 20408 55462 20460
rect 56612 20457 56640 20488
rect 58066 20476 58072 20488
rect 58124 20516 58130 20528
rect 58529 20519 58587 20525
rect 58529 20516 58541 20519
rect 58124 20488 58541 20516
rect 58124 20476 58130 20488
rect 58529 20485 58541 20488
rect 58575 20485 58587 20519
rect 58529 20479 58587 20485
rect 56597 20451 56655 20457
rect 56597 20417 56609 20451
rect 56643 20417 56655 20451
rect 56597 20411 56655 20417
rect 57072 20420 57284 20448
rect 54018 20340 54024 20392
rect 54076 20380 54082 20392
rect 55582 20389 55588 20392
rect 54113 20383 54171 20389
rect 54113 20380 54125 20383
rect 54076 20352 54125 20380
rect 54076 20340 54082 20352
rect 54113 20349 54125 20352
rect 54159 20380 54171 20383
rect 54573 20383 54631 20389
rect 54573 20380 54585 20383
rect 54159 20352 54585 20380
rect 54159 20349 54171 20352
rect 54113 20343 54171 20349
rect 54573 20349 54585 20352
rect 54619 20349 54631 20383
rect 54573 20343 54631 20349
rect 55560 20383 55588 20389
rect 55560 20349 55572 20383
rect 55560 20343 55588 20349
rect 55582 20340 55588 20343
rect 55640 20340 55646 20392
rect 55677 20383 55735 20389
rect 55677 20349 55689 20383
rect 55723 20380 55735 20383
rect 55953 20383 56011 20389
rect 55723 20352 55904 20380
rect 55723 20349 55735 20352
rect 55677 20343 55735 20349
rect 54846 20272 54852 20324
rect 54904 20272 54910 20324
rect 54478 20244 54484 20256
rect 53944 20216 54484 20244
rect 52420 20204 52426 20216
rect 54478 20204 54484 20216
rect 54536 20204 54542 20256
rect 54864 20244 54892 20272
rect 55876 20244 55904 20352
rect 55953 20349 55965 20383
rect 55999 20380 56011 20383
rect 56042 20380 56048 20392
rect 55999 20352 56048 20380
rect 55999 20349 56011 20352
rect 55953 20343 56011 20349
rect 56042 20340 56048 20352
rect 56100 20340 56106 20392
rect 56318 20340 56324 20392
rect 56376 20340 56382 20392
rect 56413 20383 56471 20389
rect 56413 20349 56425 20383
rect 56459 20380 56471 20383
rect 56962 20380 56968 20392
rect 56459 20352 56968 20380
rect 56459 20349 56471 20352
rect 56413 20343 56471 20349
rect 56962 20340 56968 20352
rect 57020 20340 57026 20392
rect 56336 20312 56364 20340
rect 57072 20312 57100 20420
rect 57256 20389 57284 20420
rect 57514 20408 57520 20460
rect 57572 20448 57578 20460
rect 57885 20451 57943 20457
rect 57885 20448 57897 20451
rect 57572 20420 57897 20448
rect 57572 20408 57578 20420
rect 57885 20417 57897 20420
rect 57931 20417 57943 20451
rect 57885 20411 57943 20417
rect 57149 20383 57207 20389
rect 57149 20349 57161 20383
rect 57195 20349 57207 20383
rect 57149 20343 57207 20349
rect 57241 20383 57299 20389
rect 57241 20349 57253 20383
rect 57287 20349 57299 20383
rect 57241 20343 57299 20349
rect 56336 20284 57100 20312
rect 57164 20312 57192 20343
rect 57422 20312 57428 20324
rect 57164 20284 57428 20312
rect 57422 20272 57428 20284
rect 57480 20272 57486 20324
rect 54864 20216 55904 20244
rect 56686 20204 56692 20256
rect 56744 20204 56750 20256
rect 1104 20154 58880 20176
rect 1104 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 22616 20154
rect 22668 20102 22680 20154
rect 22732 20102 22744 20154
rect 22796 20102 22808 20154
rect 22860 20102 22872 20154
rect 22924 20102 37060 20154
rect 37112 20102 37124 20154
rect 37176 20102 37188 20154
rect 37240 20102 37252 20154
rect 37304 20102 37316 20154
rect 37368 20102 51504 20154
rect 51556 20102 51568 20154
rect 51620 20102 51632 20154
rect 51684 20102 51696 20154
rect 51748 20102 51760 20154
rect 51812 20102 58880 20154
rect 1104 20080 58880 20102
rect 9585 20043 9643 20049
rect 9585 20009 9597 20043
rect 9631 20040 9643 20043
rect 9674 20040 9680 20052
rect 9631 20012 9680 20040
rect 9631 20009 9643 20012
rect 9585 20003 9643 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 16942 20040 16948 20052
rect 16531 20012 16948 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 19058 20000 19064 20052
rect 19116 20000 19122 20052
rect 20533 20043 20591 20049
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 21082 20040 21088 20052
rect 20579 20012 21088 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 22462 20040 22468 20052
rect 21508 20012 21772 20040
rect 21508 20000 21514 20012
rect 13909 19975 13967 19981
rect 13909 19941 13921 19975
rect 13955 19972 13967 19975
rect 13955 19944 15516 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 7834 19904 7840 19916
rect 7432 19876 7840 19904
rect 7432 19864 7438 19876
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 10229 19907 10287 19913
rect 10229 19873 10241 19907
rect 10275 19904 10287 19907
rect 10275 19876 10916 19904
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 2130 19796 2136 19848
rect 2188 19796 2194 19848
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 2869 19839 2927 19845
rect 2869 19836 2881 19839
rect 2832 19808 2881 19836
rect 2832 19796 2838 19808
rect 2869 19805 2881 19808
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 3418 19796 3424 19848
rect 3476 19796 3482 19848
rect 3510 19796 3516 19848
rect 3568 19836 3574 19848
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3568 19808 3801 19836
rect 3568 19796 3574 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 6914 19796 6920 19848
rect 6972 19796 6978 19848
rect 7558 19796 7564 19848
rect 7616 19796 7622 19848
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9824 19808 9965 19836
rect 9824 19796 9830 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 6270 19768 6276 19780
rect 3988 19740 6276 19768
rect 3988 19712 4016 19740
rect 6270 19728 6276 19740
rect 6328 19728 6334 19780
rect 10888 19712 10916 19876
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 15488 19913 15516 19944
rect 19518 19932 19524 19984
rect 19576 19972 19582 19984
rect 21744 19981 21772 20012
rect 22204 20012 22468 20040
rect 21729 19975 21787 19981
rect 19576 19944 20668 19972
rect 19576 19932 19582 19944
rect 15473 19907 15531 19913
rect 14700 19876 15424 19904
rect 14700 19864 14706 19876
rect 12526 19796 12532 19848
rect 12584 19796 12590 19848
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 14516 19808 14933 19836
rect 14516 19796 14522 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 15396 19836 15424 19876
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 17862 19864 17868 19916
rect 17920 19864 17926 19916
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 18598 19904 18604 19916
rect 18555 19876 18604 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18708 19876 19656 19904
rect 17034 19836 17040 19848
rect 15396 19808 17040 19836
rect 14921 19799 14979 19805
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 17586 19796 17592 19848
rect 17644 19845 17650 19848
rect 17644 19836 17656 19845
rect 18708 19836 18736 19876
rect 19518 19836 19524 19848
rect 17644 19808 17689 19836
rect 18156 19808 18736 19836
rect 18892 19808 19524 19836
rect 17644 19799 17656 19808
rect 17644 19796 17650 19799
rect 12796 19771 12854 19777
rect 12796 19737 12808 19771
rect 12842 19768 12854 19771
rect 13354 19768 13360 19780
rect 12842 19740 13360 19768
rect 12842 19737 12854 19740
rect 12796 19731 12854 19737
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 13740 19740 14565 19768
rect 13740 19712 13768 19740
rect 14553 19737 14565 19740
rect 14599 19737 14611 19771
rect 14553 19731 14611 19737
rect 2777 19703 2835 19709
rect 2777 19669 2789 19703
rect 2823 19700 2835 19703
rect 2958 19700 2964 19712
rect 2823 19672 2964 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 3970 19660 3976 19712
rect 4028 19660 4034 19712
rect 4433 19703 4491 19709
rect 4433 19669 4445 19703
rect 4479 19700 4491 19703
rect 4522 19700 4528 19712
rect 4479 19672 4528 19700
rect 4479 19669 4491 19672
rect 4433 19663 4491 19669
rect 4522 19660 4528 19672
rect 4580 19660 4586 19712
rect 7006 19660 7012 19712
rect 7064 19660 7070 19712
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7926 19700 7932 19712
rect 7432 19672 7932 19700
rect 7432 19660 7438 19672
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 10042 19660 10048 19712
rect 10100 19660 10106 19712
rect 10594 19660 10600 19712
rect 10652 19660 10658 19712
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 10965 19703 11023 19709
rect 10965 19700 10977 19703
rect 10928 19672 10977 19700
rect 10928 19660 10934 19672
rect 10965 19669 10977 19672
rect 11011 19669 11023 19703
rect 10965 19663 11023 19669
rect 13722 19660 13728 19712
rect 13780 19660 13786 19712
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 18156 19709 18184 19808
rect 18601 19771 18659 19777
rect 18601 19737 18613 19771
rect 18647 19768 18659 19771
rect 18782 19768 18788 19780
rect 18647 19740 18788 19768
rect 18647 19737 18659 19740
rect 18601 19731 18659 19737
rect 18782 19728 18788 19740
rect 18840 19728 18846 19780
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 18104 19672 18153 19700
rect 18104 19660 18110 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 18892 19700 18920 19808
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 19628 19836 19656 19876
rect 19702 19864 19708 19916
rect 19760 19864 19766 19916
rect 19797 19907 19855 19913
rect 19797 19873 19809 19907
rect 19843 19873 19855 19907
rect 19797 19867 19855 19873
rect 19812 19836 19840 19867
rect 20530 19864 20536 19916
rect 20588 19864 20594 19916
rect 20640 19904 20668 19944
rect 21729 19941 21741 19975
rect 21775 19972 21787 19975
rect 21775 19944 22094 19972
rect 21775 19941 21787 19944
rect 21729 19935 21787 19941
rect 21336 19907 21394 19913
rect 21336 19904 21348 19907
rect 20640 19876 21348 19904
rect 21336 19873 21348 19876
rect 21382 19873 21394 19907
rect 21336 19867 21394 19873
rect 21450 19864 21456 19916
rect 21508 19864 21514 19916
rect 19628 19808 19840 19836
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 20548 19768 20576 19864
rect 21174 19796 21180 19848
rect 21232 19796 21238 19848
rect 22066 19836 22094 19944
rect 22204 19913 22232 20012
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23716 20012 23857 20040
rect 23716 20000 23722 20012
rect 23845 20009 23857 20012
rect 23891 20009 23903 20043
rect 23845 20003 23903 20009
rect 24673 20043 24731 20049
rect 24673 20009 24685 20043
rect 24719 20040 24731 20043
rect 24854 20040 24860 20052
rect 24719 20012 24860 20040
rect 24719 20009 24731 20012
rect 24673 20003 24731 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 25593 20043 25651 20049
rect 25593 20009 25605 20043
rect 25639 20040 25651 20043
rect 26418 20040 26424 20052
rect 25639 20012 26424 20040
rect 25639 20009 25651 20012
rect 25593 20003 25651 20009
rect 26418 20000 26424 20012
rect 26476 20000 26482 20052
rect 27522 20000 27528 20052
rect 27580 20000 27586 20052
rect 30929 20043 30987 20049
rect 30929 20009 30941 20043
rect 30975 20040 30987 20043
rect 31110 20040 31116 20052
rect 30975 20012 31116 20040
rect 30975 20009 30987 20012
rect 30929 20003 30987 20009
rect 31110 20000 31116 20012
rect 31168 20000 31174 20052
rect 32493 20043 32551 20049
rect 32493 20009 32505 20043
rect 32539 20040 32551 20043
rect 32950 20040 32956 20052
rect 32539 20012 32956 20040
rect 32539 20009 32551 20012
rect 32493 20003 32551 20009
rect 32950 20000 32956 20012
rect 33008 20000 33014 20052
rect 35437 20043 35495 20049
rect 35437 20009 35449 20043
rect 35483 20040 35495 20043
rect 35802 20040 35808 20052
rect 35483 20012 35808 20040
rect 35483 20009 35495 20012
rect 35437 20003 35495 20009
rect 35802 20000 35808 20012
rect 35860 20000 35866 20052
rect 35986 20000 35992 20052
rect 36044 20000 36050 20052
rect 37461 20043 37519 20049
rect 37461 20009 37473 20043
rect 37507 20040 37519 20043
rect 37734 20040 37740 20052
rect 37507 20012 37740 20040
rect 37507 20009 37519 20012
rect 37461 20003 37519 20009
rect 37734 20000 37740 20012
rect 37792 20000 37798 20052
rect 38838 20000 38844 20052
rect 38896 20000 38902 20052
rect 39114 20000 39120 20052
rect 39172 20040 39178 20052
rect 42797 20043 42855 20049
rect 39172 20012 41460 20040
rect 39172 20000 39178 20012
rect 22296 19944 22508 19972
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 22296 19836 22324 19944
rect 22370 19864 22376 19916
rect 22428 19864 22434 19916
rect 22480 19904 22508 19944
rect 26786 19932 26792 19984
rect 26844 19932 26850 19984
rect 33873 19975 33931 19981
rect 33873 19941 33885 19975
rect 33919 19972 33931 19975
rect 35618 19972 35624 19984
rect 33919 19944 35624 19972
rect 33919 19941 33931 19944
rect 33873 19935 33931 19941
rect 35618 19932 35624 19944
rect 35676 19972 35682 19984
rect 35676 19944 35848 19972
rect 35676 19932 35682 19944
rect 35820 19916 35848 19944
rect 22480 19876 22600 19904
rect 22066 19808 22324 19836
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 19024 19740 20484 19768
rect 20548 19740 20760 19768
rect 19024 19728 19030 19740
rect 18739 19672 18920 19700
rect 19245 19703 19303 19709
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 19245 19669 19257 19703
rect 19291 19700 19303 19703
rect 19518 19700 19524 19712
rect 19291 19672 19524 19700
rect 19291 19669 19303 19672
rect 19245 19663 19303 19669
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 19628 19709 19656 19740
rect 19613 19703 19671 19709
rect 19613 19669 19625 19703
rect 19659 19669 19671 19703
rect 19613 19663 19671 19669
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20349 19703 20407 19709
rect 20349 19700 20361 19703
rect 19944 19672 20361 19700
rect 19944 19660 19950 19672
rect 20349 19669 20361 19672
rect 20395 19669 20407 19703
rect 20456 19700 20484 19740
rect 20622 19700 20628 19712
rect 20456 19672 20628 19700
rect 20349 19663 20407 19669
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 20732 19700 20760 19740
rect 21726 19700 21732 19712
rect 20732 19672 21732 19700
rect 21726 19660 21732 19672
rect 21784 19700 21790 19712
rect 22480 19700 22508 19799
rect 22572 19768 22600 19876
rect 25406 19864 25412 19916
rect 25464 19864 25470 19916
rect 26050 19864 26056 19916
rect 26108 19904 26114 19916
rect 26375 19907 26433 19913
rect 26375 19904 26387 19907
rect 26108 19876 26387 19904
rect 26108 19864 26114 19876
rect 26375 19873 26387 19876
rect 26421 19873 26433 19907
rect 26375 19867 26433 19873
rect 26510 19864 26516 19916
rect 26568 19864 26574 19916
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 26878 19904 26884 19916
rect 26752 19876 26884 19904
rect 26752 19864 26758 19876
rect 26878 19864 26884 19876
rect 26936 19904 26942 19916
rect 27249 19907 27307 19913
rect 26936 19876 27108 19904
rect 26936 19864 26942 19876
rect 22732 19839 22790 19845
rect 22732 19805 22744 19839
rect 22778 19836 22790 19839
rect 23198 19836 23204 19848
rect 22778 19808 23204 19836
rect 22778 19805 22790 19808
rect 22732 19799 22790 19805
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 26234 19796 26240 19848
rect 26292 19796 26298 19848
rect 27080 19836 27108 19876
rect 27249 19873 27261 19907
rect 27295 19904 27307 19907
rect 27798 19904 27804 19916
rect 27295 19876 27804 19904
rect 27295 19873 27307 19876
rect 27249 19867 27307 19873
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 33318 19864 33324 19916
rect 33376 19864 33382 19916
rect 33502 19913 33508 19916
rect 33480 19907 33508 19913
rect 33480 19873 33492 19907
rect 33480 19867 33508 19873
rect 33502 19864 33508 19867
rect 33560 19864 33566 19916
rect 34333 19907 34391 19913
rect 34333 19873 34345 19907
rect 34379 19904 34391 19907
rect 34379 19876 34744 19904
rect 34379 19873 34391 19876
rect 34333 19867 34391 19873
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27080 19808 27445 19836
rect 27433 19805 27445 19808
rect 27479 19805 27491 19839
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 27433 19799 27491 19805
rect 27540 19808 28917 19836
rect 24121 19771 24179 19777
rect 24121 19768 24133 19771
rect 22572 19740 24133 19768
rect 24121 19737 24133 19740
rect 24167 19768 24179 19771
rect 25038 19768 25044 19780
rect 24167 19740 25044 19768
rect 24167 19737 24179 19740
rect 24121 19731 24179 19737
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 27540 19768 27568 19808
rect 28905 19805 28917 19808
rect 28951 19836 28963 19839
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 28951 19808 29561 19836
rect 28951 19805 28963 19808
rect 28905 19799 28963 19805
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29549 19799 29607 19805
rect 29816 19839 29874 19845
rect 29816 19805 29828 19839
rect 29862 19836 29874 19839
rect 30374 19836 30380 19848
rect 29862 19808 30380 19836
rect 29862 19805 29874 19808
rect 29816 19799 29874 19805
rect 30374 19796 30380 19808
rect 30432 19796 30438 19848
rect 31386 19845 31392 19848
rect 31113 19839 31171 19845
rect 31113 19805 31125 19839
rect 31159 19805 31171 19839
rect 31380 19836 31392 19845
rect 31347 19808 31392 19836
rect 31113 19799 31171 19805
rect 31380 19799 31392 19808
rect 27448 19740 27568 19768
rect 21784 19672 22508 19700
rect 24765 19703 24823 19709
rect 21784 19660 21790 19672
rect 24765 19669 24777 19703
rect 24811 19700 24823 19703
rect 24946 19700 24952 19712
rect 24811 19672 24952 19700
rect 24811 19669 24823 19672
rect 24765 19663 24823 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 25130 19660 25136 19712
rect 25188 19660 25194 19712
rect 25225 19703 25283 19709
rect 25225 19669 25237 19703
rect 25271 19700 25283 19703
rect 26510 19700 26516 19712
rect 25271 19672 26516 19700
rect 25271 19669 25283 19672
rect 25225 19663 25283 19669
rect 26510 19660 26516 19672
rect 26568 19660 26574 19712
rect 26970 19660 26976 19712
rect 27028 19700 27034 19712
rect 27448 19700 27476 19740
rect 28442 19728 28448 19780
rect 28500 19768 28506 19780
rect 28638 19771 28696 19777
rect 28638 19768 28650 19771
rect 28500 19740 28650 19768
rect 28500 19728 28506 19740
rect 28638 19737 28650 19740
rect 28684 19737 28696 19771
rect 28638 19731 28696 19737
rect 31128 19712 31156 19799
rect 31386 19796 31392 19799
rect 31444 19796 31450 19848
rect 33594 19796 33600 19848
rect 33652 19796 33658 19848
rect 34514 19796 34520 19848
rect 34572 19796 34578 19848
rect 34716 19836 34744 19876
rect 34790 19864 34796 19916
rect 34848 19904 34854 19916
rect 35713 19907 35771 19913
rect 35713 19904 35725 19907
rect 34848 19876 35725 19904
rect 34848 19864 34854 19876
rect 35713 19873 35725 19876
rect 35759 19873 35771 19907
rect 35713 19867 35771 19873
rect 35802 19864 35808 19916
rect 35860 19864 35866 19916
rect 35069 19839 35127 19845
rect 35069 19836 35081 19839
rect 34716 19808 35081 19836
rect 35069 19805 35081 19808
rect 35115 19836 35127 19839
rect 36004 19836 36032 20000
rect 38856 19972 38884 20000
rect 40681 19975 40739 19981
rect 40681 19972 40693 19975
rect 38856 19944 40693 19972
rect 38194 19864 38200 19916
rect 38252 19904 38258 19916
rect 38381 19907 38439 19913
rect 38381 19904 38393 19907
rect 38252 19876 38393 19904
rect 38252 19864 38258 19876
rect 38381 19873 38393 19876
rect 38427 19873 38439 19907
rect 38381 19867 38439 19873
rect 38654 19864 38660 19916
rect 38712 19864 38718 19916
rect 38933 19907 38991 19913
rect 38933 19873 38945 19907
rect 38979 19904 38991 19907
rect 39022 19904 39028 19916
rect 38979 19876 39028 19904
rect 38979 19873 38991 19876
rect 38933 19867 38991 19873
rect 39022 19864 39028 19876
rect 39080 19864 39086 19916
rect 35115 19808 36032 19836
rect 36081 19839 36139 19845
rect 35115 19805 35127 19808
rect 35069 19799 35127 19805
rect 36081 19805 36093 19839
rect 36127 19836 36139 19839
rect 36170 19836 36176 19848
rect 36127 19808 36176 19836
rect 36127 19805 36139 19808
rect 36081 19799 36139 19805
rect 36170 19796 36176 19808
rect 36228 19836 36234 19848
rect 36906 19836 36912 19848
rect 36228 19808 36912 19836
rect 36228 19796 36234 19808
rect 36906 19796 36912 19808
rect 36964 19796 36970 19848
rect 38470 19796 38476 19848
rect 38528 19845 38534 19848
rect 38528 19839 38577 19845
rect 38528 19805 38531 19839
rect 38565 19805 38577 19839
rect 39316 19836 39344 19944
rect 40681 19941 40693 19944
rect 40727 19941 40739 19975
rect 40681 19935 40739 19941
rect 39393 19907 39451 19913
rect 39393 19873 39405 19907
rect 39439 19904 39451 19907
rect 39439 19876 39988 19904
rect 39439 19873 39451 19876
rect 39393 19867 39451 19873
rect 39577 19839 39635 19845
rect 39577 19836 39589 19839
rect 39316 19808 39589 19836
rect 38528 19799 38577 19805
rect 39577 19805 39589 19808
rect 39623 19805 39635 19839
rect 39960 19836 39988 19876
rect 40034 19864 40040 19916
rect 40092 19904 40098 19916
rect 40313 19907 40371 19913
rect 40313 19904 40325 19907
rect 40092 19876 40325 19904
rect 40092 19864 40098 19876
rect 40313 19873 40325 19876
rect 40359 19873 40371 19907
rect 40313 19867 40371 19873
rect 40402 19864 40408 19916
rect 40460 19904 40466 19916
rect 41432 19913 41460 20012
rect 42797 20009 42809 20043
rect 42843 20040 42855 20043
rect 43254 20040 43260 20052
rect 42843 20012 43260 20040
rect 42843 20009 42855 20012
rect 42797 20003 42855 20009
rect 43254 20000 43260 20012
rect 43312 20000 43318 20052
rect 45005 20043 45063 20049
rect 45005 20009 45017 20043
rect 45051 20040 45063 20043
rect 45278 20040 45284 20052
rect 45051 20012 45284 20040
rect 45051 20009 45063 20012
rect 45005 20003 45063 20009
rect 45278 20000 45284 20012
rect 45336 20000 45342 20052
rect 48590 20000 48596 20052
rect 48648 20000 48654 20052
rect 48685 20043 48743 20049
rect 48685 20009 48697 20043
rect 48731 20040 48743 20043
rect 49142 20040 49148 20052
rect 48731 20012 49148 20040
rect 48731 20009 48743 20012
rect 48685 20003 48743 20009
rect 49142 20000 49148 20012
rect 49200 20000 49206 20052
rect 49789 20043 49847 20049
rect 49789 20009 49801 20043
rect 49835 20040 49847 20043
rect 49835 20012 51488 20040
rect 49835 20009 49847 20012
rect 49789 20003 49847 20009
rect 42978 19932 42984 19984
rect 43036 19932 43042 19984
rect 41417 19907 41475 19913
rect 40460 19876 41184 19904
rect 40460 19864 40466 19876
rect 41046 19836 41052 19848
rect 39960 19808 41052 19836
rect 39577 19799 39635 19805
rect 38528 19796 38534 19799
rect 41046 19796 41052 19808
rect 41104 19796 41110 19848
rect 36348 19771 36406 19777
rect 36348 19737 36360 19771
rect 36394 19768 36406 19771
rect 36722 19768 36728 19780
rect 36394 19740 36728 19768
rect 36394 19737 36406 19740
rect 36348 19731 36406 19737
rect 36722 19728 36728 19740
rect 36780 19728 36786 19780
rect 40221 19771 40279 19777
rect 40221 19768 40233 19771
rect 39408 19740 40233 19768
rect 27028 19672 27476 19700
rect 27028 19660 27034 19672
rect 31110 19660 31116 19712
rect 31168 19660 31174 19712
rect 32674 19660 32680 19712
rect 32732 19660 32738 19712
rect 34882 19660 34888 19712
rect 34940 19700 34946 19712
rect 34977 19703 35035 19709
rect 34977 19700 34989 19703
rect 34940 19672 34989 19700
rect 34940 19660 34946 19672
rect 34977 19669 34989 19672
rect 35023 19669 35035 19703
rect 34977 19663 35035 19669
rect 37737 19703 37795 19709
rect 37737 19669 37749 19703
rect 37783 19700 37795 19703
rect 39408 19700 39436 19740
rect 40221 19737 40233 19740
rect 40267 19737 40279 19771
rect 40221 19731 40279 19737
rect 37783 19672 39436 19700
rect 37783 19669 37795 19672
rect 37737 19663 37795 19669
rect 39850 19660 39856 19712
rect 39908 19660 39914 19712
rect 41156 19700 41184 19876
rect 41417 19873 41429 19907
rect 41463 19873 41475 19907
rect 41417 19867 41475 19873
rect 43622 19864 43628 19916
rect 43680 19864 43686 19916
rect 43806 19913 43812 19916
rect 43784 19907 43812 19913
rect 43784 19873 43796 19907
rect 43784 19867 43812 19873
rect 43806 19864 43812 19867
rect 43864 19864 43870 19916
rect 43898 19864 43904 19916
rect 43956 19864 43962 19916
rect 44177 19907 44235 19913
rect 44177 19873 44189 19907
rect 44223 19904 44235 19907
rect 44910 19904 44916 19916
rect 44223 19876 44916 19904
rect 44223 19873 44235 19876
rect 44177 19867 44235 19873
rect 44910 19864 44916 19876
rect 44968 19904 44974 19916
rect 46385 19907 46443 19913
rect 44968 19876 45416 19904
rect 44968 19864 44974 19876
rect 41230 19796 41236 19848
rect 41288 19796 41294 19848
rect 41690 19845 41696 19848
rect 41684 19836 41696 19845
rect 41651 19808 41696 19836
rect 41684 19799 41696 19808
rect 41690 19796 41696 19799
rect 41748 19796 41754 19848
rect 44637 19839 44695 19845
rect 44637 19805 44649 19839
rect 44683 19805 44695 19839
rect 44637 19799 44695 19805
rect 44821 19839 44879 19845
rect 44821 19805 44833 19839
rect 44867 19836 44879 19839
rect 45002 19836 45008 19848
rect 44867 19808 45008 19836
rect 44867 19805 44879 19808
rect 44821 19799 44879 19805
rect 44652 19768 44680 19799
rect 45002 19796 45008 19808
rect 45060 19796 45066 19848
rect 45388 19836 45416 19876
rect 46385 19873 46397 19907
rect 46431 19904 46443 19907
rect 47210 19904 47216 19916
rect 46431 19876 47216 19904
rect 46431 19873 46443 19876
rect 46385 19867 46443 19873
rect 47210 19864 47216 19876
rect 47268 19864 47274 19916
rect 49329 19907 49387 19913
rect 49329 19873 49341 19907
rect 49375 19904 49387 19907
rect 49804 19904 49832 20003
rect 49375 19876 49832 19904
rect 49375 19873 49387 19876
rect 49329 19867 49387 19873
rect 50154 19864 50160 19916
rect 50212 19864 50218 19916
rect 51460 19904 51488 20012
rect 52362 20000 52368 20052
rect 52420 20000 52426 20052
rect 52730 20000 52736 20052
rect 52788 20000 52794 20052
rect 55030 20000 55036 20052
rect 55088 20000 55094 20052
rect 57149 20043 57207 20049
rect 55140 20012 56723 20040
rect 51537 19975 51595 19981
rect 51537 19941 51549 19975
rect 51583 19972 51595 19975
rect 51994 19972 52000 19984
rect 51583 19944 52000 19972
rect 51583 19941 51595 19944
rect 51537 19935 51595 19941
rect 51994 19932 52000 19944
rect 52052 19932 52058 19984
rect 51810 19904 51816 19916
rect 51460 19876 51816 19904
rect 51810 19864 51816 19876
rect 51868 19904 51874 19916
rect 52748 19904 52776 20000
rect 55140 19972 55168 20012
rect 53852 19944 55168 19972
rect 52825 19907 52883 19913
rect 52825 19904 52837 19907
rect 51868 19876 52684 19904
rect 52748 19876 52837 19904
rect 51868 19864 51874 19876
rect 45554 19836 45560 19848
rect 45388 19808 45560 19836
rect 45554 19796 45560 19808
rect 45612 19796 45618 19848
rect 45738 19796 45744 19848
rect 45796 19836 45802 19848
rect 47029 19839 47087 19845
rect 47029 19836 47041 19839
rect 45796 19808 47041 19836
rect 45796 19796 45802 19808
rect 47029 19805 47041 19808
rect 47075 19805 47087 19839
rect 47029 19799 47087 19805
rect 49050 19796 49056 19848
rect 49108 19796 49114 19848
rect 51997 19839 52055 19845
rect 51997 19805 52009 19839
rect 52043 19836 52055 19839
rect 52086 19836 52092 19848
rect 52043 19808 52092 19836
rect 52043 19805 52055 19808
rect 51997 19799 52055 19805
rect 52086 19796 52092 19808
rect 52144 19796 52150 19848
rect 52656 19836 52684 19876
rect 52825 19873 52837 19876
rect 52871 19873 52883 19907
rect 52825 19867 52883 19873
rect 53852 19836 53880 19944
rect 53926 19864 53932 19916
rect 53984 19904 53990 19916
rect 54389 19907 54447 19913
rect 54389 19904 54401 19907
rect 53984 19876 54401 19904
rect 53984 19864 53990 19876
rect 54389 19873 54401 19876
rect 54435 19904 54447 19907
rect 55493 19907 55551 19913
rect 55493 19904 55505 19907
rect 54435 19876 55505 19904
rect 54435 19873 54447 19876
rect 54389 19867 54447 19873
rect 55493 19873 55505 19876
rect 55539 19873 55551 19907
rect 56695 19904 56723 20012
rect 57149 20009 57161 20043
rect 57195 20040 57207 20043
rect 58158 20040 58164 20052
rect 57195 20012 58164 20040
rect 57195 20009 57207 20012
rect 57149 20003 57207 20009
rect 58158 20000 58164 20012
rect 58216 20000 58222 20052
rect 57057 19975 57115 19981
rect 57057 19941 57069 19975
rect 57103 19972 57115 19975
rect 58434 19972 58440 19984
rect 57103 19944 58440 19972
rect 57103 19941 57115 19944
rect 57057 19935 57115 19941
rect 58434 19932 58440 19944
rect 58492 19932 58498 19984
rect 57793 19907 57851 19913
rect 57793 19904 57805 19907
rect 56695 19876 57805 19904
rect 55493 19867 55551 19873
rect 57793 19873 57805 19876
rect 57839 19904 57851 19907
rect 58161 19907 58219 19913
rect 58161 19904 58173 19907
rect 57839 19876 58173 19904
rect 57839 19873 57851 19876
rect 57793 19867 57851 19873
rect 58161 19873 58173 19876
rect 58207 19873 58219 19907
rect 58161 19867 58219 19873
rect 52656 19808 53880 19836
rect 54110 19796 54116 19848
rect 54168 19836 54174 19848
rect 55674 19836 55680 19848
rect 54168 19808 55680 19836
rect 54168 19796 54174 19808
rect 55674 19796 55680 19808
rect 55732 19796 55738 19848
rect 56962 19796 56968 19848
rect 57020 19836 57026 19848
rect 57517 19839 57575 19845
rect 57517 19836 57529 19839
rect 57020 19808 57529 19836
rect 57020 19796 57026 19808
rect 57517 19805 57529 19808
rect 57563 19805 57575 19839
rect 57517 19799 57575 19805
rect 45922 19768 45928 19780
rect 44652 19740 45928 19768
rect 45922 19728 45928 19740
rect 45980 19728 45986 19780
rect 47486 19777 47492 19780
rect 46140 19771 46198 19777
rect 46140 19737 46152 19771
rect 46186 19768 46198 19771
rect 46477 19771 46535 19777
rect 46477 19768 46489 19771
rect 46186 19740 46489 19768
rect 46186 19737 46198 19740
rect 46140 19731 46198 19737
rect 46477 19737 46489 19740
rect 46523 19737 46535 19771
rect 47480 19768 47492 19777
rect 47447 19740 47492 19768
rect 46477 19731 46535 19737
rect 47480 19731 47492 19740
rect 47486 19728 47492 19731
rect 47544 19728 47550 19780
rect 50246 19728 50252 19780
rect 50304 19768 50310 19780
rect 50402 19771 50460 19777
rect 50402 19768 50414 19771
rect 50304 19740 50414 19768
rect 50304 19728 50310 19740
rect 50402 19737 50414 19740
rect 50448 19737 50460 19771
rect 50402 19731 50460 19737
rect 53092 19771 53150 19777
rect 53092 19737 53104 19771
rect 53138 19768 53150 19771
rect 54386 19768 54392 19780
rect 53138 19740 54392 19768
rect 53138 19737 53150 19740
rect 53092 19731 53150 19737
rect 54386 19728 54392 19740
rect 54444 19728 54450 19780
rect 54665 19771 54723 19777
rect 54665 19737 54677 19771
rect 54711 19768 54723 19771
rect 55582 19768 55588 19780
rect 54711 19740 55588 19768
rect 54711 19737 54723 19740
rect 54665 19731 54723 19737
rect 55582 19728 55588 19740
rect 55640 19728 55646 19780
rect 55944 19771 56002 19777
rect 55944 19737 55956 19771
rect 55990 19768 56002 19771
rect 56502 19768 56508 19780
rect 55990 19740 56508 19768
rect 55990 19737 56002 19740
rect 55944 19731 56002 19737
rect 56502 19728 56508 19740
rect 56560 19728 56566 19780
rect 44450 19700 44456 19712
rect 41156 19672 44456 19700
rect 44450 19660 44456 19672
rect 44508 19660 44514 19712
rect 48314 19660 48320 19712
rect 48372 19700 48378 19712
rect 49145 19703 49203 19709
rect 49145 19700 49157 19703
rect 48372 19672 49157 19700
rect 48372 19660 48378 19672
rect 49145 19669 49157 19672
rect 49191 19700 49203 19703
rect 49786 19700 49792 19712
rect 49191 19672 49792 19700
rect 49191 19669 49203 19672
rect 49145 19663 49203 19669
rect 49786 19660 49792 19672
rect 49844 19660 49850 19712
rect 51258 19660 51264 19712
rect 51316 19700 51322 19712
rect 51905 19703 51963 19709
rect 51905 19700 51917 19703
rect 51316 19672 51917 19700
rect 51316 19660 51322 19672
rect 51905 19669 51917 19672
rect 51951 19700 51963 19703
rect 52270 19700 52276 19712
rect 51951 19672 52276 19700
rect 51951 19669 51963 19672
rect 51905 19663 51963 19669
rect 52270 19660 52276 19672
rect 52328 19660 52334 19712
rect 54202 19660 54208 19712
rect 54260 19660 54266 19712
rect 54478 19660 54484 19712
rect 54536 19700 54542 19712
rect 54573 19703 54631 19709
rect 54573 19700 54585 19703
rect 54536 19672 54585 19700
rect 54536 19660 54542 19672
rect 54573 19669 54585 19672
rect 54619 19700 54631 19703
rect 57609 19703 57667 19709
rect 57609 19700 57621 19703
rect 54619 19672 57621 19700
rect 54619 19669 54631 19672
rect 54573 19663 54631 19669
rect 57609 19669 57621 19672
rect 57655 19700 57667 19703
rect 58066 19700 58072 19712
rect 57655 19672 58072 19700
rect 57655 19669 57667 19672
rect 57609 19663 57667 19669
rect 58066 19660 58072 19672
rect 58124 19660 58130 19712
rect 1104 19610 59040 19632
rect 1104 19558 15394 19610
rect 15446 19558 15458 19610
rect 15510 19558 15522 19610
rect 15574 19558 15586 19610
rect 15638 19558 15650 19610
rect 15702 19558 29838 19610
rect 29890 19558 29902 19610
rect 29954 19558 29966 19610
rect 30018 19558 30030 19610
rect 30082 19558 30094 19610
rect 30146 19558 44282 19610
rect 44334 19558 44346 19610
rect 44398 19558 44410 19610
rect 44462 19558 44474 19610
rect 44526 19558 44538 19610
rect 44590 19558 58726 19610
rect 58778 19558 58790 19610
rect 58842 19558 58854 19610
rect 58906 19558 58918 19610
rect 58970 19558 58982 19610
rect 59034 19558 59040 19610
rect 1104 19536 59040 19558
rect 1949 19499 2007 19505
rect 1949 19465 1961 19499
rect 1995 19496 2007 19499
rect 2130 19496 2136 19508
rect 1995 19468 2136 19496
rect 1995 19465 2007 19468
rect 1949 19459 2007 19465
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 2866 19456 2872 19508
rect 2924 19456 2930 19508
rect 3418 19456 3424 19508
rect 3476 19456 3482 19508
rect 3789 19499 3847 19505
rect 3789 19465 3801 19499
rect 3835 19496 3847 19499
rect 4522 19496 4528 19508
rect 3835 19468 4528 19496
rect 3835 19465 3847 19468
rect 3789 19459 3847 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 6270 19456 6276 19508
rect 6328 19496 6334 19508
rect 6733 19499 6791 19505
rect 6733 19496 6745 19499
rect 6328 19468 6745 19496
rect 6328 19456 6334 19468
rect 6733 19465 6745 19468
rect 6779 19465 6791 19499
rect 6733 19459 6791 19465
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7558 19496 7564 19508
rect 7147 19468 7564 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 13909 19499 13967 19505
rect 13909 19496 13921 19499
rect 13412 19468 13921 19496
rect 13412 19456 13418 19468
rect 13909 19465 13921 19468
rect 13955 19465 13967 19499
rect 13909 19459 13967 19465
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 16666 19496 16672 19508
rect 16531 19468 16672 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 17310 19456 17316 19508
rect 17368 19456 17374 19508
rect 17681 19499 17739 19505
rect 17681 19465 17693 19499
rect 17727 19496 17739 19499
rect 18230 19496 18236 19508
rect 17727 19468 18236 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 18230 19456 18236 19468
rect 18288 19456 18294 19508
rect 19886 19456 19892 19508
rect 19944 19456 19950 19508
rect 19978 19456 19984 19508
rect 20036 19456 20042 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20990 19496 20996 19508
rect 20947 19468 20996 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21361 19499 21419 19505
rect 21361 19465 21373 19499
rect 21407 19496 21419 19499
rect 22370 19496 22376 19508
rect 21407 19468 22376 19496
rect 21407 19465 21419 19468
rect 21361 19459 21419 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 23072 19468 23213 19496
rect 23072 19456 23078 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 25501 19499 25559 19505
rect 25501 19465 25513 19499
rect 25547 19496 25559 19499
rect 25774 19496 25780 19508
rect 25547 19468 25780 19496
rect 25547 19465 25559 19468
rect 25501 19459 25559 19465
rect 25774 19456 25780 19468
rect 25832 19456 25838 19508
rect 26329 19499 26387 19505
rect 26329 19465 26341 19499
rect 26375 19496 26387 19499
rect 26694 19496 26700 19508
rect 26375 19468 26700 19496
rect 26375 19465 26387 19468
rect 26329 19459 26387 19465
rect 26694 19456 26700 19468
rect 26752 19456 26758 19508
rect 26789 19499 26847 19505
rect 26789 19465 26801 19499
rect 26835 19496 26847 19499
rect 27246 19496 27252 19508
rect 26835 19468 27252 19496
rect 26835 19465 26847 19468
rect 26789 19459 26847 19465
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 28629 19499 28687 19505
rect 28629 19465 28641 19499
rect 28675 19496 28687 19499
rect 28718 19496 28724 19508
rect 28675 19468 28724 19496
rect 28675 19465 28687 19468
rect 28629 19459 28687 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 30101 19499 30159 19505
rect 30101 19496 30113 19499
rect 29932 19468 30113 19496
rect 2884 19428 2912 19456
rect 3062 19431 3120 19437
rect 3062 19428 3074 19431
rect 2884 19400 3074 19428
rect 3062 19397 3074 19400
rect 3108 19397 3120 19431
rect 3062 19391 3120 19397
rect 3878 19388 3884 19440
rect 3936 19428 3942 19440
rect 12704 19431 12762 19437
rect 3936 19400 6684 19428
rect 3936 19388 3942 19400
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 3344 19168 3372 19323
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 6656 19369 6684 19400
rect 12704 19397 12716 19431
rect 12750 19428 12762 19431
rect 12802 19428 12808 19440
rect 12750 19400 12808 19428
rect 12750 19397 12762 19400
rect 12704 19391 12762 19397
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 19904 19428 19932 19456
rect 21174 19428 21180 19440
rect 15212 19400 18644 19428
rect 19904 19400 21180 19428
rect 15212 19372 15240 19400
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 4120 19332 4261 19360
rect 4120 19320 4126 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 9769 19363 9827 19369
rect 6687 19332 7604 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 7576 19304 7604 19332
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 9858 19360 9864 19372
rect 9815 19332 9864 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 12526 19360 12532 19372
rect 12483 19332 12532 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14461 19363 14519 19369
rect 14461 19360 14473 19363
rect 14148 19332 14473 19360
rect 14148 19320 14154 19332
rect 14461 19329 14473 19332
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15194 19360 15200 19372
rect 15151 19332 15200 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15372 19363 15430 19369
rect 15372 19329 15384 19363
rect 15418 19360 15430 19363
rect 15654 19360 15660 19372
rect 15418 19332 15660 19360
rect 15418 19329 15430 19332
rect 15372 19323 15430 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 18616 19369 18644 19400
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 23934 19428 23940 19440
rect 21784 19400 23940 19428
rect 21784 19388 21790 19400
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 15896 19332 17233 19360
rect 15896 19320 15902 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 18868 19363 18926 19369
rect 18868 19329 18880 19363
rect 18914 19360 18926 19363
rect 19242 19360 19248 19372
rect 18914 19332 19248 19360
rect 18914 19329 18926 19332
rect 18868 19323 18926 19329
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 21266 19360 21272 19372
rect 20772 19332 21272 19360
rect 20772 19320 20778 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21836 19369 21864 19400
rect 23934 19388 23940 19400
rect 23992 19428 23998 19440
rect 29764 19431 29822 19437
rect 23992 19400 27016 19428
rect 23992 19388 23998 19400
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 24136 19369 24164 19400
rect 26988 19372 27016 19400
rect 27080 19400 27568 19428
rect 24394 19369 24400 19372
rect 22077 19363 22135 19369
rect 22077 19360 22089 19363
rect 21968 19332 22089 19360
rect 21968 19320 21974 19332
rect 22077 19329 22089 19332
rect 22123 19329 22135 19363
rect 22077 19323 22135 19329
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 24388 19323 24400 19369
rect 24394 19320 24400 19323
rect 24452 19320 24458 19372
rect 25130 19320 25136 19372
rect 25188 19360 25194 19372
rect 26326 19360 26332 19372
rect 25188 19332 26332 19360
rect 25188 19320 25194 19332
rect 26326 19320 26332 19332
rect 26384 19360 26390 19372
rect 26421 19363 26479 19369
rect 26421 19360 26433 19363
rect 26384 19332 26433 19360
rect 26384 19320 26390 19332
rect 26421 19329 26433 19332
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 3973 19295 4031 19301
rect 3973 19261 3985 19295
rect 4019 19261 4031 19295
rect 3973 19255 4031 19261
rect 2038 19116 2044 19168
rect 2096 19156 2102 19168
rect 3326 19156 3332 19168
rect 2096 19128 3332 19156
rect 2096 19116 2102 19128
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 3988 19156 4016 19255
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4212 19264 4813 19292
rect 4212 19252 4218 19264
rect 4801 19261 4813 19264
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 7374 19292 7380 19304
rect 6512 19264 7380 19292
rect 6512 19252 6518 19264
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7558 19252 7564 19304
rect 7616 19252 7622 19304
rect 7834 19252 7840 19304
rect 7892 19252 7898 19304
rect 9585 19295 9643 19301
rect 9585 19261 9597 19295
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 8481 19227 8539 19233
rect 8481 19224 8493 19227
rect 7668 19196 8493 19224
rect 7668 19168 7696 19196
rect 8481 19193 8493 19196
rect 8527 19193 8539 19227
rect 9600 19224 9628 19255
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 10594 19292 10600 19304
rect 9784 19264 10600 19292
rect 9784 19224 9812 19264
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19261 10839 19295
rect 10781 19255 10839 19261
rect 9600 19196 9812 19224
rect 10137 19227 10195 19233
rect 8481 19187 8539 19193
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 10796 19224 10824 19255
rect 17034 19252 17040 19304
rect 17092 19252 17098 19304
rect 21453 19295 21511 19301
rect 21453 19292 21465 19295
rect 20916 19264 21465 19292
rect 10183 19196 10824 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 20916 19168 20944 19264
rect 21453 19261 21465 19264
rect 21499 19261 21511 19295
rect 21453 19255 21511 19261
rect 26237 19295 26295 19301
rect 26237 19261 26249 19295
rect 26283 19292 26295 19295
rect 26436 19292 26464 19323
rect 26970 19320 26976 19372
rect 27028 19320 27034 19372
rect 27080 19292 27108 19400
rect 27540 19372 27568 19400
rect 29764 19397 29776 19431
rect 29810 19428 29822 19431
rect 29932 19428 29960 19468
rect 30101 19465 30113 19468
rect 30147 19465 30159 19499
rect 30101 19459 30159 19465
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19496 30527 19499
rect 31018 19496 31024 19508
rect 30515 19468 31024 19496
rect 30515 19465 30527 19468
rect 30469 19459 30527 19465
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 32674 19456 32680 19508
rect 32732 19496 32738 19508
rect 35437 19499 35495 19505
rect 35437 19496 35449 19499
rect 32732 19468 35449 19496
rect 32732 19456 32738 19468
rect 35437 19465 35449 19468
rect 35483 19465 35495 19499
rect 35437 19459 35495 19465
rect 35526 19456 35532 19508
rect 35584 19456 35590 19508
rect 35802 19456 35808 19508
rect 35860 19496 35866 19508
rect 37277 19499 37335 19505
rect 35860 19468 36308 19496
rect 35860 19456 35866 19468
rect 31110 19428 31116 19440
rect 29810 19400 29960 19428
rect 30024 19400 31116 19428
rect 29810 19397 29822 19400
rect 29764 19391 29822 19397
rect 27246 19369 27252 19372
rect 27240 19323 27252 19369
rect 27246 19320 27252 19323
rect 27304 19320 27310 19372
rect 27522 19320 27528 19372
rect 27580 19320 27586 19372
rect 30024 19369 30052 19400
rect 31110 19388 31116 19400
rect 31168 19428 31174 19440
rect 33870 19428 33876 19440
rect 31168 19400 33876 19428
rect 31168 19388 31174 19400
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19329 30067 19363
rect 30009 19323 30067 19329
rect 30558 19320 30564 19372
rect 30616 19320 30622 19372
rect 32140 19369 32168 19400
rect 33870 19388 33876 19400
rect 33928 19428 33934 19440
rect 36280 19428 36308 19468
rect 37277 19465 37289 19499
rect 37323 19496 37335 19499
rect 37550 19496 37556 19508
rect 37323 19468 37556 19496
rect 37323 19465 37335 19468
rect 37277 19459 37335 19465
rect 37550 19456 37556 19468
rect 37608 19456 37614 19508
rect 37645 19499 37703 19505
rect 37645 19465 37657 19499
rect 37691 19496 37703 19499
rect 38378 19496 38384 19508
rect 37691 19468 38384 19496
rect 37691 19465 37703 19468
rect 37645 19459 37703 19465
rect 38378 19456 38384 19468
rect 38436 19456 38442 19508
rect 39114 19456 39120 19508
rect 39172 19456 39178 19508
rect 40129 19499 40187 19505
rect 40129 19465 40141 19499
rect 40175 19496 40187 19499
rect 41230 19496 41236 19508
rect 40175 19468 41236 19496
rect 40175 19465 40187 19468
rect 40129 19459 40187 19465
rect 41230 19456 41236 19468
rect 41288 19456 41294 19508
rect 43809 19499 43867 19505
rect 43809 19465 43821 19499
rect 43855 19496 43867 19499
rect 44174 19496 44180 19508
rect 43855 19468 44180 19496
rect 43855 19465 43867 19468
rect 43809 19459 43867 19465
rect 44174 19456 44180 19468
rect 44232 19456 44238 19508
rect 45373 19499 45431 19505
rect 45373 19465 45385 19499
rect 45419 19496 45431 19499
rect 45922 19496 45928 19508
rect 45419 19468 45928 19496
rect 45419 19465 45431 19468
rect 45373 19459 45431 19465
rect 45922 19456 45928 19468
rect 45980 19456 45986 19508
rect 48961 19499 49019 19505
rect 48961 19465 48973 19499
rect 49007 19496 49019 19499
rect 49694 19496 49700 19508
rect 49007 19468 49700 19496
rect 49007 19465 49019 19468
rect 48961 19459 49019 19465
rect 49694 19456 49700 19468
rect 49752 19456 49758 19508
rect 50157 19499 50215 19505
rect 50157 19465 50169 19499
rect 50203 19496 50215 19499
rect 50246 19496 50252 19508
rect 50203 19468 50252 19496
rect 50203 19465 50215 19468
rect 50157 19459 50215 19465
rect 50246 19456 50252 19468
rect 50304 19456 50310 19508
rect 50525 19499 50583 19505
rect 50525 19465 50537 19499
rect 50571 19496 50583 19499
rect 51350 19496 51356 19508
rect 50571 19468 51356 19496
rect 50571 19465 50583 19468
rect 50525 19459 50583 19465
rect 51350 19456 51356 19468
rect 51408 19456 51414 19508
rect 51537 19499 51595 19505
rect 51537 19496 51549 19499
rect 51460 19468 51549 19496
rect 37826 19428 37832 19440
rect 33928 19400 36216 19428
rect 36280 19400 37832 19428
rect 33928 19388 33934 19400
rect 31941 19363 31999 19369
rect 31941 19329 31953 19363
rect 31987 19360 31999 19363
rect 32125 19363 32183 19369
rect 31987 19332 32076 19360
rect 31987 19329 31999 19332
rect 31941 19323 31999 19329
rect 26283 19264 26372 19292
rect 26436 19264 27108 19292
rect 26283 19261 26295 19264
rect 26237 19255 26295 19261
rect 5258 19156 5264 19168
rect 3988 19128 5264 19156
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5350 19116 5356 19168
rect 5408 19156 5414 19168
rect 5813 19159 5871 19165
rect 5813 19156 5825 19159
rect 5408 19128 5825 19156
rect 5408 19116 5414 19128
rect 5813 19125 5825 19128
rect 5859 19156 5871 19159
rect 7098 19156 7104 19168
rect 5859 19128 7104 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7190 19116 7196 19168
rect 7248 19116 7254 19168
rect 7650 19116 7656 19168
rect 7708 19116 7714 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 7984 19128 8217 19156
rect 7984 19116 7990 19128
rect 8205 19125 8217 19128
rect 8251 19156 8263 19159
rect 9398 19156 9404 19168
rect 8251 19128 9404 19156
rect 8251 19125 8263 19128
rect 8205 19119 8263 19125
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 10226 19116 10232 19168
rect 10284 19116 10290 19168
rect 13817 19159 13875 19165
rect 13817 19125 13829 19159
rect 13863 19156 13875 19159
rect 14550 19156 14556 19168
rect 13863 19128 14556 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18598 19156 18604 19168
rect 18279 19128 18604 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 20349 19159 20407 19165
rect 20349 19125 20361 19159
rect 20395 19156 20407 19159
rect 20438 19156 20444 19168
rect 20395 19128 20444 19156
rect 20395 19125 20407 19128
rect 20349 19119 20407 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20809 19159 20867 19165
rect 20809 19125 20821 19159
rect 20855 19156 20867 19159
rect 20898 19156 20904 19168
rect 20855 19128 20904 19156
rect 20855 19125 20867 19128
rect 20809 19119 20867 19125
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 23382 19116 23388 19168
rect 23440 19156 23446 19168
rect 23937 19159 23995 19165
rect 23937 19156 23949 19159
rect 23440 19128 23949 19156
rect 23440 19116 23446 19128
rect 23937 19125 23949 19128
rect 23983 19156 23995 19159
rect 25406 19156 25412 19168
rect 23983 19128 25412 19156
rect 23983 19125 23995 19128
rect 23937 19119 23995 19125
rect 25406 19116 25412 19128
rect 25464 19116 25470 19168
rect 25961 19159 26019 19165
rect 25961 19125 25973 19159
rect 26007 19156 26019 19159
rect 26050 19156 26056 19168
rect 26007 19128 26056 19156
rect 26007 19125 26019 19128
rect 25961 19119 26019 19125
rect 26050 19116 26056 19128
rect 26108 19156 26114 19168
rect 26344 19156 26372 19264
rect 30098 19252 30104 19304
rect 30156 19292 30162 19304
rect 30653 19295 30711 19301
rect 30653 19292 30665 19295
rect 30156 19264 30665 19292
rect 30156 19252 30162 19264
rect 30653 19261 30665 19264
rect 30699 19261 30711 19295
rect 30653 19255 30711 19261
rect 31386 19252 31392 19304
rect 31444 19252 31450 19304
rect 32048 19292 32076 19332
rect 32125 19329 32137 19363
rect 32171 19329 32183 19363
rect 32381 19363 32439 19369
rect 32381 19360 32393 19363
rect 32125 19323 32183 19329
rect 32232 19332 32393 19360
rect 32232 19292 32260 19332
rect 32381 19329 32393 19332
rect 32427 19329 32439 19363
rect 34146 19360 34152 19372
rect 32381 19323 32439 19329
rect 33520 19332 34152 19360
rect 32048 19264 32260 19292
rect 33520 19233 33548 19332
rect 34146 19320 34152 19332
rect 34204 19320 34210 19372
rect 34992 19369 35020 19400
rect 36188 19372 36216 19400
rect 37826 19388 37832 19400
rect 37884 19388 37890 19440
rect 39132 19428 39160 19456
rect 38764 19400 39160 19428
rect 34721 19363 34779 19369
rect 34721 19329 34733 19363
rect 34767 19360 34779 19363
rect 34977 19363 35035 19369
rect 34767 19332 34928 19360
rect 34767 19329 34779 19332
rect 34721 19323 34779 19329
rect 34900 19292 34928 19332
rect 34977 19329 34989 19363
rect 35023 19329 35035 19363
rect 35897 19363 35955 19369
rect 35897 19360 35909 19363
rect 34977 19323 35035 19329
rect 35084 19332 35909 19360
rect 35084 19292 35112 19332
rect 35897 19329 35909 19332
rect 35943 19329 35955 19363
rect 35897 19323 35955 19329
rect 36170 19320 36176 19372
rect 36228 19320 36234 19372
rect 37458 19360 37464 19372
rect 36280 19332 37464 19360
rect 34900 19264 35112 19292
rect 35618 19252 35624 19304
rect 35676 19252 35682 19304
rect 35710 19252 35716 19304
rect 35768 19252 35774 19304
rect 36078 19252 36084 19304
rect 36136 19292 36142 19304
rect 36280 19292 36308 19332
rect 37458 19320 37464 19332
rect 37516 19320 37522 19372
rect 37737 19363 37795 19369
rect 37737 19329 37749 19363
rect 37783 19360 37795 19363
rect 38470 19360 38476 19372
rect 37783 19332 38476 19360
rect 37783 19329 37795 19332
rect 37737 19323 37795 19329
rect 38470 19320 38476 19332
rect 38528 19320 38534 19372
rect 38764 19369 38792 19400
rect 39574 19388 39580 19440
rect 39632 19388 39638 19440
rect 40494 19388 40500 19440
rect 40552 19388 40558 19440
rect 40589 19431 40647 19437
rect 40589 19397 40601 19431
rect 40635 19428 40647 19431
rect 41046 19428 41052 19440
rect 40635 19400 41052 19428
rect 40635 19397 40647 19400
rect 40589 19391 40647 19397
rect 41046 19388 41052 19400
rect 41104 19388 41110 19440
rect 42444 19400 45876 19428
rect 38749 19363 38807 19369
rect 38749 19329 38761 19363
rect 38795 19329 38807 19363
rect 38749 19323 38807 19329
rect 39016 19363 39074 19369
rect 39016 19329 39028 19363
rect 39062 19360 39074 19363
rect 39592 19360 39620 19388
rect 40512 19360 40540 19388
rect 39062 19332 39620 19360
rect 40236 19332 40540 19360
rect 40681 19363 40739 19369
rect 39062 19329 39074 19332
rect 39016 19323 39074 19329
rect 36136 19264 36308 19292
rect 36136 19252 36142 19264
rect 36446 19252 36452 19304
rect 36504 19252 36510 19304
rect 37829 19295 37887 19301
rect 37829 19292 37841 19295
rect 37108 19264 37841 19292
rect 33505 19227 33563 19233
rect 27908 19196 28488 19224
rect 27908 19156 27936 19196
rect 26108 19128 27936 19156
rect 26108 19116 26114 19128
rect 28350 19116 28356 19168
rect 28408 19116 28414 19168
rect 28460 19156 28488 19196
rect 33505 19193 33517 19227
rect 33551 19193 33563 19227
rect 33505 19187 33563 19193
rect 35526 19184 35532 19236
rect 35584 19224 35590 19236
rect 35728 19224 35756 19252
rect 37108 19233 37136 19264
rect 37829 19261 37841 19264
rect 37875 19292 37887 19295
rect 37875 19264 38424 19292
rect 37875 19261 37887 19264
rect 37829 19255 37887 19261
rect 37093 19227 37151 19233
rect 37093 19224 37105 19227
rect 35584 19196 37105 19224
rect 35584 19184 35590 19196
rect 37093 19193 37105 19196
rect 37139 19193 37151 19227
rect 37093 19187 37151 19193
rect 30650 19156 30656 19168
rect 28460 19128 30656 19156
rect 30650 19116 30656 19128
rect 30708 19116 30714 19168
rect 33594 19116 33600 19168
rect 33652 19116 33658 19168
rect 35066 19116 35072 19168
rect 35124 19116 35130 19168
rect 38286 19116 38292 19168
rect 38344 19116 38350 19168
rect 38396 19156 38424 19264
rect 40236 19233 40264 19332
rect 40681 19329 40693 19363
rect 40727 19360 40739 19363
rect 40862 19360 40868 19372
rect 40727 19332 40868 19360
rect 40727 19329 40739 19332
rect 40681 19323 40739 19329
rect 40862 19320 40868 19332
rect 40920 19320 40926 19372
rect 42444 19304 42472 19400
rect 42696 19363 42754 19369
rect 42696 19329 42708 19363
rect 42742 19360 42754 19363
rect 43070 19360 43076 19372
rect 42742 19332 43076 19360
rect 42742 19329 42754 19332
rect 42696 19323 42754 19329
rect 43070 19320 43076 19332
rect 43128 19320 43134 19372
rect 43714 19320 43720 19372
rect 43772 19360 43778 19372
rect 44269 19363 44327 19369
rect 44269 19360 44281 19363
rect 43772 19332 44281 19360
rect 43772 19320 43778 19332
rect 44269 19329 44281 19332
rect 44315 19360 44327 19363
rect 45281 19363 45339 19369
rect 45281 19360 45293 19363
rect 44315 19332 45293 19360
rect 44315 19329 44327 19332
rect 44269 19323 44327 19329
rect 45281 19329 45293 19332
rect 45327 19360 45339 19363
rect 45462 19360 45468 19372
rect 45327 19332 45468 19360
rect 45327 19329 45339 19332
rect 45281 19323 45339 19329
rect 45462 19320 45468 19332
rect 45520 19320 45526 19372
rect 45738 19320 45744 19372
rect 45796 19320 45802 19372
rect 45848 19369 45876 19400
rect 47688 19400 50200 19428
rect 46106 19369 46112 19372
rect 45833 19363 45891 19369
rect 45833 19329 45845 19363
rect 45879 19329 45891 19363
rect 45833 19323 45891 19329
rect 46100 19323 46112 19369
rect 46106 19320 46112 19323
rect 46164 19320 46170 19372
rect 47210 19320 47216 19372
rect 47268 19360 47274 19372
rect 47570 19363 47628 19369
rect 47570 19360 47582 19363
rect 47268 19332 47582 19360
rect 47268 19320 47274 19332
rect 47570 19329 47582 19332
rect 47616 19360 47628 19363
rect 47688 19360 47716 19400
rect 50172 19372 50200 19400
rect 51258 19388 51264 19440
rect 51316 19428 51322 19440
rect 51460 19428 51488 19468
rect 51537 19465 51549 19468
rect 51583 19496 51595 19499
rect 51810 19496 51816 19508
rect 51583 19468 51816 19496
rect 51583 19465 51595 19468
rect 51537 19459 51595 19465
rect 51810 19456 51816 19468
rect 51868 19456 51874 19508
rect 52730 19456 52736 19508
rect 52788 19456 52794 19508
rect 54294 19456 54300 19508
rect 54352 19456 54358 19508
rect 54386 19456 54392 19508
rect 54444 19456 54450 19508
rect 55582 19456 55588 19508
rect 55640 19496 55646 19508
rect 55769 19499 55827 19505
rect 55769 19496 55781 19499
rect 55640 19468 55781 19496
rect 55640 19456 55646 19468
rect 55769 19465 55781 19468
rect 55815 19465 55827 19499
rect 55769 19459 55827 19465
rect 56686 19456 56692 19508
rect 56744 19456 56750 19508
rect 56962 19456 56968 19508
rect 57020 19496 57026 19508
rect 57885 19499 57943 19505
rect 57885 19496 57897 19499
rect 57020 19468 57897 19496
rect 57020 19456 57026 19468
rect 57885 19465 57897 19468
rect 57931 19465 57943 19499
rect 57885 19459 57943 19465
rect 51316 19400 51488 19428
rect 52748 19428 52776 19456
rect 54110 19428 54116 19440
rect 52748 19400 54116 19428
rect 51316 19388 51322 19400
rect 47854 19369 47860 19372
rect 47848 19360 47860 19369
rect 47616 19332 47716 19360
rect 47815 19332 47860 19360
rect 47616 19329 47628 19332
rect 47570 19323 47628 19329
rect 47848 19323 47860 19332
rect 47854 19320 47860 19323
rect 47912 19320 47918 19372
rect 50154 19320 50160 19372
rect 50212 19320 50218 19372
rect 50617 19363 50675 19369
rect 50617 19329 50629 19363
rect 50663 19360 50675 19363
rect 50982 19360 50988 19372
rect 50663 19332 50988 19360
rect 50663 19329 50675 19332
rect 50617 19323 50675 19329
rect 50982 19320 50988 19332
rect 51040 19320 51046 19372
rect 52748 19360 52776 19400
rect 54110 19388 54116 19400
rect 54168 19388 54174 19440
rect 56496 19431 56554 19437
rect 56496 19397 56508 19431
rect 56542 19428 56554 19431
rect 56704 19428 56732 19456
rect 56542 19400 56732 19428
rect 56542 19397 56554 19400
rect 56496 19391 56554 19397
rect 53190 19369 53196 19372
rect 52917 19363 52975 19369
rect 52917 19360 52929 19363
rect 52748 19332 52929 19360
rect 52917 19329 52929 19332
rect 52963 19329 52975 19363
rect 53184 19360 53196 19369
rect 53151 19332 53196 19360
rect 52917 19323 52975 19329
rect 53184 19323 53196 19332
rect 53190 19320 53196 19323
rect 53248 19320 53254 19372
rect 54202 19320 54208 19372
rect 54260 19320 54266 19372
rect 55030 19320 55036 19372
rect 55088 19320 55094 19372
rect 55674 19320 55680 19372
rect 55732 19360 55738 19372
rect 56226 19360 56232 19372
rect 55732 19332 56232 19360
rect 55732 19320 55738 19332
rect 56226 19320 56232 19332
rect 56284 19320 56290 19372
rect 58434 19320 58440 19372
rect 58492 19320 58498 19372
rect 40770 19252 40776 19304
rect 40828 19252 40834 19304
rect 42426 19252 42432 19304
rect 42484 19252 42490 19304
rect 43898 19252 43904 19304
rect 43956 19292 43962 19304
rect 43993 19295 44051 19301
rect 43993 19292 44005 19295
rect 43956 19264 44005 19292
rect 43956 19252 43962 19264
rect 43993 19261 44005 19264
rect 44039 19261 44051 19295
rect 43993 19255 44051 19261
rect 44177 19295 44235 19301
rect 44177 19261 44189 19295
rect 44223 19292 44235 19295
rect 45002 19292 45008 19304
rect 44223 19264 45008 19292
rect 44223 19261 44235 19264
rect 44177 19255 44235 19261
rect 40221 19227 40279 19233
rect 40221 19193 40233 19227
rect 40267 19193 40279 19227
rect 44008 19224 44036 19255
rect 45002 19252 45008 19264
rect 45060 19252 45066 19304
rect 45094 19252 45100 19304
rect 45152 19252 45158 19304
rect 45756 19233 45784 19320
rect 50709 19295 50767 19301
rect 50709 19292 50721 19295
rect 49988 19264 50721 19292
rect 45741 19227 45799 19233
rect 44008 19196 45692 19224
rect 40221 19187 40279 19193
rect 41414 19156 41420 19168
rect 38396 19128 41420 19156
rect 41414 19116 41420 19128
rect 41472 19156 41478 19168
rect 41782 19156 41788 19168
rect 41472 19128 41788 19156
rect 41472 19116 41478 19128
rect 41782 19116 41788 19128
rect 41840 19116 41846 19168
rect 44634 19116 44640 19168
rect 44692 19116 44698 19168
rect 45664 19156 45692 19196
rect 45741 19193 45753 19227
rect 45787 19193 45799 19227
rect 47394 19224 47400 19236
rect 45741 19187 45799 19193
rect 47136 19196 47400 19224
rect 47136 19156 47164 19196
rect 47394 19184 47400 19196
rect 47452 19184 47458 19236
rect 45664 19128 47164 19156
rect 47210 19116 47216 19168
rect 47268 19116 47274 19168
rect 47302 19116 47308 19168
rect 47360 19156 47366 19168
rect 49988 19165 50016 19264
rect 50709 19261 50721 19264
rect 50755 19261 50767 19295
rect 54220 19292 54248 19320
rect 55125 19295 55183 19301
rect 55125 19292 55137 19295
rect 54220 19264 55137 19292
rect 50709 19255 50767 19261
rect 55125 19261 55137 19264
rect 55171 19261 55183 19295
rect 55125 19255 55183 19261
rect 49973 19159 50031 19165
rect 49973 19156 49985 19159
rect 47360 19128 49985 19156
rect 47360 19116 47366 19128
rect 49973 19125 49985 19128
rect 50019 19125 50031 19159
rect 49973 19119 50031 19125
rect 57606 19116 57612 19168
rect 57664 19116 57670 19168
rect 1104 19066 58880 19088
rect 1104 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 22616 19066
rect 22668 19014 22680 19066
rect 22732 19014 22744 19066
rect 22796 19014 22808 19066
rect 22860 19014 22872 19066
rect 22924 19014 37060 19066
rect 37112 19014 37124 19066
rect 37176 19014 37188 19066
rect 37240 19014 37252 19066
rect 37304 19014 37316 19066
rect 37368 19014 51504 19066
rect 51556 19014 51568 19066
rect 51620 19014 51632 19066
rect 51684 19014 51696 19066
rect 51748 19014 51760 19066
rect 51812 19014 58880 19066
rect 1104 18992 58880 19014
rect 2133 18955 2191 18961
rect 2133 18921 2145 18955
rect 2179 18952 2191 18955
rect 2222 18952 2228 18964
rect 2179 18924 2228 18952
rect 2179 18921 2191 18924
rect 2133 18915 2191 18921
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 5534 18952 5540 18964
rect 3384 18924 5540 18952
rect 3384 18912 3390 18924
rect 5534 18912 5540 18924
rect 5592 18952 5598 18964
rect 5592 18924 5764 18952
rect 5592 18912 5598 18924
rect 3605 18887 3663 18893
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 4154 18884 4160 18896
rect 3651 18856 4160 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 4154 18844 4160 18856
rect 4212 18844 4218 18896
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18785 1639 18819
rect 3789 18819 3847 18825
rect 1581 18779 1639 18785
rect 1780 18788 2351 18816
rect 1596 18612 1624 18779
rect 1780 18757 1808 18788
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 2225 18751 2283 18757
rect 2225 18748 2237 18751
rect 2096 18720 2237 18748
rect 2096 18708 2102 18720
rect 2225 18717 2237 18720
rect 2271 18717 2283 18751
rect 2323 18748 2351 18788
rect 3789 18785 3801 18819
rect 3835 18816 3847 18819
rect 4062 18816 4068 18828
rect 3835 18788 4068 18816
rect 3835 18785 3847 18788
rect 3789 18779 3847 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4430 18776 4436 18828
rect 4488 18776 4494 18828
rect 4522 18776 4528 18828
rect 4580 18816 4586 18828
rect 4826 18819 4884 18825
rect 4826 18816 4838 18819
rect 4580 18788 4838 18816
rect 4580 18776 4586 18788
rect 4826 18785 4838 18788
rect 4872 18785 4884 18819
rect 4826 18779 4884 18785
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5350 18816 5356 18828
rect 5031 18788 5356 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 5736 18825 5764 18924
rect 6914 18912 6920 18964
rect 6972 18952 6978 18964
rect 7101 18955 7159 18961
rect 7101 18952 7113 18955
rect 6972 18924 7113 18952
rect 6972 18912 6978 18924
rect 7101 18921 7113 18924
rect 7147 18921 7159 18955
rect 7101 18915 7159 18921
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 7892 18924 7941 18952
rect 7892 18912 7898 18924
rect 7929 18921 7941 18924
rect 7975 18921 7987 18955
rect 7929 18915 7987 18921
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 10134 18952 10140 18964
rect 9732 18924 10140 18952
rect 9732 18912 9738 18924
rect 10134 18912 10140 18924
rect 10192 18952 10198 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 10192 18924 10517 18952
rect 10192 18912 10198 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 15654 18912 15660 18964
rect 15712 18952 15718 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15712 18924 16037 18952
rect 15712 18912 15718 18924
rect 16025 18921 16037 18924
rect 16071 18921 16083 18955
rect 16025 18915 16083 18921
rect 17034 18912 17040 18964
rect 17092 18912 17098 18964
rect 19242 18912 19248 18964
rect 19300 18912 19306 18964
rect 21082 18912 21088 18964
rect 21140 18912 21146 18964
rect 24394 18912 24400 18964
rect 24452 18952 24458 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 24452 18924 24593 18952
rect 24452 18912 24458 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 26970 18912 26976 18964
rect 27028 18952 27034 18964
rect 27065 18955 27123 18961
rect 27065 18952 27077 18955
rect 27028 18924 27077 18952
rect 27028 18912 27034 18924
rect 27065 18921 27077 18924
rect 27111 18921 27123 18955
rect 27065 18915 27123 18921
rect 29086 18912 29092 18964
rect 29144 18952 29150 18964
rect 30009 18955 30067 18961
rect 30009 18952 30021 18955
rect 29144 18924 30021 18952
rect 29144 18912 29150 18924
rect 30009 18921 30021 18924
rect 30055 18952 30067 18955
rect 30098 18952 30104 18964
rect 30055 18924 30104 18952
rect 30055 18921 30067 18924
rect 30009 18915 30067 18921
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 31386 18912 31392 18964
rect 31444 18952 31450 18964
rect 32033 18955 32091 18961
rect 32033 18952 32045 18955
rect 31444 18924 32045 18952
rect 31444 18912 31450 18924
rect 32033 18921 32045 18924
rect 32079 18921 32091 18955
rect 32033 18915 32091 18921
rect 34241 18955 34299 18961
rect 34241 18921 34253 18955
rect 34287 18952 34299 18955
rect 36446 18952 36452 18964
rect 34287 18924 36452 18952
rect 34287 18921 34299 18924
rect 34241 18915 34299 18921
rect 36446 18912 36452 18924
rect 36504 18912 36510 18964
rect 38654 18912 38660 18964
rect 38712 18952 38718 18964
rect 39117 18955 39175 18961
rect 39117 18952 39129 18955
rect 38712 18924 39129 18952
rect 38712 18912 38718 18924
rect 39117 18921 39129 18924
rect 39163 18921 39175 18955
rect 39117 18915 39175 18921
rect 40129 18955 40187 18961
rect 40129 18921 40141 18955
rect 40175 18952 40187 18955
rect 40770 18952 40776 18964
rect 40175 18924 40776 18952
rect 40175 18921 40187 18924
rect 40129 18915 40187 18921
rect 40770 18912 40776 18924
rect 40828 18912 40834 18964
rect 45002 18912 45008 18964
rect 45060 18912 45066 18964
rect 46017 18955 46075 18961
rect 46017 18921 46029 18955
rect 46063 18952 46075 18955
rect 46106 18952 46112 18964
rect 46063 18924 46112 18952
rect 46063 18921 46075 18924
rect 46017 18915 46075 18921
rect 46106 18912 46112 18924
rect 46164 18912 46170 18964
rect 54110 18912 54116 18964
rect 54168 18912 54174 18964
rect 56502 18912 56508 18964
rect 56560 18952 56566 18964
rect 57333 18955 57391 18961
rect 57333 18952 57345 18955
rect 56560 18924 57345 18952
rect 56560 18912 56566 18924
rect 57333 18921 57345 18924
rect 57379 18921 57391 18955
rect 57333 18915 57391 18921
rect 10413 18887 10471 18893
rect 10413 18853 10425 18887
rect 10459 18853 10471 18887
rect 21100 18884 21128 18912
rect 29454 18884 29460 18896
rect 21100 18856 21956 18884
rect 10413 18847 10471 18853
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18785 5779 18819
rect 5721 18779 5779 18785
rect 7377 18819 7435 18825
rect 7377 18785 7389 18819
rect 7423 18816 7435 18819
rect 7650 18816 7656 18828
rect 7423 18788 7656 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 10428 18816 10456 18847
rect 11057 18819 11115 18825
rect 11057 18816 11069 18819
rect 10428 18788 11069 18816
rect 11057 18785 11069 18788
rect 11103 18785 11115 18819
rect 11057 18779 11115 18785
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15933 18819 15991 18825
rect 15933 18816 15945 18819
rect 15344 18788 15945 18816
rect 15344 18776 15350 18788
rect 15933 18785 15945 18788
rect 15979 18816 15991 18819
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 15979 18788 16589 18816
rect 15979 18785 15991 18788
rect 15933 18779 15991 18785
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 19518 18776 19524 18828
rect 19576 18816 19582 18828
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19576 18788 19809 18816
rect 19576 18776 19582 18788
rect 19797 18785 19809 18788
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 2958 18748 2964 18760
rect 2323 18720 2964 18748
rect 2225 18711 2283 18717
rect 2958 18708 2964 18720
rect 3016 18748 3022 18760
rect 3016 18720 3924 18748
rect 3016 18708 3022 18720
rect 1673 18683 1731 18689
rect 1673 18649 1685 18683
rect 1719 18680 1731 18683
rect 2492 18683 2550 18689
rect 1719 18652 2452 18680
rect 1719 18649 1731 18652
rect 1673 18643 1731 18649
rect 1854 18612 1860 18624
rect 1596 18584 1860 18612
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 2424 18612 2452 18652
rect 2492 18649 2504 18683
rect 2538 18680 2550 18683
rect 3786 18680 3792 18692
rect 2538 18652 3792 18680
rect 2538 18649 2550 18652
rect 2492 18643 2550 18649
rect 3786 18640 3792 18652
rect 3844 18640 3850 18692
rect 3694 18612 3700 18624
rect 2424 18584 3700 18612
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 3896 18612 3924 18720
rect 3970 18708 3976 18760
rect 4028 18708 4034 18760
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 5988 18751 6046 18757
rect 5988 18717 6000 18751
rect 6034 18748 6046 18751
rect 7006 18748 7012 18760
rect 6034 18720 7012 18748
rect 6034 18717 6046 18720
rect 5988 18711 6046 18717
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7558 18708 7564 18760
rect 7616 18708 7622 18760
rect 8018 18708 8024 18760
rect 8076 18708 8082 18760
rect 9030 18708 9036 18760
rect 9088 18708 9094 18760
rect 9300 18751 9358 18757
rect 9300 18717 9312 18751
rect 9346 18748 9358 18751
rect 10226 18748 10232 18760
rect 9346 18720 10232 18748
rect 9346 18717 9358 18720
rect 9300 18711 9358 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18748 16451 18751
rect 17402 18748 17408 18760
rect 16439 18720 17408 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 21928 18748 21956 18856
rect 28000 18856 29460 18884
rect 22278 18776 22284 18828
rect 22336 18776 22342 18828
rect 22373 18819 22431 18825
rect 22373 18785 22385 18819
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 21928 18720 22201 18748
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 22379 18748 22407 18779
rect 24946 18776 24952 18828
rect 25004 18816 25010 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 25004 18788 25145 18816
rect 25004 18776 25010 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 27154 18776 27160 18828
rect 27212 18816 27218 18828
rect 28000 18825 28028 18856
rect 29454 18844 29460 18856
rect 29512 18844 29518 18896
rect 36078 18884 36084 18896
rect 32692 18856 36084 18884
rect 27985 18819 28043 18825
rect 27985 18816 27997 18819
rect 27212 18788 27997 18816
rect 27212 18776 27218 18788
rect 27985 18785 27997 18788
rect 28031 18785 28043 18819
rect 27985 18779 28043 18785
rect 28350 18776 28356 18828
rect 28408 18816 28414 18828
rect 28813 18819 28871 18825
rect 28813 18816 28825 18819
rect 28408 18788 28825 18816
rect 28408 18776 28414 18788
rect 28813 18785 28825 18788
rect 28859 18785 28871 18819
rect 28813 18779 28871 18785
rect 31938 18776 31944 18828
rect 31996 18816 32002 18828
rect 32692 18825 32720 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 37645 18887 37703 18893
rect 37645 18853 37657 18887
rect 37691 18884 37703 18887
rect 43993 18887 44051 18893
rect 37691 18856 38516 18884
rect 37691 18853 37703 18856
rect 37645 18847 37703 18853
rect 32677 18819 32735 18825
rect 32677 18816 32689 18819
rect 31996 18788 32689 18816
rect 31996 18776 32002 18788
rect 32677 18785 32689 18788
rect 32723 18785 32735 18819
rect 32677 18779 32735 18785
rect 33413 18819 33471 18825
rect 33413 18785 33425 18819
rect 33459 18816 33471 18819
rect 33689 18819 33747 18825
rect 33689 18816 33701 18819
rect 33459 18788 33701 18816
rect 33459 18785 33471 18788
rect 33413 18779 33471 18785
rect 33689 18785 33701 18788
rect 33735 18785 33747 18819
rect 33689 18779 33747 18785
rect 33781 18819 33839 18825
rect 33781 18785 33793 18819
rect 33827 18816 33839 18819
rect 34514 18816 34520 18828
rect 33827 18788 34520 18816
rect 33827 18785 33839 18788
rect 33781 18779 33839 18785
rect 26602 18748 26608 18760
rect 22379 18720 26608 18748
rect 7469 18683 7527 18689
rect 7469 18649 7481 18683
rect 7515 18680 7527 18683
rect 8665 18683 8723 18689
rect 8665 18680 8677 18683
rect 7515 18652 8677 18680
rect 7515 18649 7527 18652
rect 7469 18643 7527 18649
rect 8665 18649 8677 18652
rect 8711 18680 8723 18683
rect 9214 18680 9220 18692
rect 8711 18652 9220 18680
rect 8711 18649 8723 18652
rect 8665 18643 8723 18649
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 9398 18640 9404 18692
rect 9456 18680 9462 18692
rect 11698 18680 11704 18692
rect 9456 18652 11704 18680
rect 9456 18640 9462 18652
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 22379 18680 22407 18720
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 27798 18708 27804 18760
rect 27856 18748 27862 18760
rect 28261 18751 28319 18757
rect 28261 18748 28273 18751
rect 27856 18720 28273 18748
rect 27856 18708 27862 18720
rect 28261 18717 28273 18720
rect 28307 18717 28319 18751
rect 28261 18711 28319 18717
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18748 32551 18751
rect 33502 18748 33508 18760
rect 32539 18720 33508 18748
rect 32539 18717 32551 18720
rect 32493 18711 32551 18717
rect 33502 18708 33508 18720
rect 33560 18708 33566 18760
rect 33704 18748 33732 18779
rect 34514 18776 34520 18788
rect 34572 18776 34578 18828
rect 35066 18776 35072 18828
rect 35124 18816 35130 18828
rect 35253 18819 35311 18825
rect 35253 18816 35265 18819
rect 35124 18788 35265 18816
rect 35124 18776 35130 18788
rect 35253 18785 35265 18788
rect 35299 18785 35311 18819
rect 35253 18779 35311 18785
rect 36170 18776 36176 18828
rect 36228 18816 36234 18828
rect 36265 18819 36323 18825
rect 36265 18816 36277 18819
rect 36228 18788 36277 18816
rect 36228 18776 36234 18788
rect 36265 18785 36277 18788
rect 36311 18785 36323 18819
rect 36265 18779 36323 18785
rect 38010 18776 38016 18828
rect 38068 18816 38074 18828
rect 38488 18825 38516 18856
rect 43993 18853 44005 18887
rect 44039 18884 44051 18887
rect 44039 18856 45600 18884
rect 44039 18853 44051 18856
rect 43993 18847 44051 18853
rect 38289 18819 38347 18825
rect 38289 18816 38301 18819
rect 38068 18788 38301 18816
rect 38068 18776 38074 18788
rect 38289 18785 38301 18788
rect 38335 18785 38347 18819
rect 38289 18779 38347 18785
rect 38473 18819 38531 18825
rect 38473 18785 38485 18819
rect 38519 18785 38531 18819
rect 38473 18779 38531 18785
rect 44634 18776 44640 18828
rect 44692 18776 44698 18828
rect 45572 18825 45600 18856
rect 45557 18819 45615 18825
rect 45557 18785 45569 18819
rect 45603 18785 45615 18819
rect 45557 18779 45615 18785
rect 46106 18776 46112 18828
rect 46164 18816 46170 18828
rect 46569 18819 46627 18825
rect 46569 18816 46581 18819
rect 46164 18788 46581 18816
rect 46164 18776 46170 18788
rect 46569 18785 46581 18788
rect 46615 18816 46627 18819
rect 47302 18816 47308 18828
rect 46615 18788 47308 18816
rect 46615 18785 46627 18788
rect 46569 18779 46627 18785
rect 47302 18776 47308 18788
rect 47360 18776 47366 18828
rect 57977 18819 58035 18825
rect 57977 18785 57989 18819
rect 58023 18816 58035 18819
rect 58158 18816 58164 18828
rect 58023 18788 58164 18816
rect 58023 18785 58035 18788
rect 57977 18779 58035 18785
rect 58158 18776 58164 18788
rect 58216 18776 58222 18828
rect 38102 18748 38108 18760
rect 33704 18720 38108 18748
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 42426 18708 42432 18760
rect 42484 18748 42490 18760
rect 42613 18751 42671 18757
rect 42613 18748 42625 18751
rect 42484 18720 42625 18748
rect 42484 18708 42490 18720
rect 42613 18717 42625 18720
rect 42659 18717 42671 18751
rect 42613 18711 42671 18717
rect 46385 18751 46443 18757
rect 46385 18717 46397 18751
rect 46431 18748 46443 18751
rect 46658 18748 46664 18760
rect 46431 18720 46664 18748
rect 46431 18717 46443 18720
rect 46385 18711 46443 18717
rect 46658 18708 46664 18720
rect 46716 18708 46722 18760
rect 51810 18708 51816 18760
rect 51868 18708 51874 18760
rect 52454 18708 52460 18760
rect 52512 18708 52518 18760
rect 52546 18708 52552 18760
rect 52604 18748 52610 18760
rect 52825 18751 52883 18757
rect 52825 18748 52837 18751
rect 52604 18720 52837 18748
rect 52604 18708 52610 18720
rect 52825 18717 52837 18720
rect 52871 18717 52883 18751
rect 52825 18711 52883 18717
rect 57146 18708 57152 18760
rect 57204 18708 57210 18760
rect 21652 18652 22407 18680
rect 4706 18612 4712 18624
rect 3896 18584 4712 18612
rect 4706 18572 4712 18584
rect 4764 18572 4770 18624
rect 5629 18615 5687 18621
rect 5629 18581 5641 18615
rect 5675 18612 5687 18615
rect 10686 18612 10692 18624
rect 5675 18584 10692 18612
rect 5675 18581 5687 18584
rect 5629 18575 5687 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 16482 18572 16488 18624
rect 16540 18572 16546 18624
rect 21450 18572 21456 18624
rect 21508 18612 21514 18624
rect 21652 18621 21680 18652
rect 25222 18640 25228 18692
rect 25280 18680 25286 18692
rect 25593 18683 25651 18689
rect 25593 18680 25605 18683
rect 25280 18652 25605 18680
rect 25280 18640 25286 18652
rect 25593 18649 25605 18652
rect 25639 18680 25651 18683
rect 25958 18680 25964 18692
rect 25639 18652 25964 18680
rect 25639 18649 25651 18652
rect 25593 18643 25651 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 32401 18683 32459 18689
rect 32401 18649 32413 18683
rect 32447 18680 32459 18683
rect 32582 18680 32588 18692
rect 32447 18652 32588 18680
rect 32447 18649 32459 18652
rect 32401 18643 32459 18649
rect 32582 18640 32588 18652
rect 32640 18680 32646 18692
rect 33873 18683 33931 18689
rect 33873 18680 33885 18683
rect 32640 18652 33885 18680
rect 32640 18640 32646 18652
rect 33873 18649 33885 18652
rect 33919 18680 33931 18683
rect 36532 18683 36590 18689
rect 33919 18652 34928 18680
rect 33919 18649 33931 18652
rect 33873 18643 33931 18649
rect 34900 18624 34928 18652
rect 36532 18649 36544 18683
rect 36578 18680 36590 18683
rect 37737 18683 37795 18689
rect 37737 18680 37749 18683
rect 36578 18652 37749 18680
rect 36578 18649 36590 18652
rect 36532 18643 36590 18649
rect 37737 18649 37749 18652
rect 37783 18649 37795 18683
rect 37737 18643 37795 18649
rect 42880 18683 42938 18689
rect 42880 18649 42892 18683
rect 42926 18680 42938 18683
rect 44085 18683 44143 18689
rect 44085 18680 44097 18683
rect 42926 18652 44097 18680
rect 42926 18649 42938 18652
rect 42880 18643 42938 18649
rect 44085 18649 44097 18652
rect 44131 18649 44143 18683
rect 44085 18643 44143 18649
rect 21637 18615 21695 18621
rect 21637 18612 21649 18615
rect 21508 18584 21649 18612
rect 21508 18572 21514 18584
rect 21637 18581 21649 18584
rect 21683 18581 21695 18615
rect 21637 18575 21695 18581
rect 21821 18615 21879 18621
rect 21821 18581 21833 18615
rect 21867 18612 21879 18615
rect 22186 18612 22192 18624
rect 21867 18584 22192 18612
rect 21867 18581 21879 18584
rect 21821 18575 21879 18581
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 27430 18572 27436 18624
rect 27488 18572 27494 18624
rect 27522 18572 27528 18624
rect 27580 18612 27586 18624
rect 27893 18615 27951 18621
rect 27893 18612 27905 18615
rect 27580 18584 27905 18612
rect 27580 18572 27586 18584
rect 27893 18581 27905 18584
rect 27939 18581 27951 18615
rect 27893 18575 27951 18581
rect 34698 18572 34704 18624
rect 34756 18572 34762 18624
rect 34882 18572 34888 18624
rect 34940 18572 34946 18624
rect 35618 18572 35624 18624
rect 35676 18612 35682 18624
rect 40402 18612 40408 18624
rect 35676 18584 40408 18612
rect 35676 18572 35682 18584
rect 40402 18572 40408 18584
rect 40460 18572 40466 18624
rect 46474 18572 46480 18624
rect 46532 18572 46538 18624
rect 51166 18572 51172 18624
rect 51224 18572 51230 18624
rect 51902 18572 51908 18624
rect 51960 18572 51966 18624
rect 56594 18572 56600 18624
rect 56652 18572 56658 18624
rect 1104 18522 59040 18544
rect 1104 18470 15394 18522
rect 15446 18470 15458 18522
rect 15510 18470 15522 18522
rect 15574 18470 15586 18522
rect 15638 18470 15650 18522
rect 15702 18470 29838 18522
rect 29890 18470 29902 18522
rect 29954 18470 29966 18522
rect 30018 18470 30030 18522
rect 30082 18470 30094 18522
rect 30146 18470 44282 18522
rect 44334 18470 44346 18522
rect 44398 18470 44410 18522
rect 44462 18470 44474 18522
rect 44526 18470 44538 18522
rect 44590 18470 58726 18522
rect 58778 18470 58790 18522
rect 58842 18470 58854 18522
rect 58906 18470 58918 18522
rect 58970 18470 58982 18522
rect 59034 18470 59040 18522
rect 1104 18448 59040 18470
rect 3329 18411 3387 18417
rect 3329 18377 3341 18411
rect 3375 18408 3387 18411
rect 3510 18408 3516 18420
rect 3375 18380 3516 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 3878 18408 3884 18420
rect 3752 18380 3884 18408
rect 3752 18368 3758 18380
rect 3878 18368 3884 18380
rect 3936 18408 3942 18420
rect 3973 18411 4031 18417
rect 3973 18408 3985 18411
rect 3936 18380 3985 18408
rect 3936 18368 3942 18380
rect 3973 18377 3985 18380
rect 4019 18377 4031 18411
rect 3973 18371 4031 18377
rect 4062 18368 4068 18420
rect 4120 18368 4126 18420
rect 7837 18411 7895 18417
rect 7837 18377 7849 18411
rect 7883 18408 7895 18411
rect 8018 18408 8024 18420
rect 7883 18380 8024 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8110 18368 8116 18420
rect 8168 18368 8174 18420
rect 8297 18411 8355 18417
rect 8297 18377 8309 18411
rect 8343 18408 8355 18411
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 8343 18380 10609 18408
rect 8343 18377 8355 18380
rect 8297 18371 8355 18377
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 10686 18368 10692 18420
rect 10744 18368 10750 18420
rect 17034 18368 17040 18420
rect 17092 18408 17098 18420
rect 20257 18411 20315 18417
rect 20257 18408 20269 18411
rect 17092 18380 20269 18408
rect 17092 18368 17098 18380
rect 20257 18377 20269 18380
rect 20303 18408 20315 18411
rect 20714 18408 20720 18420
rect 20303 18380 20720 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 27246 18368 27252 18420
rect 27304 18408 27310 18420
rect 27341 18411 27399 18417
rect 27341 18408 27353 18411
rect 27304 18380 27353 18408
rect 27304 18368 27310 18380
rect 27341 18377 27353 18380
rect 27387 18377 27399 18411
rect 27341 18371 27399 18377
rect 27430 18368 27436 18420
rect 27488 18368 27494 18420
rect 33781 18411 33839 18417
rect 33781 18377 33793 18411
rect 33827 18408 33839 18411
rect 34514 18408 34520 18420
rect 33827 18380 34520 18408
rect 33827 18377 33839 18380
rect 33781 18371 33839 18377
rect 34514 18368 34520 18380
rect 34572 18368 34578 18420
rect 34885 18411 34943 18417
rect 34885 18377 34897 18411
rect 34931 18408 34943 18411
rect 35802 18408 35808 18420
rect 34931 18380 35808 18408
rect 34931 18377 34943 18380
rect 34885 18371 34943 18377
rect 35802 18368 35808 18380
rect 35860 18368 35866 18420
rect 51810 18368 51816 18420
rect 51868 18368 51874 18420
rect 51902 18368 51908 18420
rect 51960 18368 51966 18420
rect 52546 18368 52552 18420
rect 52604 18408 52610 18420
rect 52917 18411 52975 18417
rect 52917 18408 52929 18411
rect 52604 18380 52929 18408
rect 52604 18368 52610 18380
rect 52917 18377 52929 18380
rect 52963 18377 52975 18411
rect 52917 18371 52975 18377
rect 56597 18411 56655 18417
rect 56597 18377 56609 18411
rect 56643 18408 56655 18411
rect 57146 18408 57152 18420
rect 56643 18380 57152 18408
rect 56643 18377 56655 18380
rect 56597 18371 56655 18377
rect 57146 18368 57152 18380
rect 57204 18368 57210 18420
rect 2216 18343 2274 18349
rect 2216 18309 2228 18343
rect 2262 18340 2274 18343
rect 2774 18340 2780 18352
rect 2262 18312 2780 18340
rect 2262 18309 2274 18312
rect 2216 18303 2274 18309
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 6724 18343 6782 18349
rect 6724 18309 6736 18343
rect 6770 18340 6782 18343
rect 7190 18340 7196 18352
rect 6770 18312 7196 18340
rect 6770 18309 6782 18312
rect 6724 18303 6782 18309
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 1949 18275 2007 18281
rect 1949 18241 1961 18275
rect 1995 18272 2007 18275
rect 2038 18272 2044 18284
rect 1995 18244 2044 18272
rect 1995 18241 2007 18244
rect 1949 18235 2007 18241
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 4430 18232 4436 18284
rect 4488 18272 4494 18284
rect 4488 18244 4844 18272
rect 4488 18232 4494 18244
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4203 18176 4752 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18136 4252 18148
rect 3528 18108 4252 18136
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 3528 18068 3556 18108
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 4724 18080 4752 18176
rect 4816 18136 4844 18244
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 8128 18272 8156 18368
rect 7156 18244 8156 18272
rect 7156 18232 7162 18244
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 6457 18207 6515 18213
rect 6457 18204 6469 18207
rect 5592 18176 6469 18204
rect 5592 18164 5598 18176
rect 6457 18173 6469 18176
rect 6503 18173 6515 18207
rect 8128 18204 8156 18244
rect 9214 18232 9220 18284
rect 9272 18232 9278 18284
rect 10134 18232 10140 18284
rect 10192 18232 10198 18284
rect 27448 18272 27476 18368
rect 50700 18343 50758 18349
rect 50700 18309 50712 18343
rect 50746 18340 50758 18343
rect 51920 18340 51948 18368
rect 50746 18312 51948 18340
rect 50746 18309 50758 18312
rect 50700 18303 50758 18309
rect 27893 18275 27951 18281
rect 27893 18272 27905 18275
rect 27448 18244 27905 18272
rect 27893 18241 27905 18244
rect 27939 18241 27951 18275
rect 27893 18235 27951 18241
rect 33594 18232 33600 18284
rect 33652 18272 33658 18284
rect 34333 18275 34391 18281
rect 34333 18272 34345 18275
rect 33652 18244 34345 18272
rect 33652 18232 33658 18244
rect 34333 18241 34345 18244
rect 34379 18241 34391 18275
rect 34333 18235 34391 18241
rect 39393 18275 39451 18281
rect 39393 18241 39405 18275
rect 39439 18272 39451 18275
rect 39850 18272 39856 18284
rect 39439 18244 39856 18272
rect 39439 18241 39451 18244
rect 39393 18235 39451 18241
rect 39850 18232 39856 18244
rect 39908 18232 39914 18284
rect 50154 18232 50160 18284
rect 50212 18272 50218 18284
rect 50433 18275 50491 18281
rect 50433 18272 50445 18275
rect 50212 18244 50445 18272
rect 50212 18232 50218 18244
rect 50433 18241 50445 18244
rect 50479 18241 50491 18275
rect 50433 18235 50491 18241
rect 56962 18232 56968 18284
rect 57020 18272 57026 18284
rect 57885 18275 57943 18281
rect 57885 18272 57897 18275
rect 57020 18244 57897 18272
rect 57020 18232 57026 18244
rect 57885 18241 57897 18244
rect 57931 18241 57943 18275
rect 57885 18235 57943 18241
rect 9122 18213 9128 18216
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8128 18176 8953 18204
rect 6457 18167 6515 18173
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 9100 18207 9128 18213
rect 9100 18173 9112 18207
rect 9100 18167 9128 18173
rect 9122 18164 9128 18167
rect 9180 18164 9186 18216
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9456 18176 9505 18204
rect 9456 18164 9462 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 9950 18164 9956 18216
rect 10008 18164 10014 18216
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 10919 18176 11376 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 10888 18136 10916 18167
rect 11348 18145 11376 18176
rect 12986 18164 12992 18216
rect 13044 18164 13050 18216
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18204 13323 18207
rect 13354 18204 13360 18216
rect 13311 18176 13360 18204
rect 13311 18173 13323 18176
rect 13265 18167 13323 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 15565 18207 15623 18213
rect 15565 18204 15577 18207
rect 15160 18176 15577 18204
rect 15160 18164 15166 18176
rect 15565 18173 15577 18176
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15804 18176 15853 18204
rect 15804 18164 15810 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 19150 18164 19156 18216
rect 19208 18164 19214 18216
rect 44634 18164 44640 18216
rect 44692 18164 44698 18216
rect 48406 18164 48412 18216
rect 48464 18164 48470 18216
rect 48774 18164 48780 18216
rect 48832 18164 48838 18216
rect 52546 18164 52552 18216
rect 52604 18164 52610 18216
rect 53834 18164 53840 18216
rect 53892 18204 53898 18216
rect 54113 18207 54171 18213
rect 54113 18204 54125 18207
rect 53892 18176 54125 18204
rect 53892 18164 53898 18176
rect 54113 18173 54125 18176
rect 54159 18173 54171 18207
rect 54113 18167 54171 18173
rect 56870 18164 56876 18216
rect 56928 18204 56934 18216
rect 57057 18207 57115 18213
rect 57057 18204 57069 18207
rect 56928 18176 57069 18204
rect 56928 18164 56934 18176
rect 57057 18173 57069 18176
rect 57103 18173 57115 18207
rect 57057 18167 57115 18173
rect 57149 18207 57207 18213
rect 57149 18173 57161 18207
rect 57195 18173 57207 18207
rect 57149 18167 57207 18173
rect 4816 18108 6040 18136
rect 1912 18040 3556 18068
rect 3605 18071 3663 18077
rect 1912 18028 1918 18040
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4338 18068 4344 18080
rect 3651 18040 4344 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 4706 18028 4712 18080
rect 4764 18028 4770 18080
rect 6012 18077 6040 18108
rect 9646 18108 10916 18136
rect 11333 18139 11391 18145
rect 5997 18071 6055 18077
rect 5997 18037 6009 18071
rect 6043 18068 6055 18071
rect 6086 18068 6092 18080
rect 6043 18040 6092 18068
rect 6043 18037 6055 18040
rect 5997 18031 6055 18037
rect 6086 18028 6092 18040
rect 6144 18068 6150 18080
rect 7926 18068 7932 18080
rect 6144 18040 7932 18068
rect 6144 18028 6150 18040
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9646 18068 9674 18108
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 13906 18136 13912 18148
rect 11379 18108 13912 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 22002 18136 22008 18148
rect 20772 18108 22008 18136
rect 20772 18096 20778 18108
rect 22002 18096 22008 18108
rect 22060 18136 22066 18148
rect 26694 18136 26700 18148
rect 22060 18108 26700 18136
rect 22060 18096 22066 18108
rect 26694 18096 26700 18108
rect 26752 18136 26758 18148
rect 27154 18136 27160 18148
rect 26752 18108 27160 18136
rect 26752 18096 26758 18108
rect 27154 18096 27160 18108
rect 27212 18096 27218 18148
rect 45833 18139 45891 18145
rect 45833 18136 45845 18139
rect 40052 18108 45845 18136
rect 40052 18080 40080 18108
rect 45833 18105 45845 18108
rect 45879 18136 45891 18139
rect 46106 18136 46112 18148
rect 45879 18108 46112 18136
rect 45879 18105 45891 18108
rect 45833 18099 45891 18105
rect 46106 18096 46112 18108
rect 46164 18096 46170 18148
rect 56502 18096 56508 18148
rect 56560 18136 56566 18148
rect 57164 18136 57192 18167
rect 57698 18164 57704 18216
rect 57756 18204 57762 18216
rect 58437 18207 58495 18213
rect 58437 18204 58449 18207
rect 57756 18176 58449 18204
rect 57756 18164 57762 18176
rect 58437 18173 58449 18176
rect 58483 18173 58495 18207
rect 58437 18167 58495 18173
rect 56560 18108 57192 18136
rect 56560 18096 56566 18108
rect 8812 18040 9674 18068
rect 8812 18028 8818 18040
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 12437 18071 12495 18077
rect 12437 18037 12449 18071
rect 12483 18068 12495 18071
rect 12618 18068 12624 18080
rect 12483 18040 12624 18068
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14918 18068 14924 18080
rect 13872 18040 14924 18068
rect 13872 18028 13878 18040
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15010 18028 15016 18080
rect 15068 18028 15074 18080
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 16485 18071 16543 18077
rect 16485 18068 16497 18071
rect 16448 18040 16497 18068
rect 16448 18028 16454 18040
rect 16485 18037 16497 18040
rect 16531 18037 16543 18071
rect 16485 18031 16543 18037
rect 19794 18028 19800 18080
rect 19852 18028 19858 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 25222 18068 25228 18080
rect 20956 18040 25228 18068
rect 20956 18028 20962 18040
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 25501 18071 25559 18077
rect 25501 18037 25513 18071
rect 25547 18068 25559 18071
rect 25958 18068 25964 18080
rect 25547 18040 25964 18068
rect 25547 18037 25559 18040
rect 25501 18031 25559 18037
rect 25958 18028 25964 18040
rect 26016 18028 26022 18080
rect 37550 18028 37556 18080
rect 37608 18028 37614 18080
rect 38746 18028 38752 18080
rect 38804 18028 38810 18080
rect 40034 18028 40040 18080
rect 40092 18028 40098 18080
rect 43162 18028 43168 18080
rect 43220 18068 43226 18080
rect 43717 18071 43775 18077
rect 43717 18068 43729 18071
rect 43220 18040 43729 18068
rect 43220 18028 43226 18040
rect 43717 18037 43729 18040
rect 43763 18068 43775 18071
rect 43898 18068 43904 18080
rect 43763 18040 43904 18068
rect 43763 18037 43775 18040
rect 43717 18031 43775 18037
rect 43898 18028 43904 18040
rect 43956 18028 43962 18080
rect 44082 18028 44088 18080
rect 44140 18028 44146 18080
rect 44174 18028 44180 18080
rect 44232 18068 44238 18080
rect 45005 18071 45063 18077
rect 45005 18068 45017 18071
rect 44232 18040 45017 18068
rect 44232 18028 44238 18040
rect 45005 18037 45017 18040
rect 45051 18037 45063 18071
rect 45005 18031 45063 18037
rect 45370 18028 45376 18080
rect 45428 18028 45434 18080
rect 47854 18028 47860 18080
rect 47912 18028 47918 18080
rect 49326 18028 49332 18080
rect 49384 18028 49390 18080
rect 51902 18028 51908 18080
rect 51960 18028 51966 18080
rect 53374 18028 53380 18080
rect 53432 18068 53438 18080
rect 53561 18071 53619 18077
rect 53561 18068 53573 18071
rect 53432 18040 53573 18068
rect 53432 18028 53438 18040
rect 53561 18037 53573 18040
rect 53607 18037 53619 18071
rect 53561 18031 53619 18037
rect 1104 17978 58880 18000
rect 1104 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 22616 17978
rect 22668 17926 22680 17978
rect 22732 17926 22744 17978
rect 22796 17926 22808 17978
rect 22860 17926 22872 17978
rect 22924 17926 37060 17978
rect 37112 17926 37124 17978
rect 37176 17926 37188 17978
rect 37240 17926 37252 17978
rect 37304 17926 37316 17978
rect 37368 17926 51504 17978
rect 51556 17926 51568 17978
rect 51620 17926 51632 17978
rect 51684 17926 51696 17978
rect 51748 17926 51760 17978
rect 51812 17926 58880 17978
rect 1104 17904 58880 17926
rect 3786 17824 3792 17876
rect 3844 17824 3850 17876
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 8570 17864 8576 17876
rect 4764 17836 8576 17864
rect 4764 17824 4770 17836
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 9858 17864 9864 17876
rect 8680 17836 9864 17864
rect 7558 17756 7564 17808
rect 7616 17796 7622 17808
rect 8680 17796 8708 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10008 17836 10701 17864
rect 10008 17824 10014 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 12529 17867 12587 17873
rect 12529 17833 12541 17867
rect 12575 17864 12587 17867
rect 12986 17864 12992 17876
rect 12575 17836 12992 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 14826 17864 14832 17876
rect 13964 17836 14832 17864
rect 13964 17824 13970 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15252 17836 15884 17864
rect 15252 17824 15258 17836
rect 7616 17768 8708 17796
rect 12437 17799 12495 17805
rect 7616 17756 7622 17768
rect 12437 17765 12449 17799
rect 12483 17796 12495 17799
rect 13078 17796 13084 17808
rect 12483 17768 13084 17796
rect 12483 17765 12495 17768
rect 12437 17759 12495 17765
rect 13078 17756 13084 17768
rect 13136 17796 13142 17808
rect 14461 17799 14519 17805
rect 13136 17768 13216 17796
rect 13136 17756 13142 17768
rect 4338 17688 4344 17740
rect 4396 17688 4402 17740
rect 5534 17688 5540 17740
rect 5592 17688 5598 17740
rect 7742 17728 7748 17740
rect 7024 17700 7748 17728
rect 5552 17660 5580 17688
rect 7024 17669 7052 17700
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 9030 17728 9036 17740
rect 7800 17700 9036 17728
rect 7800 17688 7806 17700
rect 9030 17688 9036 17700
rect 9088 17728 9094 17740
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 9088 17700 9229 17728
rect 9088 17688 9094 17700
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 12526 17728 12532 17740
rect 9217 17691 9275 17697
rect 10244 17700 12532 17728
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 5552 17632 7021 17660
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7009 17623 7067 17629
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17629 8815 17663
rect 9232 17660 9260 17691
rect 10244 17660 10272 17700
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 13188 17737 13216 17768
rect 14461 17765 14473 17799
rect 14507 17765 14519 17799
rect 14461 17759 14519 17765
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17728 13231 17731
rect 13538 17728 13544 17740
rect 13219 17700 13544 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 9232 17632 10272 17660
rect 10612 17632 11253 17660
rect 8757 17623 8815 17629
rect 5804 17595 5862 17601
rect 5804 17561 5816 17595
rect 5850 17592 5862 17595
rect 6270 17592 6276 17604
rect 5850 17564 6276 17592
rect 5850 17561 5862 17564
rect 5804 17555 5862 17561
rect 6270 17552 6276 17564
rect 6328 17552 6334 17604
rect 8772 17536 8800 17623
rect 9490 17601 9496 17604
rect 9484 17555 9496 17601
rect 9490 17552 9496 17555
rect 9548 17552 9554 17604
rect 6914 17484 6920 17536
rect 6972 17484 6978 17536
rect 8754 17484 8760 17536
rect 8812 17484 8818 17536
rect 10612 17533 10640 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17660 12955 17663
rect 13814 17660 13820 17672
rect 12943 17632 13820 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14476 17660 14504 17759
rect 15856 17737 15884 17836
rect 25222 17824 25228 17876
rect 25280 17864 25286 17876
rect 26050 17864 26056 17876
rect 25280 17836 26056 17864
rect 25280 17824 25286 17836
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 47857 17867 47915 17873
rect 47857 17833 47869 17867
rect 47903 17864 47915 17867
rect 48406 17864 48412 17876
rect 47903 17836 48412 17864
rect 47903 17833 47915 17836
rect 47857 17827 47915 17833
rect 48406 17824 48412 17836
rect 48464 17824 48470 17876
rect 51629 17867 51687 17873
rect 48516 17836 51212 17864
rect 37550 17756 37556 17808
rect 37608 17796 37614 17808
rect 40034 17796 40040 17808
rect 37608 17768 40040 17796
rect 37608 17756 37614 17768
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17728 15899 17731
rect 17310 17728 17316 17740
rect 15887 17700 17316 17728
rect 15887 17697 15899 17700
rect 15841 17691 15899 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 37936 17737 37964 17768
rect 40034 17756 40040 17768
rect 40092 17756 40098 17808
rect 43809 17799 43867 17805
rect 43809 17765 43821 17799
rect 43855 17796 43867 17799
rect 48516 17796 48544 17836
rect 43855 17768 43944 17796
rect 43855 17765 43867 17768
rect 43809 17759 43867 17765
rect 43916 17737 43944 17768
rect 47780 17768 48581 17796
rect 47780 17740 47808 17768
rect 37921 17731 37979 17737
rect 37921 17697 37933 17731
rect 37967 17697 37979 17731
rect 43901 17731 43959 17737
rect 37921 17691 37979 17697
rect 39684 17700 42564 17728
rect 15746 17660 15752 17672
rect 14476 17632 15752 17660
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 16758 17620 16764 17672
rect 16816 17620 16822 17672
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 18966 17620 18972 17672
rect 19024 17620 19030 17672
rect 20254 17620 20260 17672
rect 20312 17620 20318 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21634 17620 21640 17672
rect 21692 17620 21698 17672
rect 25866 17620 25872 17672
rect 25924 17620 25930 17672
rect 26234 17620 26240 17672
rect 26292 17660 26298 17672
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 26292 17632 26617 17660
rect 26292 17620 26298 17632
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 26605 17623 26663 17629
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 30432 17632 30573 17660
rect 30432 17620 30438 17632
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 30834 17620 30840 17672
rect 30892 17620 30898 17672
rect 33042 17620 33048 17672
rect 33100 17620 33106 17672
rect 33778 17620 33784 17672
rect 33836 17620 33842 17672
rect 36354 17620 36360 17672
rect 36412 17620 36418 17672
rect 36630 17620 36636 17672
rect 36688 17620 36694 17672
rect 37645 17663 37703 17669
rect 37645 17629 37657 17663
rect 37691 17660 37703 17663
rect 38746 17660 38752 17672
rect 37691 17632 38752 17660
rect 37691 17629 37703 17632
rect 37645 17623 37703 17629
rect 38746 17620 38752 17632
rect 38804 17620 38810 17672
rect 15596 17595 15654 17601
rect 15596 17561 15608 17595
rect 15642 17592 15654 17595
rect 16209 17595 16267 17601
rect 16209 17592 16221 17595
rect 15642 17564 16221 17592
rect 15642 17561 15654 17564
rect 15596 17555 15654 17561
rect 16209 17561 16221 17564
rect 16255 17561 16267 17595
rect 16209 17555 16267 17561
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 23382 17592 23388 17604
rect 18104 17564 23388 17592
rect 18104 17552 18110 17564
rect 23382 17552 23388 17564
rect 23440 17552 23446 17604
rect 37182 17552 37188 17604
rect 37240 17592 37246 17604
rect 37240 17564 38608 17592
rect 37240 17552 37246 17564
rect 38580 17536 38608 17564
rect 39684 17536 39712 17700
rect 40402 17620 40408 17672
rect 40460 17620 40466 17672
rect 41138 17620 41144 17672
rect 41196 17620 41202 17672
rect 41322 17620 41328 17672
rect 41380 17620 41386 17672
rect 41877 17663 41935 17669
rect 41877 17629 41889 17663
rect 41923 17629 41935 17663
rect 41877 17623 41935 17629
rect 40126 17552 40132 17604
rect 40184 17592 40190 17604
rect 41892 17592 41920 17623
rect 42426 17620 42432 17672
rect 42484 17620 42490 17672
rect 42536 17660 42564 17700
rect 43901 17697 43913 17731
rect 43947 17697 43959 17731
rect 45370 17728 45376 17740
rect 43901 17691 43959 17697
rect 44008 17700 45376 17728
rect 44008 17660 44036 17700
rect 45370 17688 45376 17700
rect 45428 17688 45434 17740
rect 47762 17688 47768 17740
rect 47820 17688 47826 17740
rect 48516 17737 48544 17768
rect 48682 17756 48688 17808
rect 48740 17756 48746 17808
rect 50154 17796 50160 17808
rect 49068 17768 50160 17796
rect 48501 17731 48559 17737
rect 48501 17697 48513 17731
rect 48547 17697 48559 17731
rect 48501 17691 48559 17697
rect 42536 17632 44036 17660
rect 44818 17620 44824 17672
rect 44876 17660 44882 17672
rect 45005 17663 45063 17669
rect 45005 17660 45017 17663
rect 44876 17632 45017 17660
rect 44876 17620 44882 17632
rect 45005 17629 45017 17632
rect 45051 17629 45063 17663
rect 45005 17623 45063 17629
rect 47670 17620 47676 17672
rect 47728 17660 47734 17672
rect 48958 17660 48964 17672
rect 47728 17632 48964 17660
rect 47728 17620 47734 17632
rect 48958 17620 48964 17632
rect 49016 17620 49022 17672
rect 49068 17669 49096 17768
rect 50154 17756 50160 17768
rect 50212 17756 50218 17808
rect 49234 17688 49240 17740
rect 49292 17728 49298 17740
rect 49697 17731 49755 17737
rect 49697 17728 49709 17731
rect 49292 17700 49709 17728
rect 49292 17688 49298 17700
rect 49697 17697 49709 17700
rect 49743 17697 49755 17731
rect 51184 17728 51212 17836
rect 51629 17833 51641 17867
rect 51675 17864 51687 17867
rect 52546 17864 52552 17876
rect 51675 17836 52552 17864
rect 51675 17833 51687 17836
rect 51629 17827 51687 17833
rect 52546 17824 52552 17836
rect 52604 17824 52610 17876
rect 53653 17867 53711 17873
rect 53653 17833 53665 17867
rect 53699 17864 53711 17867
rect 53834 17864 53840 17876
rect 53699 17836 53840 17864
rect 53699 17833 53711 17836
rect 53653 17827 53711 17833
rect 53834 17824 53840 17836
rect 53892 17824 53898 17876
rect 57698 17824 57704 17876
rect 57756 17824 57762 17876
rect 51537 17799 51595 17805
rect 51537 17765 51549 17799
rect 51583 17796 51595 17799
rect 51583 17768 53052 17796
rect 51583 17765 51595 17768
rect 51537 17759 51595 17765
rect 52273 17731 52331 17737
rect 51184 17700 52040 17728
rect 49697 17691 49755 17697
rect 49053 17663 49111 17669
rect 49053 17629 49065 17663
rect 49099 17629 49111 17663
rect 49053 17623 49111 17629
rect 49142 17620 49148 17672
rect 49200 17660 49206 17672
rect 50157 17663 50215 17669
rect 50157 17660 50169 17663
rect 49200 17632 50169 17660
rect 49200 17620 49206 17632
rect 50157 17629 50169 17632
rect 50203 17629 50215 17663
rect 50157 17623 50215 17629
rect 50424 17663 50482 17669
rect 50424 17629 50436 17663
rect 50470 17660 50482 17663
rect 51902 17660 51908 17672
rect 50470 17632 51908 17660
rect 50470 17629 50482 17632
rect 50424 17623 50482 17629
rect 51902 17620 51908 17632
rect 51960 17620 51966 17672
rect 52012 17660 52040 17700
rect 52273 17697 52285 17731
rect 52319 17728 52331 17731
rect 52546 17728 52552 17740
rect 52319 17700 52552 17728
rect 52319 17697 52331 17700
rect 52273 17691 52331 17697
rect 52546 17688 52552 17700
rect 52604 17688 52610 17740
rect 53024 17737 53052 17768
rect 53009 17731 53067 17737
rect 53009 17697 53021 17731
rect 53055 17697 53067 17731
rect 53009 17691 53067 17697
rect 53561 17731 53619 17737
rect 53561 17697 53573 17731
rect 53607 17728 53619 17731
rect 54205 17731 54263 17737
rect 54205 17728 54217 17731
rect 53607 17700 54217 17728
rect 53607 17697 53619 17700
rect 53561 17691 53619 17697
rect 54205 17697 54217 17700
rect 54251 17697 54263 17731
rect 54205 17691 54263 17697
rect 53576 17660 53604 17691
rect 56226 17688 56232 17740
rect 56284 17728 56290 17740
rect 56321 17731 56379 17737
rect 56321 17728 56333 17731
rect 56284 17700 56333 17728
rect 56284 17688 56290 17700
rect 56321 17697 56333 17700
rect 56367 17697 56379 17731
rect 56321 17691 56379 17697
rect 52012 17632 53604 17660
rect 54478 17620 54484 17672
rect 54536 17620 54542 17672
rect 56594 17669 56600 17672
rect 56588 17660 56600 17669
rect 56555 17632 56600 17660
rect 56588 17623 56600 17632
rect 56594 17620 56600 17623
rect 56652 17620 56658 17672
rect 40184 17564 41920 17592
rect 42696 17595 42754 17601
rect 40184 17552 40190 17564
rect 42696 17561 42708 17595
rect 42742 17592 42754 17595
rect 43254 17592 43260 17604
rect 42742 17564 43260 17592
rect 42742 17561 42754 17564
rect 42696 17555 42754 17561
rect 43254 17552 43260 17564
rect 43312 17552 43318 17604
rect 48225 17595 48283 17601
rect 48225 17561 48237 17595
rect 48271 17592 48283 17595
rect 49326 17592 49332 17604
rect 48271 17564 49332 17592
rect 48271 17561 48283 17564
rect 48225 17555 48283 17561
rect 49326 17552 49332 17564
rect 49384 17552 49390 17604
rect 54021 17595 54079 17601
rect 54021 17561 54033 17595
rect 54067 17592 54079 17595
rect 55125 17595 55183 17601
rect 55125 17592 55137 17595
rect 54067 17564 55137 17592
rect 54067 17561 54079 17564
rect 54021 17555 54079 17561
rect 55125 17561 55137 17564
rect 55171 17592 55183 17595
rect 55950 17592 55956 17604
rect 55171 17564 55956 17592
rect 55171 17561 55183 17564
rect 55125 17555 55183 17561
rect 55950 17552 55956 17564
rect 56008 17552 56014 17604
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17493 10655 17527
rect 10597 17487 10655 17493
rect 12989 17527 13047 17533
rect 12989 17493 13001 17527
rect 13035 17524 13047 17527
rect 13906 17524 13912 17536
rect 13035 17496 13912 17524
rect 13035 17493 13047 17496
rect 12989 17487 13047 17493
rect 13906 17484 13912 17496
rect 13964 17484 13970 17536
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 18417 17527 18475 17533
rect 18417 17493 18429 17527
rect 18463 17524 18475 17527
rect 18506 17524 18512 17536
rect 18463 17496 18512 17524
rect 18463 17493 18475 17496
rect 18417 17487 18475 17493
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 19610 17484 19616 17536
rect 19668 17484 19674 17536
rect 20346 17484 20352 17536
rect 20404 17484 20410 17536
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 20864 17496 21097 17524
rect 20864 17484 20870 17496
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 25314 17484 25320 17536
rect 25372 17484 25378 17536
rect 26053 17527 26111 17533
rect 26053 17493 26065 17527
rect 26099 17524 26111 17527
rect 26326 17524 26332 17536
rect 26099 17496 26332 17524
rect 26099 17493 26111 17496
rect 26053 17487 26111 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 29730 17484 29736 17536
rect 29788 17524 29794 17536
rect 30009 17527 30067 17533
rect 30009 17524 30021 17527
rect 29788 17496 30021 17524
rect 29788 17484 29794 17496
rect 30009 17493 30021 17496
rect 30055 17493 30067 17527
rect 30009 17487 30067 17493
rect 31202 17484 31208 17536
rect 31260 17524 31266 17536
rect 31389 17527 31447 17533
rect 31389 17524 31401 17527
rect 31260 17496 31401 17524
rect 31260 17484 31266 17496
rect 31389 17493 31401 17496
rect 31435 17493 31447 17527
rect 31389 17487 31447 17493
rect 33134 17484 33140 17536
rect 33192 17524 33198 17536
rect 33689 17527 33747 17533
rect 33689 17524 33701 17527
rect 33192 17496 33701 17524
rect 33192 17484 33198 17496
rect 33689 17493 33701 17496
rect 33735 17493 33747 17527
rect 33689 17487 33747 17493
rect 34422 17484 34428 17536
rect 34480 17484 34486 17536
rect 35710 17484 35716 17536
rect 35768 17524 35774 17536
rect 35805 17527 35863 17533
rect 35805 17524 35817 17527
rect 35768 17496 35817 17524
rect 35768 17484 35774 17496
rect 35805 17493 35817 17496
rect 35851 17493 35863 17527
rect 35805 17487 35863 17493
rect 37277 17527 37335 17533
rect 37277 17493 37289 17527
rect 37323 17524 37335 17527
rect 37366 17524 37372 17536
rect 37323 17496 37372 17524
rect 37323 17493 37335 17496
rect 37277 17487 37335 17493
rect 37366 17484 37372 17496
rect 37424 17484 37430 17536
rect 37737 17527 37795 17533
rect 37737 17493 37749 17527
rect 37783 17524 37795 17527
rect 38378 17524 38384 17536
rect 37783 17496 38384 17524
rect 37783 17493 37795 17496
rect 37737 17487 37795 17493
rect 38378 17484 38384 17496
rect 38436 17484 38442 17536
rect 38562 17484 38568 17536
rect 38620 17484 38626 17536
rect 39666 17484 39672 17536
rect 39724 17484 39730 17536
rect 39850 17484 39856 17536
rect 39908 17484 39914 17536
rect 40586 17484 40592 17536
rect 40644 17484 40650 17536
rect 40678 17484 40684 17536
rect 40736 17524 40742 17536
rect 44174 17524 44180 17536
rect 40736 17496 44180 17524
rect 40736 17484 40742 17496
rect 44174 17484 44180 17496
rect 44232 17484 44238 17536
rect 44545 17527 44603 17533
rect 44545 17493 44557 17527
rect 44591 17524 44603 17527
rect 44726 17524 44732 17536
rect 44591 17496 44732 17524
rect 44591 17493 44603 17496
rect 44545 17487 44603 17493
rect 44726 17484 44732 17496
rect 44784 17484 44790 17536
rect 45278 17484 45284 17536
rect 45336 17524 45342 17536
rect 45649 17527 45707 17533
rect 45649 17524 45661 17527
rect 45336 17496 45661 17524
rect 45336 17484 45342 17496
rect 45649 17493 45661 17496
rect 45695 17493 45707 17527
rect 45649 17487 45707 17493
rect 48314 17484 48320 17536
rect 48372 17524 48378 17536
rect 49145 17527 49203 17533
rect 49145 17524 49157 17527
rect 48372 17496 49157 17524
rect 48372 17484 48378 17496
rect 49145 17493 49157 17496
rect 49191 17493 49203 17527
rect 49145 17487 49203 17493
rect 49510 17484 49516 17536
rect 49568 17524 49574 17536
rect 50246 17524 50252 17536
rect 49568 17496 50252 17524
rect 49568 17484 49574 17496
rect 50246 17484 50252 17496
rect 50304 17484 50310 17536
rect 51902 17484 51908 17536
rect 51960 17524 51966 17536
rect 51997 17527 52055 17533
rect 51997 17524 52009 17527
rect 51960 17496 52009 17524
rect 51960 17484 51966 17496
rect 51997 17493 52009 17496
rect 52043 17493 52055 17527
rect 51997 17487 52055 17493
rect 52086 17484 52092 17536
rect 52144 17524 52150 17536
rect 52457 17527 52515 17533
rect 52457 17524 52469 17527
rect 52144 17496 52469 17524
rect 52144 17484 52150 17496
rect 52457 17493 52469 17496
rect 52503 17493 52515 17527
rect 52457 17487 52515 17493
rect 54113 17527 54171 17533
rect 54113 17493 54125 17527
rect 54159 17524 54171 17527
rect 54202 17524 54208 17536
rect 54159 17496 54208 17524
rect 54159 17493 54171 17496
rect 54113 17487 54171 17493
rect 54202 17484 54208 17496
rect 54260 17484 54266 17536
rect 55214 17484 55220 17536
rect 55272 17524 55278 17536
rect 56594 17524 56600 17536
rect 55272 17496 56600 17524
rect 55272 17484 55278 17496
rect 56594 17484 56600 17496
rect 56652 17484 56658 17536
rect 1104 17434 59040 17456
rect 1104 17382 15394 17434
rect 15446 17382 15458 17434
rect 15510 17382 15522 17434
rect 15574 17382 15586 17434
rect 15638 17382 15650 17434
rect 15702 17382 29838 17434
rect 29890 17382 29902 17434
rect 29954 17382 29966 17434
rect 30018 17382 30030 17434
rect 30082 17382 30094 17434
rect 30146 17382 44282 17434
rect 44334 17382 44346 17434
rect 44398 17382 44410 17434
rect 44462 17382 44474 17434
rect 44526 17382 44538 17434
rect 44590 17382 58726 17434
rect 58778 17382 58790 17434
rect 58842 17382 58854 17434
rect 58906 17382 58918 17434
rect 58970 17382 58982 17434
rect 59034 17382 59040 17434
rect 1104 17360 59040 17382
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 4706 17320 4712 17332
rect 4396 17292 4712 17320
rect 4396 17280 4402 17292
rect 4706 17280 4712 17292
rect 4764 17320 4770 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4764 17292 4997 17320
rect 4764 17280 4770 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 6914 17280 6920 17332
rect 6972 17280 6978 17332
rect 7101 17323 7159 17329
rect 7101 17289 7113 17323
rect 7147 17320 7159 17323
rect 8665 17323 8723 17329
rect 7147 17292 8248 17320
rect 7147 17289 7159 17292
rect 7101 17283 7159 17289
rect 6932 17252 6960 17280
rect 8220 17261 8248 17292
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 8754 17320 8760 17332
rect 8711 17292 8760 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 8754 17280 8760 17292
rect 8812 17320 8818 17332
rect 10134 17320 10140 17332
rect 8812 17292 10140 17320
rect 8812 17280 8818 17292
rect 10134 17280 10140 17292
rect 10192 17320 10198 17332
rect 14182 17320 14188 17332
rect 10192 17292 14188 17320
rect 10192 17280 10198 17292
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14274 17280 14280 17332
rect 14332 17320 14338 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 14332 17292 14473 17320
rect 14332 17280 14338 17292
rect 14461 17289 14473 17292
rect 14507 17289 14519 17323
rect 14461 17283 14519 17289
rect 16669 17323 16727 17329
rect 16669 17289 16681 17323
rect 16715 17320 16727 17323
rect 16758 17320 16764 17332
rect 16715 17292 16764 17320
rect 16715 17289 16727 17292
rect 16669 17283 16727 17289
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 18049 17323 18107 17329
rect 18049 17289 18061 17323
rect 18095 17320 18107 17323
rect 18230 17320 18236 17332
rect 18095 17292 18236 17320
rect 18095 17289 18107 17292
rect 18049 17283 18107 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 20162 17320 20168 17332
rect 18564 17292 20168 17320
rect 18564 17280 18570 17292
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 20312 17292 20361 17320
rect 20312 17280 20318 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 20806 17280 20812 17332
rect 20864 17280 20870 17332
rect 20990 17280 20996 17332
rect 21048 17320 21054 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 21048 17292 21189 17320
rect 21048 17280 21054 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 21177 17283 21235 17289
rect 23842 17280 23848 17332
rect 23900 17320 23906 17332
rect 23937 17323 23995 17329
rect 23937 17320 23949 17323
rect 23900 17292 23949 17320
rect 23900 17280 23906 17292
rect 23937 17289 23949 17292
rect 23983 17320 23995 17323
rect 24762 17320 24768 17332
rect 23983 17292 24768 17320
rect 23983 17289 23995 17292
rect 23937 17283 23995 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 25866 17320 25872 17332
rect 25455 17292 25872 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 27338 17280 27344 17332
rect 27396 17280 27402 17332
rect 29730 17280 29736 17332
rect 29788 17280 29794 17332
rect 30834 17280 30840 17332
rect 30892 17320 30898 17332
rect 30929 17323 30987 17329
rect 30929 17320 30941 17323
rect 30892 17292 30941 17320
rect 30892 17280 30898 17292
rect 30929 17289 30941 17292
rect 30975 17289 30987 17323
rect 30929 17283 30987 17289
rect 33505 17323 33563 17329
rect 33505 17289 33517 17323
rect 33551 17320 33563 17323
rect 33778 17320 33784 17332
rect 33551 17292 33784 17320
rect 33551 17289 33563 17292
rect 33505 17283 33563 17289
rect 33778 17280 33784 17292
rect 33836 17280 33842 17332
rect 34333 17323 34391 17329
rect 34333 17289 34345 17323
rect 34379 17320 34391 17323
rect 34698 17320 34704 17332
rect 34379 17292 34704 17320
rect 34379 17289 34391 17292
rect 34333 17283 34391 17289
rect 34698 17280 34704 17292
rect 34756 17280 34762 17332
rect 35897 17323 35955 17329
rect 35897 17289 35909 17323
rect 35943 17320 35955 17323
rect 36354 17320 36360 17332
rect 35943 17292 36360 17320
rect 35943 17289 35955 17292
rect 35897 17283 35955 17289
rect 36354 17280 36360 17292
rect 36412 17280 36418 17332
rect 36722 17280 36728 17332
rect 36780 17320 36786 17332
rect 36909 17323 36967 17329
rect 36909 17320 36921 17323
rect 36780 17292 36921 17320
rect 36780 17280 36786 17292
rect 36909 17289 36921 17292
rect 36955 17289 36967 17323
rect 36909 17283 36967 17289
rect 39669 17323 39727 17329
rect 39669 17289 39681 17323
rect 39715 17320 39727 17323
rect 39850 17320 39856 17332
rect 39715 17292 39856 17320
rect 39715 17289 39727 17292
rect 39669 17283 39727 17289
rect 39850 17280 39856 17292
rect 39908 17280 39914 17332
rect 40126 17280 40132 17332
rect 40184 17280 40190 17332
rect 40957 17323 41015 17329
rect 40957 17289 40969 17323
rect 41003 17320 41015 17323
rect 41138 17320 41144 17332
rect 41003 17292 41144 17320
rect 41003 17289 41015 17292
rect 40957 17283 41015 17289
rect 41138 17280 41144 17292
rect 41196 17280 41202 17332
rect 42245 17323 42303 17329
rect 42245 17289 42257 17323
rect 42291 17320 42303 17323
rect 42518 17320 42524 17332
rect 42291 17292 42524 17320
rect 42291 17289 42303 17292
rect 42245 17283 42303 17289
rect 8205 17255 8263 17261
rect 6932 17224 7604 17252
rect 7576 17193 7604 17224
rect 8205 17221 8217 17255
rect 8251 17252 8263 17255
rect 9122 17252 9128 17264
rect 8251 17224 9128 17252
rect 8251 17221 8263 17224
rect 8205 17215 8263 17221
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 9401 17255 9459 17261
rect 9401 17221 9413 17255
rect 9447 17252 9459 17255
rect 9490 17252 9496 17264
rect 9447 17224 9496 17252
rect 9447 17221 9459 17224
rect 9401 17215 9459 17221
rect 9490 17212 9496 17224
rect 9548 17212 9554 17264
rect 9861 17255 9919 17261
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 9950 17252 9956 17264
rect 9907 17224 9956 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 9950 17212 9956 17224
rect 10008 17212 10014 17264
rect 12526 17252 12532 17264
rect 11992 17224 12532 17252
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 10226 17144 10232 17196
rect 10284 17184 10290 17196
rect 11992 17193 12020 17224
rect 12526 17212 12532 17224
rect 12584 17252 12590 17264
rect 14912 17255 14970 17261
rect 12584 17224 14688 17252
rect 12584 17212 12590 17224
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 10284 17156 10885 17184
rect 10284 17144 10290 17156
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12244 17187 12302 17193
rect 12244 17153 12256 17187
rect 12290 17184 12302 17187
rect 12618 17184 12624 17196
rect 12290 17156 12624 17184
rect 12290 17153 12302 17156
rect 12244 17147 12302 17153
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 13814 17144 13820 17196
rect 13872 17144 13878 17196
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 14660 17193 14688 17224
rect 14912 17221 14924 17255
rect 14958 17252 14970 17255
rect 15010 17252 15016 17264
rect 14958 17224 15016 17252
rect 14958 17221 14970 17224
rect 14912 17215 14970 17221
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 17310 17212 17316 17264
rect 17368 17252 17374 17264
rect 19518 17252 19524 17264
rect 17368 17224 19524 17252
rect 17368 17212 17374 17224
rect 14645 17187 14703 17193
rect 13964 17156 14596 17184
rect 13964 17144 13970 17156
rect 3970 17076 3976 17128
rect 4028 17076 4034 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17085 7251 17119
rect 7193 17079 7251 17085
rect 4706 17008 4712 17060
rect 4764 17048 4770 17060
rect 5258 17048 5264 17060
rect 4764 17020 5264 17048
rect 4764 17008 4770 17020
rect 5258 17008 5264 17020
rect 5316 17048 5322 17060
rect 7208 17048 7236 17079
rect 7374 17076 7380 17128
rect 7432 17076 7438 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 8895 17088 9536 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 7558 17048 7564 17060
rect 5316 17020 6868 17048
rect 7208 17020 7564 17048
rect 5316 17008 5322 17020
rect 3418 16940 3424 16992
rect 3476 16940 3482 16992
rect 6730 16940 6736 16992
rect 6788 16940 6794 16992
rect 6840 16980 6868 17020
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 9508 17057 9536 17088
rect 9950 17076 9956 17128
rect 10008 17076 10014 17128
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10410 17116 10416 17128
rect 10183 17088 10416 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13280 17088 14105 17116
rect 9493 17051 9551 17057
rect 9493 17017 9505 17051
rect 9539 17017 9551 17051
rect 9493 17011 9551 17017
rect 9600 17020 10456 17048
rect 9600 16980 9628 17020
rect 6840 16952 9628 16980
rect 10318 16940 10324 16992
rect 10376 16940 10382 16992
rect 10428 16980 10456 17020
rect 13280 16980 13308 17088
rect 14093 17085 14105 17088
rect 14139 17116 14151 17119
rect 14274 17116 14280 17128
rect 14139 17088 14280 17116
rect 14139 17085 14151 17088
rect 14093 17079 14151 17085
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14568 17116 14596 17156
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 16114 17184 16120 17196
rect 14645 17147 14703 17153
rect 14752 17156 16120 17184
rect 14752 17116 14780 17156
rect 16114 17144 16120 17156
rect 16172 17184 16178 17196
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16172 17156 17049 17184
rect 16172 17144 16178 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 18984 17193 19012 17224
rect 19518 17212 19524 17224
rect 19576 17252 19582 17264
rect 19576 17224 21496 17252
rect 19576 17212 19582 17224
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 19236 17187 19294 17193
rect 19236 17153 19248 17187
rect 19282 17184 19294 17187
rect 19794 17184 19800 17196
rect 19282 17156 19800 17184
rect 19282 17153 19294 17156
rect 19236 17147 19294 17153
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 21468 17184 21496 17224
rect 21542 17212 21548 17264
rect 21600 17252 21606 17264
rect 25958 17252 25964 17264
rect 21600 17224 25964 17252
rect 21600 17212 21606 17224
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26988 17224 29592 17252
rect 26988 17196 27016 17224
rect 29564 17196 29592 17224
rect 21818 17184 21824 17196
rect 21468 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 22094 17193 22100 17196
rect 22077 17187 22100 17193
rect 22077 17153 22089 17187
rect 22077 17147 22100 17153
rect 22094 17144 22100 17147
rect 22152 17144 22158 17196
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17184 24087 17187
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 24075 17156 25053 17184
rect 24075 17153 24087 17156
rect 24029 17147 24087 17153
rect 25041 17153 25053 17156
rect 25087 17184 25099 17187
rect 25406 17184 25412 17196
rect 25087 17156 25412 17184
rect 25087 17153 25099 17156
rect 25041 17147 25099 17153
rect 25406 17144 25412 17156
rect 25464 17144 25470 17196
rect 25777 17187 25835 17193
rect 25777 17153 25789 17187
rect 25823 17153 25835 17187
rect 25777 17147 25835 17153
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17184 25927 17187
rect 25915 17156 26372 17184
rect 25915 17153 25927 17156
rect 25869 17147 25927 17153
rect 14568 17088 14780 17116
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 16390 17116 16396 17128
rect 15988 17088 16396 17116
rect 15988 17076 15994 17088
rect 16390 17076 16396 17088
rect 16448 17116 16454 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 16448 17088 17141 17116
rect 16448 17076 16454 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17085 17279 17119
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17221 17079 17279 17085
rect 18064 17088 18613 17116
rect 13354 17008 13360 17060
rect 13412 17008 13418 17060
rect 17236 17048 17264 17079
rect 16592 17020 17264 17048
rect 16592 16992 16620 17020
rect 18064 16992 18092 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 20640 17116 20668 17144
rect 20579 17088 20668 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 20714 17076 20720 17128
rect 20772 17076 20778 17128
rect 23382 17076 23388 17128
rect 23440 17116 23446 17128
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23440 17088 24133 17116
rect 23440 17076 23446 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24121 17079 24179 17085
rect 24394 17076 24400 17128
rect 24452 17076 24458 17128
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25792 17116 25820 17147
rect 26344 17128 26372 17156
rect 26970 17144 26976 17196
rect 27028 17144 27034 17196
rect 29546 17144 29552 17196
rect 29604 17144 29610 17196
rect 29748 17184 29776 17280
rect 30466 17212 30472 17264
rect 30524 17252 30530 17264
rect 33045 17255 33103 17261
rect 33045 17252 33057 17255
rect 30524 17224 33057 17252
rect 30524 17212 30530 17224
rect 33045 17221 33057 17224
rect 33091 17221 33103 17255
rect 33045 17215 33103 17221
rect 35802 17212 35808 17264
rect 35860 17252 35866 17264
rect 40678 17252 40684 17264
rect 35860 17224 39252 17252
rect 35860 17212 35866 17224
rect 29805 17187 29863 17193
rect 29805 17184 29817 17187
rect 29748 17156 29817 17184
rect 29805 17153 29817 17156
rect 29851 17153 29863 17187
rect 33134 17184 33140 17196
rect 29805 17147 29863 17153
rect 32692 17156 33140 17184
rect 24820 17088 25820 17116
rect 24820 17076 24826 17088
rect 26050 17076 26056 17128
rect 26108 17076 26114 17128
rect 26326 17076 26332 17128
rect 26384 17076 26390 17128
rect 27430 17076 27436 17128
rect 27488 17076 27494 17128
rect 27525 17119 27583 17125
rect 27525 17085 27537 17119
rect 27571 17085 27583 17119
rect 27525 17079 27583 17085
rect 23201 17051 23259 17057
rect 23201 17017 23213 17051
rect 23247 17048 23259 17051
rect 24946 17048 24952 17060
rect 23247 17020 24952 17048
rect 23247 17017 23259 17020
rect 23201 17011 23259 17017
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 26786 17008 26792 17060
rect 26844 17048 26850 17060
rect 27540 17048 27568 17079
rect 28810 17076 28816 17128
rect 28868 17076 28874 17128
rect 29086 17076 29092 17128
rect 29144 17076 29150 17128
rect 31570 17076 31576 17128
rect 31628 17076 31634 17128
rect 29104 17048 29132 17076
rect 31846 17048 31852 17060
rect 26844 17020 29132 17048
rect 30484 17020 31852 17048
rect 26844 17008 26850 17020
rect 10428 16952 13308 16980
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 16022 16940 16028 16992
rect 16080 16940 16086 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 16485 16983 16543 16989
rect 16485 16980 16497 16983
rect 16264 16952 16497 16980
rect 16264 16940 16270 16952
rect 16485 16949 16497 16952
rect 16531 16980 16543 16983
rect 16574 16980 16580 16992
rect 16531 16952 16580 16980
rect 16531 16949 16543 16952
rect 16485 16943 16543 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 17957 16983 18015 16989
rect 17957 16949 17969 16983
rect 18003 16980 18015 16983
rect 18046 16980 18052 16992
rect 18003 16952 18052 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 21542 16980 21548 16992
rect 21048 16952 21548 16980
rect 21048 16940 21054 16952
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 23569 16983 23627 16989
rect 23569 16949 23581 16983
rect 23615 16980 23627 16983
rect 23934 16980 23940 16992
rect 23615 16952 23940 16980
rect 23615 16949 23627 16952
rect 23569 16943 23627 16949
rect 23934 16940 23940 16952
rect 23992 16940 23998 16992
rect 26878 16940 26884 16992
rect 26936 16980 26942 16992
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 26936 16952 26985 16980
rect 26936 16940 26942 16952
rect 26973 16949 26985 16952
rect 27019 16949 27031 16983
rect 26973 16943 27031 16949
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 30484 16980 30512 17020
rect 31846 17008 31852 17020
rect 31904 17008 31910 17060
rect 32692 16992 32720 17156
rect 33134 17144 33140 17156
rect 33192 17144 33198 17196
rect 36265 17187 36323 17193
rect 34164 17156 34376 17184
rect 34164 17125 34192 17156
rect 34348 17128 34376 17156
rect 36265 17153 36277 17187
rect 36311 17184 36323 17187
rect 37182 17184 37188 17196
rect 36311 17156 37188 17184
rect 36311 17153 36323 17156
rect 36265 17147 36323 17153
rect 37182 17144 37188 17156
rect 37240 17144 37246 17196
rect 37292 17193 37320 17224
rect 37277 17187 37335 17193
rect 37277 17153 37289 17187
rect 37323 17153 37335 17187
rect 37277 17147 37335 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37533 17187 37591 17193
rect 37533 17184 37545 17187
rect 37424 17156 37545 17184
rect 37424 17144 37430 17156
rect 37533 17153 37545 17156
rect 37579 17153 37591 17187
rect 37533 17147 37591 17153
rect 39224 17128 39252 17224
rect 39500 17224 40684 17252
rect 39500 17128 39528 17224
rect 40678 17212 40684 17224
rect 40736 17212 40742 17264
rect 42444 17261 42472 17292
rect 42518 17280 42524 17292
rect 42576 17280 42582 17332
rect 44361 17323 44419 17329
rect 44361 17289 44373 17323
rect 44407 17320 44419 17323
rect 44634 17320 44640 17332
rect 44407 17292 44640 17320
rect 44407 17289 44419 17292
rect 44361 17283 44419 17289
rect 44634 17280 44640 17292
rect 44692 17280 44698 17332
rect 44821 17323 44879 17329
rect 44821 17289 44833 17323
rect 44867 17320 44879 17323
rect 45278 17320 45284 17332
rect 44867 17292 45284 17320
rect 44867 17289 44879 17292
rect 44821 17283 44879 17289
rect 45278 17280 45284 17292
rect 45336 17280 45342 17332
rect 45925 17323 45983 17329
rect 45925 17289 45937 17323
rect 45971 17320 45983 17323
rect 45971 17292 46888 17320
rect 45971 17289 45983 17292
rect 45925 17283 45983 17289
rect 42429 17255 42487 17261
rect 42429 17221 42441 17255
rect 42475 17252 42487 17255
rect 42475 17224 42509 17252
rect 42475 17221 42487 17224
rect 42429 17215 42487 17221
rect 39761 17187 39819 17193
rect 39761 17184 39773 17187
rect 39592 17156 39773 17184
rect 32953 17119 33011 17125
rect 32953 17085 32965 17119
rect 32999 17116 33011 17119
rect 34149 17119 34207 17125
rect 32999 17088 33916 17116
rect 32999 17085 33011 17088
rect 32953 17079 33011 17085
rect 33888 17048 33916 17088
rect 34149 17085 34161 17119
rect 34195 17085 34207 17119
rect 34149 17079 34207 17085
rect 34238 17076 34244 17128
rect 34296 17076 34302 17128
rect 34330 17076 34336 17128
rect 34388 17076 34394 17128
rect 36357 17119 36415 17125
rect 36357 17085 36369 17119
rect 36403 17085 36415 17119
rect 36357 17079 36415 17085
rect 34790 17048 34796 17060
rect 33888 17020 34796 17048
rect 29512 16952 30512 16980
rect 29512 16940 29518 16952
rect 30926 16940 30932 16992
rect 30984 16980 30990 16992
rect 31021 16983 31079 16989
rect 31021 16980 31033 16983
rect 30984 16952 31033 16980
rect 30984 16940 30990 16952
rect 31021 16949 31033 16952
rect 31067 16949 31079 16983
rect 31021 16943 31079 16949
rect 32674 16940 32680 16992
rect 32732 16940 32738 16992
rect 33888 16989 33916 17020
rect 34790 17008 34796 17020
rect 34848 17008 34854 17060
rect 33873 16983 33931 16989
rect 33873 16949 33885 16983
rect 33919 16980 33931 16983
rect 34054 16980 34060 16992
rect 33919 16952 34060 16980
rect 33919 16949 33931 16952
rect 33873 16943 33931 16949
rect 34054 16940 34060 16952
rect 34112 16940 34118 16992
rect 34698 16940 34704 16992
rect 34756 16940 34762 16992
rect 35250 16940 35256 16992
rect 35308 16980 35314 16992
rect 35713 16983 35771 16989
rect 35713 16980 35725 16983
rect 35308 16952 35725 16980
rect 35308 16940 35314 16952
rect 35713 16949 35725 16952
rect 35759 16980 35771 16983
rect 35894 16980 35900 16992
rect 35759 16952 35900 16980
rect 35759 16949 35771 16952
rect 35713 16943 35771 16949
rect 35894 16940 35900 16952
rect 35952 16980 35958 16992
rect 36262 16980 36268 16992
rect 35952 16952 36268 16980
rect 35952 16940 35958 16952
rect 36262 16940 36268 16952
rect 36320 16940 36326 16992
rect 36372 16980 36400 17079
rect 36446 17076 36452 17128
rect 36504 17076 36510 17128
rect 39206 17076 39212 17128
rect 39264 17076 39270 17128
rect 39482 17076 39488 17128
rect 39540 17076 39546 17128
rect 39592 17048 39620 17156
rect 39761 17153 39773 17156
rect 39807 17153 39819 17187
rect 39761 17147 39819 17153
rect 40589 17187 40647 17193
rect 40589 17153 40601 17187
rect 40635 17153 40647 17187
rect 40589 17147 40647 17153
rect 39666 17076 39672 17128
rect 39724 17116 39730 17128
rect 40313 17119 40371 17125
rect 40313 17116 40325 17119
rect 39724 17088 40325 17116
rect 39724 17076 39730 17088
rect 40313 17085 40325 17088
rect 40359 17085 40371 17119
rect 40313 17079 40371 17085
rect 40497 17119 40555 17125
rect 40497 17085 40509 17119
rect 40543 17085 40555 17119
rect 40497 17079 40555 17085
rect 40512 17048 40540 17079
rect 38580 17020 40540 17048
rect 37458 16980 37464 16992
rect 36372 16952 37464 16980
rect 37458 16940 37464 16952
rect 37516 16980 37522 16992
rect 38580 16980 38608 17020
rect 37516 16952 38608 16980
rect 37516 16940 37522 16952
rect 38654 16940 38660 16992
rect 38712 16940 38718 16992
rect 39114 16940 39120 16992
rect 39172 16980 39178 16992
rect 39209 16983 39267 16989
rect 39209 16980 39221 16983
rect 39172 16952 39221 16980
rect 39172 16940 39178 16952
rect 39209 16949 39221 16952
rect 39255 16980 39267 16983
rect 39390 16980 39396 16992
rect 39255 16952 39396 16980
rect 39255 16949 39267 16952
rect 39209 16943 39267 16949
rect 39390 16940 39396 16952
rect 39448 16940 39454 16992
rect 39482 16940 39488 16992
rect 39540 16980 39546 16992
rect 40604 16980 40632 17147
rect 42794 17144 42800 17196
rect 42852 17184 42858 17196
rect 44729 17187 44787 17193
rect 44729 17184 44741 17187
rect 42852 17156 44741 17184
rect 42852 17144 42858 17156
rect 44729 17153 44741 17156
rect 44775 17184 44787 17187
rect 45465 17187 45523 17193
rect 45465 17184 45477 17187
rect 44775 17156 45477 17184
rect 44775 17153 44787 17156
rect 44729 17147 44787 17153
rect 45465 17153 45477 17156
rect 45511 17153 45523 17187
rect 45465 17147 45523 17153
rect 45554 17144 45560 17196
rect 45612 17184 45618 17196
rect 46753 17187 46811 17193
rect 46753 17184 46765 17187
rect 45612 17156 46765 17184
rect 45612 17144 45618 17156
rect 46753 17153 46765 17156
rect 46799 17153 46811 17187
rect 46753 17147 46811 17153
rect 41506 17076 41512 17128
rect 41564 17116 41570 17128
rect 41601 17119 41659 17125
rect 41601 17116 41613 17119
rect 41564 17088 41613 17116
rect 41564 17076 41570 17088
rect 41601 17085 41613 17088
rect 41647 17085 41659 17119
rect 41601 17079 41659 17085
rect 44174 17076 44180 17128
rect 44232 17116 44238 17128
rect 44913 17119 44971 17125
rect 44913 17116 44925 17119
rect 44232 17088 44925 17116
rect 44232 17076 44238 17088
rect 44913 17085 44925 17088
rect 44959 17085 44971 17119
rect 44913 17079 44971 17085
rect 45370 17076 45376 17128
rect 45428 17116 45434 17128
rect 46661 17119 46719 17125
rect 45428 17088 46244 17116
rect 45428 17076 45434 17088
rect 41049 16983 41107 16989
rect 41049 16980 41061 16983
rect 39540 16952 41061 16980
rect 39540 16940 39546 16952
rect 41049 16949 41061 16952
rect 41095 16949 41107 16983
rect 41049 16943 41107 16949
rect 43717 16983 43775 16989
rect 43717 16949 43729 16983
rect 43763 16980 43775 16983
rect 43806 16980 43812 16992
rect 43763 16952 43812 16980
rect 43763 16949 43775 16952
rect 43717 16943 43775 16949
rect 43806 16940 43812 16952
rect 43864 16940 43870 16992
rect 46014 16940 46020 16992
rect 46072 16940 46078 16992
rect 46216 16980 46244 17088
rect 46661 17085 46673 17119
rect 46707 17116 46719 17119
rect 46860 17116 46888 17292
rect 48774 17280 48780 17332
rect 48832 17320 48838 17332
rect 48961 17323 49019 17329
rect 48961 17320 48973 17323
rect 48832 17292 48973 17320
rect 48832 17280 48838 17292
rect 48961 17289 48973 17292
rect 49007 17289 49019 17323
rect 51813 17323 51871 17329
rect 51813 17320 51825 17323
rect 48961 17283 49019 17289
rect 51184 17292 51825 17320
rect 47854 17261 47860 17264
rect 47848 17252 47860 17261
rect 47815 17224 47860 17252
rect 47848 17215 47860 17224
rect 47854 17212 47860 17215
rect 47912 17212 47918 17264
rect 48590 17212 48596 17264
rect 48648 17252 48654 17264
rect 49234 17252 49240 17264
rect 48648 17224 49240 17252
rect 48648 17212 48654 17224
rect 49234 17212 49240 17224
rect 49292 17212 49298 17264
rect 49329 17255 49387 17261
rect 49329 17221 49341 17255
rect 49375 17252 49387 17255
rect 49510 17252 49516 17264
rect 49375 17224 49516 17252
rect 49375 17221 49387 17224
rect 49329 17215 49387 17221
rect 49510 17212 49516 17224
rect 49568 17212 49574 17264
rect 51184 17196 51212 17292
rect 51813 17289 51825 17292
rect 51859 17289 51871 17323
rect 51813 17283 51871 17289
rect 52086 17280 52092 17332
rect 52144 17280 52150 17332
rect 52181 17323 52239 17329
rect 52181 17289 52193 17323
rect 52227 17320 52239 17323
rect 52454 17320 52460 17332
rect 52227 17292 52460 17320
rect 52227 17289 52239 17292
rect 52181 17283 52239 17289
rect 52454 17280 52460 17292
rect 52512 17280 52518 17332
rect 52564 17292 54248 17320
rect 52104 17252 52132 17280
rect 51368 17224 52132 17252
rect 47581 17187 47639 17193
rect 47581 17153 47593 17187
rect 47627 17184 47639 17187
rect 47670 17184 47676 17196
rect 47627 17156 47676 17184
rect 47627 17153 47639 17156
rect 47581 17147 47639 17153
rect 47670 17144 47676 17156
rect 47728 17144 47734 17196
rect 50154 17144 50160 17196
rect 50212 17144 50218 17196
rect 50430 17144 50436 17196
rect 50488 17144 50494 17196
rect 51166 17144 51172 17196
rect 51224 17144 51230 17196
rect 51368 17193 51396 17224
rect 51353 17187 51411 17193
rect 51353 17153 51365 17187
rect 51399 17153 51411 17187
rect 52564 17184 52592 17292
rect 54220 17252 54248 17292
rect 54478 17280 54484 17332
rect 54536 17280 54542 17332
rect 56502 17320 56508 17332
rect 54588 17292 56508 17320
rect 54588 17252 54616 17292
rect 56502 17280 56508 17292
rect 56560 17280 56566 17332
rect 53116 17224 54156 17252
rect 54220 17224 54616 17252
rect 53116 17193 53144 17224
rect 54128 17196 54156 17224
rect 54938 17212 54944 17264
rect 54996 17252 55002 17264
rect 55214 17252 55220 17264
rect 54996 17224 55220 17252
rect 54996 17212 55002 17224
rect 55214 17212 55220 17224
rect 55272 17212 55278 17264
rect 53374 17193 53380 17196
rect 51353 17147 51411 17153
rect 51644 17156 52592 17184
rect 53101 17187 53159 17193
rect 46707 17088 46888 17116
rect 46707 17085 46719 17088
rect 46661 17079 46719 17085
rect 47026 17076 47032 17128
rect 47084 17116 47090 17128
rect 47305 17119 47363 17125
rect 47305 17116 47317 17119
rect 47084 17088 47317 17116
rect 47084 17076 47090 17088
rect 47305 17085 47317 17088
rect 47351 17085 47363 17119
rect 47305 17079 47363 17085
rect 49326 17076 49332 17128
rect 49384 17116 49390 17128
rect 50295 17119 50353 17125
rect 50295 17116 50307 17119
rect 49384 17088 50307 17116
rect 49384 17076 49390 17088
rect 50295 17085 50307 17088
rect 50341 17085 50353 17119
rect 50295 17079 50353 17085
rect 50614 17076 50620 17128
rect 50672 17116 50678 17128
rect 51644 17125 51672 17156
rect 53101 17153 53113 17187
rect 53147 17153 53159 17187
rect 53368 17184 53380 17193
rect 53335 17156 53380 17184
rect 53101 17147 53159 17153
rect 53368 17147 53380 17156
rect 53374 17144 53380 17147
rect 53432 17144 53438 17196
rect 54110 17144 54116 17196
rect 54168 17144 54174 17196
rect 55950 17144 55956 17196
rect 56008 17193 56014 17196
rect 56008 17187 56057 17193
rect 56008 17153 56011 17187
rect 56045 17153 56057 17187
rect 56008 17147 56057 17153
rect 56873 17187 56931 17193
rect 56873 17153 56885 17187
rect 56919 17184 56931 17187
rect 56962 17184 56968 17196
rect 56919 17156 56968 17184
rect 56919 17153 56931 17156
rect 56873 17147 56931 17153
rect 56008 17144 56014 17147
rect 56962 17144 56968 17156
rect 57020 17144 57026 17196
rect 50709 17119 50767 17125
rect 50709 17116 50721 17119
rect 50672 17088 50721 17116
rect 50672 17076 50678 17088
rect 50709 17085 50721 17088
rect 50755 17085 50767 17119
rect 50709 17079 50767 17085
rect 51629 17119 51687 17125
rect 51629 17085 51641 17119
rect 51675 17085 51687 17119
rect 51629 17079 51687 17085
rect 51721 17119 51779 17125
rect 51721 17085 51733 17119
rect 51767 17116 51779 17119
rect 51902 17116 51908 17128
rect 51767 17088 51908 17116
rect 51767 17085 51779 17088
rect 51721 17079 51779 17085
rect 51350 17008 51356 17060
rect 51408 17048 51414 17060
rect 51644 17048 51672 17079
rect 51902 17076 51908 17088
rect 51960 17116 51966 17128
rect 52178 17116 52184 17128
rect 51960 17088 52184 17116
rect 51960 17076 51966 17088
rect 52178 17076 52184 17088
rect 52236 17076 52242 17128
rect 55490 17076 55496 17128
rect 55548 17116 55554 17128
rect 55861 17119 55919 17125
rect 55861 17116 55873 17119
rect 55548 17088 55873 17116
rect 55548 17076 55554 17088
rect 55861 17085 55873 17088
rect 55907 17085 55919 17119
rect 55861 17079 55919 17085
rect 56137 17119 56195 17125
rect 56137 17085 56149 17119
rect 56183 17116 56195 17119
rect 56318 17116 56324 17128
rect 56183 17088 56324 17116
rect 56183 17085 56195 17088
rect 56137 17079 56195 17085
rect 56318 17076 56324 17088
rect 56376 17076 56382 17128
rect 56413 17119 56471 17125
rect 56413 17085 56425 17119
rect 56459 17116 56471 17119
rect 56502 17116 56508 17128
rect 56459 17088 56508 17116
rect 56459 17085 56471 17088
rect 56413 17079 56471 17085
rect 56502 17076 56508 17088
rect 56560 17076 56566 17128
rect 57054 17076 57060 17128
rect 57112 17076 57118 17128
rect 55398 17048 55404 17060
rect 51408 17020 51672 17048
rect 54312 17020 55404 17048
rect 51408 17008 51414 17020
rect 48774 16980 48780 16992
rect 46216 16952 48780 16980
rect 48774 16940 48780 16952
rect 48832 16940 48838 16992
rect 49513 16983 49571 16989
rect 49513 16949 49525 16983
rect 49559 16980 49571 16983
rect 50246 16980 50252 16992
rect 49559 16952 50252 16980
rect 49559 16949 49571 16952
rect 49513 16943 49571 16949
rect 50246 16940 50252 16952
rect 50304 16940 50310 16992
rect 52546 16940 52552 16992
rect 52604 16980 52610 16992
rect 54312 16980 54340 17020
rect 55398 17008 55404 17020
rect 55456 17008 55462 17060
rect 52604 16952 54340 16980
rect 55217 16983 55275 16989
rect 52604 16940 52610 16952
rect 55217 16949 55229 16983
rect 55263 16980 55275 16983
rect 56502 16980 56508 16992
rect 55263 16952 56508 16980
rect 55263 16949 55275 16952
rect 55217 16943 55275 16949
rect 56502 16940 56508 16952
rect 56560 16940 56566 16992
rect 1104 16890 58880 16912
rect 1104 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 22616 16890
rect 22668 16838 22680 16890
rect 22732 16838 22744 16890
rect 22796 16838 22808 16890
rect 22860 16838 22872 16890
rect 22924 16838 37060 16890
rect 37112 16838 37124 16890
rect 37176 16838 37188 16890
rect 37240 16838 37252 16890
rect 37304 16838 37316 16890
rect 37368 16838 51504 16890
rect 51556 16838 51568 16890
rect 51620 16838 51632 16890
rect 51684 16838 51696 16890
rect 51748 16838 51760 16890
rect 51812 16838 58880 16890
rect 1104 16816 58880 16838
rect 6270 16736 6276 16788
rect 6328 16736 6334 16788
rect 6730 16736 6736 16788
rect 6788 16736 6794 16788
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 7432 16748 7573 16776
rect 7432 16736 7438 16748
rect 7561 16745 7573 16748
rect 7607 16745 7619 16779
rect 7561 16739 7619 16745
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 12526 16776 12532 16788
rect 11900 16748 12532 16776
rect 3789 16711 3847 16717
rect 3789 16677 3801 16711
rect 3835 16677 3847 16711
rect 3789 16671 3847 16677
rect 3605 16643 3663 16649
rect 3605 16609 3617 16643
rect 3651 16640 3663 16643
rect 3804 16640 3832 16671
rect 3651 16612 3832 16640
rect 3651 16609 3663 16612
rect 3605 16603 3663 16609
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 4212 16612 4261 16640
rect 4212 16600 4218 16612
rect 4249 16609 4261 16612
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4706 16640 4712 16652
rect 4479 16612 4712 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 6748 16640 6776 16736
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6748 16612 6837 16640
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 9766 16600 9772 16652
rect 9824 16600 9830 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10686 16640 10692 16652
rect 9999 16612 10692 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 11900 16649 11928 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 18966 16776 18972 16788
rect 18831 16748 18972 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 19702 16776 19708 16788
rect 19291 16748 19708 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20806 16736 20812 16788
rect 20864 16736 20870 16788
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 21876 16748 22477 16776
rect 21876 16736 21882 16748
rect 22465 16745 22477 16748
rect 22511 16776 22523 16779
rect 22554 16776 22560 16788
rect 22511 16748 22560 16776
rect 22511 16745 22523 16748
rect 22465 16739 22523 16745
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 26234 16736 26240 16788
rect 26292 16736 26298 16788
rect 26970 16776 26976 16788
rect 26620 16748 26976 16776
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10836 16612 11069 16640
rect 10836 16600 10842 16612
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16640 13967 16643
rect 14090 16640 14096 16652
rect 13955 16612 14096 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14090 16600 14096 16612
rect 14148 16640 14154 16652
rect 14918 16649 14924 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14148 16612 14749 16640
rect 14148 16600 14154 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14896 16643 14924 16649
rect 14896 16609 14908 16643
rect 14896 16603 14924 16609
rect 14918 16600 14924 16603
rect 14976 16600 14982 16652
rect 15286 16600 15292 16652
rect 15344 16600 15350 16652
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 16040 16640 16068 16736
rect 19058 16668 19064 16720
rect 19116 16708 19122 16720
rect 19116 16680 19564 16708
rect 19116 16668 19122 16680
rect 16577 16643 16635 16649
rect 16577 16640 16589 16643
rect 16040 16612 16589 16640
rect 16577 16609 16589 16612
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 17368 16612 17417 16640
rect 17368 16600 17374 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 19536 16640 19564 16680
rect 20027 16643 20085 16649
rect 20027 16640 20039 16643
rect 19536 16612 20039 16640
rect 17405 16603 17463 16609
rect 20027 16609 20039 16612
rect 20073 16609 20085 16643
rect 20027 16603 20085 16609
rect 20162 16600 20168 16652
rect 20220 16600 20226 16652
rect 20438 16600 20444 16652
rect 20496 16600 20502 16652
rect 20824 16640 20852 16736
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20824 16612 20913 16640
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 21085 16643 21143 16649
rect 21085 16640 21097 16643
rect 20901 16603 20959 16609
rect 21008 16612 21097 16640
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10318 16572 10324 16584
rect 9723 16544 10324 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 17678 16581 17684 16584
rect 17672 16572 17684 16581
rect 15804 16544 16068 16572
rect 17639 16544 17684 16572
rect 15804 16532 15810 16544
rect 4157 16507 4215 16513
rect 4157 16473 4169 16507
rect 4203 16504 4215 16507
rect 4890 16504 4896 16516
rect 4203 16476 4896 16504
rect 4203 16473 4215 16476
rect 4157 16467 4215 16473
rect 4890 16464 4896 16476
rect 4948 16504 4954 16516
rect 5261 16507 5319 16513
rect 5261 16504 5273 16507
rect 4948 16476 5273 16504
rect 4948 16464 4954 16476
rect 5261 16473 5273 16476
rect 5307 16473 5319 16507
rect 5261 16467 5319 16473
rect 12152 16507 12210 16513
rect 12152 16473 12164 16507
rect 12198 16504 12210 16507
rect 12802 16504 12808 16516
rect 12198 16476 12808 16504
rect 12198 16473 12210 16476
rect 12152 16467 12210 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 16040 16513 16068 16544
rect 17672 16535 17684 16544
rect 17678 16532 17684 16535
rect 17736 16532 17742 16584
rect 19886 16532 19892 16584
rect 19944 16532 19950 16584
rect 21008 16572 21036 16612
rect 21085 16609 21097 16612
rect 21131 16609 21143 16643
rect 22572 16640 22600 16736
rect 24854 16640 24860 16652
rect 22572 16612 24860 16640
rect 21085 16603 21143 16609
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 25958 16600 25964 16652
rect 26016 16640 26022 16652
rect 26234 16640 26240 16652
rect 26016 16612 26240 16640
rect 26016 16600 26022 16612
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 26620 16649 26648 16748
rect 26970 16736 26976 16748
rect 27028 16736 27034 16788
rect 29638 16736 29644 16788
rect 29696 16776 29702 16788
rect 29917 16779 29975 16785
rect 29917 16776 29929 16779
rect 29696 16748 29929 16776
rect 29696 16736 29702 16748
rect 29917 16745 29929 16748
rect 29963 16776 29975 16779
rect 30098 16776 30104 16788
rect 29963 16748 30104 16776
rect 29963 16745 29975 16748
rect 29917 16739 29975 16745
rect 30098 16736 30104 16748
rect 30156 16776 30162 16788
rect 30650 16776 30656 16788
rect 30156 16748 30656 16776
rect 30156 16736 30162 16748
rect 30650 16736 30656 16748
rect 30708 16736 30714 16788
rect 30926 16736 30932 16788
rect 30984 16736 30990 16788
rect 32674 16776 32680 16788
rect 31036 16748 32680 16776
rect 26605 16643 26663 16649
rect 26605 16609 26617 16643
rect 26651 16609 26663 16643
rect 26605 16603 26663 16609
rect 28442 16600 28448 16652
rect 28500 16640 28506 16652
rect 29181 16643 29239 16649
rect 29181 16640 29193 16643
rect 28500 16612 29193 16640
rect 28500 16600 28506 16612
rect 29181 16609 29193 16612
rect 29227 16609 29239 16643
rect 29181 16603 29239 16609
rect 30098 16600 30104 16652
rect 30156 16600 30162 16652
rect 30285 16643 30343 16649
rect 30285 16609 30297 16643
rect 30331 16640 30343 16643
rect 30837 16643 30895 16649
rect 30837 16640 30849 16643
rect 30331 16612 30849 16640
rect 30331 16609 30343 16612
rect 30285 16603 30343 16609
rect 30837 16609 30849 16612
rect 30883 16640 30895 16643
rect 30944 16640 30972 16736
rect 31036 16649 31064 16748
rect 32674 16736 32680 16748
rect 32732 16736 32738 16788
rect 32769 16779 32827 16785
rect 32769 16745 32781 16779
rect 32815 16776 32827 16779
rect 33042 16776 33048 16788
rect 32815 16748 33048 16776
rect 32815 16745 32827 16748
rect 32769 16739 32827 16745
rect 33042 16736 33048 16748
rect 33100 16736 33106 16788
rect 33870 16736 33876 16788
rect 33928 16776 33934 16788
rect 33928 16748 34192 16776
rect 33928 16736 33934 16748
rect 31220 16680 31616 16708
rect 31220 16652 31248 16680
rect 30883 16612 30972 16640
rect 31021 16643 31079 16649
rect 30883 16609 30895 16612
rect 30837 16603 30895 16609
rect 31021 16609 31033 16643
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 31202 16600 31208 16652
rect 31260 16600 31266 16652
rect 31478 16600 31484 16652
rect 31536 16600 31542 16652
rect 31588 16640 31616 16680
rect 31757 16643 31815 16649
rect 31757 16640 31769 16643
rect 31588 16612 31769 16640
rect 31757 16609 31769 16612
rect 31803 16609 31815 16643
rect 31757 16603 31815 16609
rect 31846 16600 31852 16652
rect 31904 16649 31910 16652
rect 31904 16643 31932 16649
rect 31920 16609 31932 16643
rect 31904 16603 31932 16609
rect 31904 16600 31910 16603
rect 32674 16600 32680 16652
rect 32732 16600 32738 16652
rect 34164 16649 34192 16748
rect 34330 16736 34336 16788
rect 34388 16776 34394 16788
rect 34517 16779 34575 16785
rect 34517 16776 34529 16779
rect 34388 16748 34529 16776
rect 34388 16736 34394 16748
rect 34517 16745 34529 16748
rect 34563 16776 34575 16779
rect 34563 16748 36584 16776
rect 34563 16745 34575 16748
rect 34517 16739 34575 16745
rect 36556 16708 36584 16748
rect 36630 16736 36636 16788
rect 36688 16776 36694 16788
rect 36817 16779 36875 16785
rect 36817 16776 36829 16779
rect 36688 16748 36829 16776
rect 36688 16736 36694 16748
rect 36817 16745 36829 16748
rect 36863 16745 36875 16779
rect 36817 16739 36875 16745
rect 37550 16736 37556 16788
rect 37608 16736 37614 16788
rect 37829 16779 37887 16785
rect 37829 16745 37841 16779
rect 37875 16776 37887 16779
rect 38930 16776 38936 16788
rect 37875 16748 38936 16776
rect 37875 16745 37887 16748
rect 37829 16739 37887 16745
rect 38930 16736 38936 16748
rect 38988 16736 38994 16788
rect 39206 16736 39212 16788
rect 39264 16776 39270 16788
rect 42426 16776 42432 16788
rect 39264 16748 41276 16776
rect 39264 16736 39270 16748
rect 37568 16708 37596 16736
rect 36556 16680 37596 16708
rect 39022 16668 39028 16720
rect 39080 16668 39086 16720
rect 39850 16668 39856 16720
rect 39908 16668 39914 16720
rect 34149 16643 34207 16649
rect 34149 16609 34161 16643
rect 34195 16609 34207 16643
rect 34149 16603 34207 16609
rect 36722 16600 36728 16652
rect 36780 16640 36786 16652
rect 37001 16643 37059 16649
rect 37001 16640 37013 16643
rect 36780 16612 37013 16640
rect 36780 16600 36786 16612
rect 37001 16609 37013 16612
rect 37047 16609 37059 16643
rect 37001 16603 37059 16609
rect 37185 16643 37243 16649
rect 37185 16609 37197 16643
rect 37231 16640 37243 16643
rect 37458 16640 37464 16652
rect 37231 16612 37464 16640
rect 37231 16609 37243 16612
rect 37185 16603 37243 16609
rect 37458 16600 37464 16612
rect 37516 16600 37522 16652
rect 38286 16600 38292 16652
rect 38344 16640 38350 16652
rect 38344 16612 38516 16640
rect 38344 16600 38350 16612
rect 20916 16544 21036 16572
rect 16025 16507 16083 16513
rect 16025 16473 16037 16507
rect 16071 16473 16083 16507
rect 16025 16467 16083 16473
rect 2958 16396 2964 16448
rect 3016 16396 3022 16448
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 11701 16439 11759 16445
rect 11701 16436 11713 16439
rect 11480 16408 11713 16436
rect 11480 16396 11486 16408
rect 11701 16405 11713 16408
rect 11747 16405 11759 16439
rect 11701 16399 11759 16405
rect 13262 16396 13268 16448
rect 13320 16396 13326 16448
rect 14093 16439 14151 16445
rect 14093 16405 14105 16439
rect 14139 16436 14151 16439
rect 15194 16436 15200 16448
rect 14139 16408 15200 16436
rect 14139 16405 14151 16408
rect 14093 16399 14151 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 20916 16436 20944 16544
rect 23934 16532 23940 16584
rect 23992 16532 23998 16584
rect 26878 16581 26884 16584
rect 26872 16572 26884 16581
rect 26839 16544 26884 16572
rect 26872 16535 26884 16544
rect 26878 16532 26884 16535
rect 26936 16532 26942 16584
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16572 29055 16575
rect 29454 16572 29460 16584
rect 29043 16544 29460 16572
rect 29043 16541 29055 16544
rect 28997 16535 29055 16541
rect 29454 16532 29460 16544
rect 29512 16532 29518 16584
rect 30377 16575 30435 16581
rect 30377 16541 30389 16575
rect 30423 16572 30435 16575
rect 30466 16572 30472 16584
rect 30423 16544 30472 16572
rect 30423 16541 30435 16544
rect 30377 16535 30435 16541
rect 20990 16464 20996 16516
rect 21048 16504 21054 16516
rect 21177 16507 21235 16513
rect 21177 16504 21189 16507
rect 21048 16476 21189 16504
rect 21048 16464 21054 16476
rect 21177 16473 21189 16476
rect 21223 16473 21235 16507
rect 21177 16467 21235 16473
rect 25124 16507 25182 16513
rect 25124 16473 25136 16507
rect 25170 16504 25182 16507
rect 25314 16504 25320 16516
rect 25170 16476 25320 16504
rect 25170 16473 25182 16476
rect 25124 16467 25182 16473
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 29089 16507 29147 16513
rect 29089 16473 29101 16507
rect 29135 16504 29147 16507
rect 30392 16504 30420 16535
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 32030 16532 32036 16584
rect 32088 16532 32094 16584
rect 33893 16575 33951 16581
rect 33893 16541 33905 16575
rect 33939 16572 33951 16575
rect 34422 16572 34428 16584
rect 33939 16544 34428 16572
rect 33939 16541 33951 16544
rect 33893 16535 33951 16541
rect 34422 16532 34428 16544
rect 34480 16532 34486 16584
rect 38488 16581 38516 16612
rect 39482 16600 39488 16652
rect 39540 16600 39546 16652
rect 39669 16643 39727 16649
rect 39669 16609 39681 16643
rect 39715 16640 39727 16643
rect 39868 16640 39896 16668
rect 41248 16649 41276 16748
rect 41708 16748 42432 16776
rect 41708 16649 41736 16748
rect 42426 16736 42432 16748
rect 42484 16776 42490 16788
rect 43806 16776 43812 16788
rect 42484 16748 43812 16776
rect 42484 16736 42490 16748
rect 43456 16649 43484 16748
rect 43806 16736 43812 16748
rect 43864 16776 43870 16788
rect 47670 16776 47676 16788
rect 43864 16748 47676 16776
rect 43864 16736 43870 16748
rect 44818 16668 44824 16720
rect 44876 16668 44882 16720
rect 45020 16649 45048 16748
rect 47320 16649 47348 16748
rect 47670 16736 47676 16748
rect 47728 16736 47734 16788
rect 48774 16736 48780 16788
rect 48832 16776 48838 16788
rect 51350 16776 51356 16788
rect 48832 16748 51356 16776
rect 48832 16736 48838 16748
rect 51350 16736 51356 16748
rect 51408 16736 51414 16788
rect 54110 16776 54116 16788
rect 53392 16748 54116 16776
rect 49789 16711 49847 16717
rect 49789 16677 49801 16711
rect 49835 16708 49847 16711
rect 50062 16708 50068 16720
rect 49835 16680 50068 16708
rect 49835 16677 49847 16680
rect 49789 16671 49847 16677
rect 39715 16612 39896 16640
rect 41233 16643 41291 16649
rect 39715 16609 39727 16612
rect 39669 16603 39727 16609
rect 41233 16609 41245 16643
rect 41279 16640 41291 16643
rect 41693 16643 41751 16649
rect 41693 16640 41705 16643
rect 41279 16612 41705 16640
rect 41279 16609 41291 16612
rect 41233 16603 41291 16609
rect 41693 16609 41705 16612
rect 41739 16609 41751 16643
rect 41693 16603 41751 16609
rect 43441 16643 43499 16649
rect 43441 16609 43453 16643
rect 43487 16609 43499 16643
rect 43441 16603 43499 16609
rect 45005 16643 45063 16649
rect 45005 16609 45017 16643
rect 45051 16609 45063 16643
rect 45005 16603 45063 16609
rect 47305 16643 47363 16649
rect 47305 16609 47317 16643
rect 47351 16609 47363 16643
rect 47305 16603 47363 16609
rect 48682 16600 48688 16652
rect 48740 16640 48746 16652
rect 49329 16643 49387 16649
rect 49329 16640 49341 16643
rect 48740 16612 49341 16640
rect 48740 16600 48746 16612
rect 49329 16609 49341 16612
rect 49375 16609 49387 16643
rect 49329 16603 49387 16609
rect 35437 16575 35495 16581
rect 35437 16541 35449 16575
rect 35483 16572 35495 16575
rect 37277 16575 37335 16581
rect 35483 16544 35848 16572
rect 35483 16541 35495 16544
rect 35437 16535 35495 16541
rect 35820 16516 35848 16544
rect 37277 16541 37289 16575
rect 37323 16541 37335 16575
rect 37277 16535 37335 16541
rect 38473 16575 38531 16581
rect 38473 16541 38485 16575
rect 38519 16541 38531 16575
rect 38473 16535 38531 16541
rect 35710 16513 35716 16516
rect 35704 16504 35716 16513
rect 29135 16476 30420 16504
rect 35671 16476 35716 16504
rect 29135 16473 29147 16476
rect 29089 16467 29147 16473
rect 35704 16467 35716 16476
rect 35710 16464 35716 16467
rect 35768 16464 35774 16516
rect 35802 16464 35808 16516
rect 35860 16464 35866 16516
rect 37292 16504 37320 16535
rect 38562 16532 38568 16584
rect 38620 16581 38626 16584
rect 38620 16575 38669 16581
rect 38620 16541 38623 16575
rect 38657 16541 38669 16575
rect 38620 16535 38669 16541
rect 38620 16532 38626 16535
rect 38746 16532 38752 16584
rect 38804 16532 38810 16584
rect 40402 16532 40408 16584
rect 40460 16532 40466 16584
rect 40977 16575 41035 16581
rect 40977 16541 40989 16575
rect 41023 16572 41035 16575
rect 41322 16572 41328 16584
rect 41023 16544 41328 16572
rect 41023 16541 41035 16544
rect 40977 16535 41035 16541
rect 41322 16532 41328 16544
rect 41380 16532 41386 16584
rect 43708 16575 43766 16581
rect 43708 16541 43720 16575
rect 43754 16572 43766 16575
rect 44082 16572 44088 16584
rect 43754 16544 44088 16572
rect 43754 16541 43766 16544
rect 43708 16535 43766 16541
rect 44082 16532 44088 16544
rect 44140 16532 44146 16584
rect 45272 16575 45330 16581
rect 45272 16541 45284 16575
rect 45318 16572 45330 16575
rect 46014 16572 46020 16584
rect 45318 16544 46020 16572
rect 45318 16541 45330 16544
rect 45272 16535 45330 16541
rect 46014 16532 46020 16544
rect 46072 16532 46078 16584
rect 47026 16532 47032 16584
rect 47084 16532 47090 16584
rect 48130 16532 48136 16584
rect 48188 16572 48194 16584
rect 49804 16572 49832 16671
rect 50062 16668 50068 16680
rect 50120 16668 50126 16720
rect 50706 16600 50712 16652
rect 50764 16640 50770 16652
rect 51445 16643 51503 16649
rect 51445 16640 51457 16643
rect 50764 16612 51457 16640
rect 50764 16600 50770 16612
rect 51445 16609 51457 16612
rect 51491 16609 51503 16643
rect 51445 16603 51503 16609
rect 52362 16600 52368 16652
rect 52420 16640 52426 16652
rect 53392 16649 53420 16748
rect 54110 16736 54116 16748
rect 54168 16736 54174 16788
rect 55125 16779 55183 16785
rect 55125 16745 55137 16779
rect 55171 16776 55183 16779
rect 55490 16776 55496 16788
rect 55171 16748 55496 16776
rect 55171 16745 55183 16748
rect 55125 16739 55183 16745
rect 55490 16736 55496 16748
rect 55548 16736 55554 16788
rect 53377 16643 53435 16649
rect 53377 16640 53389 16643
rect 52420 16612 53389 16640
rect 52420 16600 52426 16612
rect 53377 16609 53389 16612
rect 53423 16609 53435 16643
rect 53377 16603 53435 16609
rect 56134 16600 56140 16652
rect 56192 16600 56198 16652
rect 57146 16600 57152 16652
rect 57204 16640 57210 16652
rect 58161 16643 58219 16649
rect 58161 16640 58173 16643
rect 57204 16612 58173 16640
rect 57204 16600 57210 16612
rect 58161 16609 58173 16612
rect 58207 16609 58219 16643
rect 58161 16603 58219 16609
rect 48188 16544 49832 16572
rect 48188 16532 48194 16544
rect 55858 16532 55864 16584
rect 55916 16532 55922 16584
rect 37292 16476 38056 16504
rect 19668 16408 20944 16436
rect 19668 16396 19674 16408
rect 23382 16396 23388 16448
rect 23440 16396 23446 16448
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16436 24731 16439
rect 24762 16436 24768 16448
rect 24719 16408 24768 16436
rect 24719 16405 24731 16408
rect 24673 16399 24731 16405
rect 24762 16396 24768 16408
rect 24820 16396 24826 16448
rect 27982 16396 27988 16448
rect 28040 16396 28046 16448
rect 28626 16396 28632 16448
rect 28684 16396 28690 16448
rect 30742 16396 30748 16448
rect 30800 16396 30806 16448
rect 37642 16396 37648 16448
rect 37700 16396 37706 16448
rect 38028 16436 38056 16476
rect 38746 16436 38752 16448
rect 38028 16408 38752 16436
rect 38746 16396 38752 16408
rect 38804 16396 38810 16448
rect 39853 16439 39911 16445
rect 39853 16405 39865 16439
rect 39899 16436 39911 16439
rect 40420 16436 40448 16532
rect 41598 16464 41604 16516
rect 41656 16504 41662 16516
rect 41938 16507 41996 16513
rect 41938 16504 41950 16507
rect 41656 16476 41950 16504
rect 41656 16464 41662 16476
rect 41938 16473 41950 16476
rect 41984 16473 41996 16507
rect 41938 16467 41996 16473
rect 39899 16408 40448 16436
rect 39899 16405 39911 16408
rect 39853 16399 39911 16405
rect 43070 16396 43076 16448
rect 43128 16396 43134 16448
rect 46385 16439 46443 16445
rect 46385 16405 46397 16439
rect 46431 16436 46443 16439
rect 47044 16436 47072 16532
rect 47572 16507 47630 16513
rect 47572 16473 47584 16507
rect 47618 16504 47630 16507
rect 48777 16507 48835 16513
rect 48777 16504 48789 16507
rect 47618 16476 48789 16504
rect 47618 16473 47630 16476
rect 47572 16467 47630 16473
rect 48777 16473 48789 16476
rect 48823 16473 48835 16507
rect 48777 16467 48835 16473
rect 53644 16507 53702 16513
rect 53644 16473 53656 16507
rect 53690 16504 53702 16507
rect 55309 16507 55367 16513
rect 55309 16504 55321 16507
rect 53690 16476 55321 16504
rect 53690 16473 53702 16476
rect 53644 16467 53702 16473
rect 55309 16473 55321 16476
rect 55355 16473 55367 16507
rect 55309 16467 55367 16473
rect 56404 16507 56462 16513
rect 56404 16473 56416 16507
rect 56450 16504 56462 16507
rect 57609 16507 57667 16513
rect 57609 16504 57621 16507
rect 56450 16476 57621 16504
rect 56450 16473 56462 16476
rect 56404 16467 56462 16473
rect 57609 16473 57621 16476
rect 57655 16473 57667 16507
rect 57609 16467 57667 16473
rect 46431 16408 47072 16436
rect 46431 16405 46443 16408
rect 46385 16399 46443 16405
rect 48682 16396 48688 16448
rect 48740 16396 48746 16448
rect 52086 16396 52092 16448
rect 52144 16396 52150 16448
rect 54754 16396 54760 16448
rect 54812 16396 54818 16448
rect 57514 16396 57520 16448
rect 57572 16396 57578 16448
rect 1104 16346 59040 16368
rect 1104 16294 15394 16346
rect 15446 16294 15458 16346
rect 15510 16294 15522 16346
rect 15574 16294 15586 16346
rect 15638 16294 15650 16346
rect 15702 16294 29838 16346
rect 29890 16294 29902 16346
rect 29954 16294 29966 16346
rect 30018 16294 30030 16346
rect 30082 16294 30094 16346
rect 30146 16294 44282 16346
rect 44334 16294 44346 16346
rect 44398 16294 44410 16346
rect 44462 16294 44474 16346
rect 44526 16294 44538 16346
rect 44590 16294 58726 16346
rect 58778 16294 58790 16346
rect 58842 16294 58854 16346
rect 58906 16294 58918 16346
rect 58970 16294 58982 16346
rect 59034 16294 59040 16346
rect 1104 16272 59040 16294
rect 2958 16232 2964 16244
rect 2746 16204 2964 16232
rect 2308 16167 2366 16173
rect 2308 16133 2320 16167
rect 2354 16164 2366 16167
rect 2746 16164 2774 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3970 16232 3976 16244
rect 3743 16204 3976 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4065 16235 4123 16241
rect 4065 16201 4077 16235
rect 4111 16232 4123 16235
rect 4154 16232 4160 16244
rect 4111 16204 4160 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4154 16192 4160 16204
rect 4212 16232 4218 16244
rect 4430 16232 4436 16244
rect 4212 16204 4436 16232
rect 4212 16192 4218 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 9306 16192 9312 16244
rect 9364 16192 9370 16244
rect 12802 16192 12808 16244
rect 12860 16192 12866 16244
rect 13262 16192 13268 16244
rect 13320 16192 13326 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 13872 16204 14289 16232
rect 13872 16192 13878 16204
rect 14277 16201 14289 16204
rect 14323 16232 14335 16235
rect 14918 16232 14924 16244
rect 14323 16204 14924 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 15102 16192 15108 16244
rect 15160 16192 15166 16244
rect 15473 16235 15531 16241
rect 15473 16201 15485 16235
rect 15519 16232 15531 16235
rect 15746 16232 15752 16244
rect 15519 16204 15752 16232
rect 15519 16201 15531 16204
rect 15473 16195 15531 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 16114 16192 16120 16244
rect 16172 16192 16178 16244
rect 17310 16192 17316 16244
rect 17368 16192 17374 16244
rect 19061 16235 19119 16241
rect 19061 16201 19073 16235
rect 19107 16232 19119 16235
rect 19150 16232 19156 16244
rect 19107 16204 19156 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 19521 16235 19579 16241
rect 19521 16201 19533 16235
rect 19567 16232 19579 16235
rect 19610 16232 19616 16244
rect 19567 16204 19616 16232
rect 19567 16201 19579 16204
rect 19521 16195 19579 16201
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 20622 16232 20628 16244
rect 19720 16204 20628 16232
rect 2354 16136 2774 16164
rect 7500 16167 7558 16173
rect 2354 16133 2366 16136
rect 2308 16127 2366 16133
rect 7500 16133 7512 16167
rect 7546 16164 7558 16167
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 7546 16136 7849 16164
rect 7546 16133 7558 16136
rect 7500 16127 7558 16133
rect 7837 16133 7849 16136
rect 7883 16133 7895 16167
rect 7837 16127 7895 16133
rect 9208 16167 9266 16173
rect 9208 16133 9220 16167
rect 9254 16164 9266 16167
rect 9324 16164 9352 16192
rect 9254 16136 9352 16164
rect 13280 16164 13308 16192
rect 15565 16167 15623 16173
rect 13280 16136 13676 16164
rect 9254 16133 9266 16136
rect 9208 16127 9266 16133
rect 4154 16056 4160 16108
rect 4212 16096 4218 16108
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 4212 16068 4537 16096
rect 4212 16056 4218 16068
rect 4525 16065 4537 16068
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8941 16099 8999 16105
rect 8941 16096 8953 16099
rect 7800 16068 8953 16096
rect 7800 16056 7806 16068
rect 8941 16065 8953 16068
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13446 16056 13452 16108
rect 13504 16056 13510 16108
rect 13648 16105 13676 16136
rect 15565 16133 15577 16167
rect 15611 16164 15623 16167
rect 16132 16164 16160 16192
rect 17328 16164 17356 16192
rect 15611 16136 16160 16164
rect 17052 16136 17356 16164
rect 15611 16133 15623 16136
rect 15565 16127 15623 16133
rect 17052 16105 17080 16136
rect 18414 16124 18420 16176
rect 18472 16164 18478 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18472 16136 19441 16164
rect 18472 16124 18478 16136
rect 19429 16133 19441 16136
rect 19475 16164 19487 16167
rect 19720 16164 19748 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 21269 16235 21327 16241
rect 21269 16201 21281 16235
rect 21315 16232 21327 16235
rect 21634 16232 21640 16244
rect 21315 16204 21640 16232
rect 21315 16201 21327 16204
rect 21269 16195 21327 16201
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16232 21879 16235
rect 22094 16232 22100 16244
rect 21867 16204 22100 16232
rect 21867 16201 21879 16204
rect 21821 16195 21879 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22186 16192 22192 16244
rect 22244 16192 22250 16244
rect 23382 16192 23388 16244
rect 23440 16192 23446 16244
rect 24213 16235 24271 16241
rect 24213 16201 24225 16235
rect 24259 16232 24271 16235
rect 24394 16232 24400 16244
rect 24259 16204 24400 16232
rect 24259 16201 24271 16204
rect 24213 16195 24271 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 25314 16232 25320 16244
rect 24504 16204 25320 16232
rect 19475 16136 19748 16164
rect 20156 16167 20214 16173
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 20156 16133 20168 16167
rect 20202 16164 20214 16167
rect 20346 16164 20352 16176
rect 20202 16136 20352 16164
rect 20202 16133 20214 16136
rect 20156 16127 20214 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 23100 16167 23158 16173
rect 23100 16133 23112 16167
rect 23146 16164 23158 16167
rect 23400 16164 23428 16192
rect 23146 16136 23428 16164
rect 23146 16133 23158 16136
rect 23100 16127 23158 16133
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17304 16099 17362 16105
rect 17304 16065 17316 16099
rect 17350 16096 17362 16099
rect 17586 16096 17592 16108
rect 17350 16068 17592 16096
rect 17350 16065 17362 16068
rect 17304 16059 17362 16065
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19576 16068 19901 16096
rect 19576 16056 19582 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 21637 16099 21695 16105
rect 21637 16065 21649 16099
rect 21683 16096 21695 16099
rect 24504 16096 24532 16204
rect 25314 16192 25320 16204
rect 25372 16232 25378 16244
rect 26786 16232 26792 16244
rect 25372 16204 26792 16232
rect 25372 16192 25378 16204
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 27246 16192 27252 16244
rect 27304 16192 27310 16244
rect 28537 16235 28595 16241
rect 28537 16201 28549 16235
rect 28583 16232 28595 16235
rect 28810 16232 28816 16244
rect 28583 16204 28816 16232
rect 28583 16201 28595 16204
rect 28537 16195 28595 16201
rect 28810 16192 28816 16204
rect 28868 16192 28874 16244
rect 29546 16192 29552 16244
rect 29604 16192 29610 16244
rect 31389 16235 31447 16241
rect 31389 16201 31401 16235
rect 31435 16232 31447 16235
rect 31570 16232 31576 16244
rect 31435 16204 31576 16232
rect 31435 16201 31447 16204
rect 31389 16195 31447 16201
rect 31570 16192 31576 16204
rect 31628 16192 31634 16244
rect 32030 16192 32036 16244
rect 32088 16232 32094 16244
rect 32769 16235 32827 16241
rect 32769 16232 32781 16235
rect 32088 16204 32781 16232
rect 32088 16192 32094 16204
rect 32769 16201 32781 16204
rect 32815 16201 32827 16235
rect 32769 16195 32827 16201
rect 37642 16192 37648 16244
rect 37700 16192 37706 16244
rect 38657 16235 38715 16241
rect 38657 16201 38669 16235
rect 38703 16232 38715 16235
rect 38746 16232 38752 16244
rect 38703 16204 38752 16232
rect 38703 16201 38715 16204
rect 38657 16195 38715 16201
rect 38746 16192 38752 16204
rect 38804 16192 38810 16244
rect 40497 16235 40555 16241
rect 40497 16201 40509 16235
rect 40543 16232 40555 16235
rect 41506 16232 41512 16244
rect 40543 16204 41512 16232
rect 40543 16201 40555 16204
rect 40497 16195 40555 16201
rect 41506 16192 41512 16204
rect 41564 16192 41570 16244
rect 41598 16192 41604 16244
rect 41656 16192 41662 16244
rect 47762 16232 47768 16244
rect 43640 16204 47768 16232
rect 27341 16167 27399 16173
rect 27341 16164 27353 16167
rect 26160 16136 27353 16164
rect 21683 16068 24532 16096
rect 21683 16065 21695 16068
rect 21637 16059 21695 16065
rect 2038 15988 2044 16040
rect 2096 15988 2102 16040
rect 4338 15988 4344 16040
rect 4396 15988 4402 16040
rect 4614 15988 4620 16040
rect 4672 15988 4678 16040
rect 5074 15988 5080 16040
rect 5132 15988 5138 16040
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 4632 15960 4660 15988
rect 3467 15932 4660 15960
rect 6196 15960 6224 15991
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 7892 16000 8401 16028
rect 7892 15988 7898 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 13188 16028 13216 16056
rect 14458 16028 14464 16040
rect 13188 16000 14464 16028
rect 8389 15991 8447 15997
rect 14458 15988 14464 16000
rect 14516 16028 14522 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14516 16000 14933 16028
rect 14516 15988 14522 16000
rect 14921 15997 14933 16000
rect 14967 16028 14979 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 14967 16000 15669 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 19610 15988 19616 16040
rect 19668 15988 19674 16040
rect 22278 15988 22284 16040
rect 22336 15988 22342 16040
rect 22480 16037 22508 16068
rect 25406 16056 25412 16108
rect 25464 16056 25470 16108
rect 26160 16105 26188 16136
rect 27341 16133 27353 16136
rect 27387 16164 27399 16167
rect 27801 16167 27859 16173
rect 27801 16164 27813 16167
rect 27387 16136 27813 16164
rect 27387 16133 27399 16136
rect 27341 16127 27399 16133
rect 27801 16133 27813 16136
rect 27847 16133 27859 16167
rect 29564 16164 29592 16192
rect 34548 16167 34606 16173
rect 29564 16136 29960 16164
rect 27801 16127 27859 16133
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 26326 16056 26332 16108
rect 26384 16056 26390 16108
rect 26694 16056 26700 16108
rect 26752 16056 26758 16108
rect 29362 16056 29368 16108
rect 29420 16096 29426 16108
rect 29932 16105 29960 16136
rect 34548 16133 34560 16167
rect 34594 16164 34606 16167
rect 34698 16164 34704 16176
rect 34594 16136 34704 16164
rect 34594 16133 34606 16136
rect 34548 16127 34606 16133
rect 34698 16124 34704 16136
rect 34756 16124 34762 16176
rect 29650 16099 29708 16105
rect 29650 16096 29662 16099
rect 29420 16068 29662 16096
rect 29420 16056 29426 16068
rect 29650 16065 29662 16068
rect 29696 16065 29708 16099
rect 29650 16059 29708 16065
rect 29917 16099 29975 16105
rect 29917 16065 29929 16099
rect 29963 16096 29975 16099
rect 30009 16099 30067 16105
rect 30009 16096 30021 16099
rect 29963 16068 30021 16096
rect 29963 16065 29975 16068
rect 29917 16059 29975 16065
rect 30009 16065 30021 16068
rect 30055 16065 30067 16099
rect 30009 16059 30067 16065
rect 30276 16099 30334 16105
rect 30276 16065 30288 16099
rect 30322 16096 30334 16099
rect 30834 16096 30840 16108
rect 30322 16068 30840 16096
rect 30322 16065 30334 16068
rect 30276 16059 30334 16065
rect 30834 16056 30840 16068
rect 30892 16056 30898 16108
rect 34793 16099 34851 16105
rect 34793 16065 34805 16099
rect 34839 16096 34851 16099
rect 35713 16099 35771 16105
rect 35713 16096 35725 16099
rect 34839 16068 35725 16096
rect 34839 16065 34851 16068
rect 34793 16059 34851 16065
rect 35713 16065 35725 16068
rect 35759 16096 35771 16099
rect 35802 16096 35808 16108
rect 35759 16068 35808 16096
rect 35759 16065 35771 16068
rect 35713 16059 35771 16065
rect 35802 16056 35808 16068
rect 35860 16056 35866 16108
rect 35980 16099 36038 16105
rect 35980 16065 35992 16099
rect 36026 16096 36038 16099
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 36026 16068 37289 16096
rect 36026 16065 36038 16068
rect 35980 16059 36038 16065
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37660 16096 37688 16192
rect 39384 16167 39442 16173
rect 39384 16133 39396 16167
rect 39430 16164 39442 16167
rect 40586 16164 40592 16176
rect 39430 16136 40592 16164
rect 39430 16133 39442 16136
rect 39384 16127 39442 16133
rect 40586 16124 40592 16136
rect 40644 16124 40650 16176
rect 42334 16124 42340 16176
rect 42392 16164 42398 16176
rect 42392 16136 43116 16164
rect 42392 16124 42398 16136
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37660 16068 37841 16096
rect 37277 16059 37335 16065
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 39117 16099 39175 16105
rect 39117 16065 39129 16099
rect 39163 16096 39175 16099
rect 39206 16096 39212 16108
rect 39163 16068 39212 16096
rect 39163 16065 39175 16068
rect 39117 16059 39175 16065
rect 39206 16056 39212 16068
rect 39264 16056 39270 16108
rect 42797 16099 42855 16105
rect 42797 16065 42809 16099
rect 42843 16096 42855 16099
rect 42978 16096 42984 16108
rect 42843 16068 42984 16096
rect 42843 16065 42855 16068
rect 42797 16059 42855 16065
rect 42978 16056 42984 16068
rect 43036 16056 43042 16108
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22612 16000 22845 16028
rect 22612 15988 22618 16000
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 24762 15988 24768 16040
rect 24820 16028 24826 16040
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24820 16000 25145 16028
rect 24820 15988 24826 16000
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 25222 15988 25228 16040
rect 25280 16037 25286 16040
rect 25280 16031 25329 16037
rect 25280 15997 25283 16031
rect 25317 15997 25329 16031
rect 26712 16028 26740 16056
rect 27065 16031 27123 16037
rect 27065 16028 27077 16031
rect 26712 16000 27077 16028
rect 25280 15991 25329 15997
rect 27065 15997 27077 16000
rect 27111 15997 27123 16031
rect 27065 15991 27123 15997
rect 25280 15988 25286 15991
rect 27614 15988 27620 16040
rect 27672 16028 27678 16040
rect 43088 16037 43116 16136
rect 28353 16031 28411 16037
rect 28353 16028 28365 16031
rect 27672 16000 28365 16028
rect 27672 15988 27678 16000
rect 28353 15997 28365 16000
rect 28399 15997 28411 16031
rect 38013 16031 38071 16037
rect 38013 16028 38025 16031
rect 28353 15991 28411 15997
rect 37108 16000 38025 16028
rect 6365 15963 6423 15969
rect 6365 15960 6377 15963
rect 6196 15932 6377 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 6365 15929 6377 15932
rect 6411 15929 6423 15963
rect 6365 15923 6423 15929
rect 25682 15920 25688 15972
rect 25740 15920 25746 15972
rect 37108 15969 37136 16000
rect 38013 15997 38025 16000
rect 38059 15997 38071 16031
rect 38013 15991 38071 15997
rect 42245 16031 42303 16037
rect 42245 15997 42257 16031
rect 42291 15997 42303 16031
rect 42889 16031 42947 16037
rect 42889 16028 42901 16031
rect 42245 15991 42303 15997
rect 42812 16000 42901 16028
rect 37093 15963 37151 15969
rect 37093 15929 37105 15963
rect 37139 15929 37151 15963
rect 42260 15960 42288 15991
rect 42429 15963 42487 15969
rect 42429 15960 42441 15963
rect 42260 15932 42441 15960
rect 37093 15923 37151 15929
rect 42429 15929 42441 15932
rect 42475 15929 42487 15963
rect 42429 15923 42487 15929
rect 42812 15904 42840 16000
rect 42889 15997 42901 16000
rect 42935 15997 42947 16031
rect 42889 15991 42947 15997
rect 43073 16031 43131 16037
rect 43073 15997 43085 16031
rect 43119 16028 43131 16031
rect 43640 16028 43668 16204
rect 47762 16192 47768 16204
rect 47820 16192 47826 16244
rect 48682 16192 48688 16244
rect 48740 16192 48746 16244
rect 49605 16235 49663 16241
rect 49605 16201 49617 16235
rect 49651 16232 49663 16235
rect 50338 16232 50344 16244
rect 49651 16204 50344 16232
rect 49651 16201 49663 16204
rect 49605 16195 49663 16201
rect 50338 16192 50344 16204
rect 50396 16192 50402 16244
rect 51258 16192 51264 16244
rect 51316 16232 51322 16244
rect 52273 16235 52331 16241
rect 52273 16232 52285 16235
rect 51316 16204 52285 16232
rect 51316 16192 51322 16204
rect 52273 16201 52285 16204
rect 52319 16201 52331 16235
rect 52273 16195 52331 16201
rect 54297 16235 54355 16241
rect 54297 16201 54309 16235
rect 54343 16232 54355 16235
rect 55401 16235 55459 16241
rect 55401 16232 55413 16235
rect 54343 16204 55413 16232
rect 54343 16201 54355 16204
rect 54297 16195 54355 16201
rect 55401 16201 55413 16204
rect 55447 16232 55459 16235
rect 56318 16232 56324 16244
rect 55447 16204 56324 16232
rect 55447 16201 55459 16204
rect 55401 16195 55459 16201
rect 56318 16192 56324 16204
rect 56376 16192 56382 16244
rect 57146 16192 57152 16244
rect 57204 16192 57210 16244
rect 57514 16192 57520 16244
rect 57572 16192 57578 16244
rect 44266 16056 44272 16108
rect 44324 16105 44330 16108
rect 44324 16099 44373 16105
rect 44324 16065 44327 16099
rect 44361 16065 44373 16099
rect 44324 16059 44373 16065
rect 44324 16056 44330 16059
rect 45278 16056 45284 16108
rect 45336 16096 45342 16108
rect 45373 16099 45431 16105
rect 45373 16096 45385 16099
rect 45336 16068 45385 16096
rect 45336 16056 45342 16068
rect 45373 16065 45385 16068
rect 45419 16065 45431 16099
rect 45373 16059 45431 16065
rect 45554 16056 45560 16108
rect 45612 16056 45618 16108
rect 47210 16056 47216 16108
rect 47268 16096 47274 16108
rect 48133 16099 48191 16105
rect 48133 16096 48145 16099
rect 47268 16068 48145 16096
rect 47268 16056 47274 16068
rect 48133 16065 48145 16068
rect 48179 16065 48191 16099
rect 48700 16096 48728 16192
rect 54754 16124 54760 16176
rect 54812 16164 54818 16176
rect 54812 16136 54892 16164
rect 54812 16124 54818 16136
rect 48961 16099 49019 16105
rect 48961 16096 48973 16099
rect 48700 16068 48973 16096
rect 48133 16059 48191 16065
rect 48961 16065 48973 16068
rect 49007 16065 49019 16099
rect 48961 16059 49019 16065
rect 49694 16056 49700 16108
rect 49752 16056 49758 16108
rect 51994 16056 52000 16108
rect 52052 16056 52058 16108
rect 54864 16105 54892 16136
rect 54849 16099 54907 16105
rect 54849 16065 54861 16099
rect 54895 16065 54907 16099
rect 54849 16059 54907 16065
rect 56781 16099 56839 16105
rect 56781 16065 56793 16099
rect 56827 16096 56839 16099
rect 56870 16096 56876 16108
rect 56827 16068 56876 16096
rect 56827 16065 56839 16068
rect 56781 16059 56839 16065
rect 56870 16056 56876 16068
rect 56928 16056 56934 16108
rect 57532 16096 57560 16192
rect 58437 16099 58495 16105
rect 58437 16096 58449 16099
rect 57532 16068 58449 16096
rect 58437 16065 58449 16068
rect 58483 16065 58495 16099
rect 58437 16059 58495 16065
rect 43119 16000 43668 16028
rect 43119 15997 43131 16000
rect 43073 15991 43131 15997
rect 44174 15988 44180 16040
rect 44232 15988 44238 16040
rect 44453 16031 44511 16037
rect 44453 15997 44465 16031
rect 44499 16028 44511 16031
rect 44634 16028 44640 16040
rect 44499 16000 44640 16028
rect 44499 15997 44511 16000
rect 44453 15991 44511 15997
rect 44634 15988 44640 16000
rect 44692 15988 44698 16040
rect 45189 16031 45247 16037
rect 45189 15997 45201 16031
rect 45235 16028 45247 16031
rect 45572 16028 45600 16056
rect 45235 16000 45600 16028
rect 45235 15997 45247 16000
rect 45189 15991 45247 15997
rect 49510 15988 49516 16040
rect 49568 15988 49574 16040
rect 50614 15988 50620 16040
rect 50672 16028 50678 16040
rect 50985 16031 51043 16037
rect 50985 16028 50997 16031
rect 50672 16000 50997 16028
rect 50672 15988 50678 16000
rect 50985 15997 50997 16000
rect 51031 15997 51043 16031
rect 54021 16031 54079 16037
rect 54021 16028 54033 16031
rect 50985 15991 51043 15997
rect 53760 16000 54033 16028
rect 44729 15963 44787 15969
rect 44729 15929 44741 15963
rect 44775 15960 44787 15963
rect 44818 15960 44824 15972
rect 44775 15932 44824 15960
rect 44775 15929 44787 15932
rect 44729 15923 44787 15929
rect 44818 15920 44824 15932
rect 44876 15960 44882 15972
rect 46382 15960 46388 15972
rect 44876 15932 46388 15960
rect 44876 15920 44882 15932
rect 46382 15920 46388 15932
rect 46440 15960 46446 15972
rect 49528 15960 49556 15988
rect 53760 15969 53788 16000
rect 54021 15997 54033 16000
rect 54067 15997 54079 16031
rect 54021 15991 54079 15997
rect 54202 15988 54208 16040
rect 54260 15988 54266 16040
rect 55858 16028 55864 16040
rect 54680 16000 55864 16028
rect 54680 15969 54708 16000
rect 55858 15988 55864 16000
rect 55916 15988 55922 16040
rect 56505 16031 56563 16037
rect 56505 16028 56517 16031
rect 56244 16000 56517 16028
rect 53745 15963 53803 15969
rect 53745 15960 53757 15963
rect 46440 15932 49556 15960
rect 50264 15932 53757 15960
rect 46440 15920 46446 15932
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 4120 15864 5549 15892
rect 4120 15852 4126 15864
rect 5537 15861 5549 15864
rect 5583 15892 5595 15895
rect 6546 15892 6552 15904
rect 5583 15864 6552 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 10321 15895 10379 15901
rect 10321 15861 10333 15895
rect 10367 15892 10379 15895
rect 10686 15892 10692 15904
rect 10367 15864 10692 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 14645 15895 14703 15901
rect 14645 15861 14657 15895
rect 14691 15892 14703 15895
rect 14918 15892 14924 15904
rect 14691 15864 14924 15892
rect 14691 15861 14703 15864
rect 14645 15855 14703 15861
rect 14918 15852 14924 15864
rect 14976 15892 14982 15904
rect 15286 15892 15292 15904
rect 14976 15864 15292 15892
rect 14976 15852 14982 15864
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 18414 15852 18420 15904
rect 18472 15852 18478 15904
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 19886 15892 19892 15904
rect 19024 15864 19892 15892
rect 19024 15852 19030 15864
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 24489 15895 24547 15901
rect 24489 15861 24501 15895
rect 24535 15892 24547 15895
rect 25958 15892 25964 15904
rect 24535 15864 25964 15892
rect 24535 15861 24547 15864
rect 24489 15855 24547 15861
rect 25958 15852 25964 15864
rect 26016 15852 26022 15904
rect 27706 15852 27712 15904
rect 27764 15852 27770 15904
rect 33134 15852 33140 15904
rect 33192 15852 33198 15904
rect 33413 15895 33471 15901
rect 33413 15861 33425 15895
rect 33459 15892 33471 15895
rect 34514 15892 34520 15904
rect 33459 15864 34520 15892
rect 33459 15861 33471 15864
rect 33413 15855 33471 15861
rect 34514 15852 34520 15864
rect 34572 15852 34578 15904
rect 42794 15852 42800 15904
rect 42852 15852 42858 15904
rect 43533 15895 43591 15901
rect 43533 15861 43545 15895
rect 43579 15892 43591 15895
rect 45278 15892 45284 15904
rect 43579 15864 45284 15892
rect 43579 15861 43591 15864
rect 43533 15855 43591 15861
rect 45278 15852 45284 15864
rect 45336 15852 45342 15904
rect 47118 15852 47124 15904
rect 47176 15892 47182 15904
rect 47581 15895 47639 15901
rect 47581 15892 47593 15895
rect 47176 15864 47593 15892
rect 47176 15852 47182 15864
rect 47581 15861 47593 15864
rect 47627 15861 47639 15895
rect 47581 15855 47639 15861
rect 48590 15852 48596 15904
rect 48648 15892 48654 15904
rect 50264 15892 50292 15932
rect 53745 15929 53757 15932
rect 53791 15929 53803 15963
rect 53745 15923 53803 15929
rect 54665 15963 54723 15969
rect 54665 15929 54677 15963
rect 54711 15929 54723 15963
rect 54665 15923 54723 15929
rect 48648 15864 50292 15892
rect 48648 15852 48654 15864
rect 50338 15852 50344 15904
rect 50396 15852 50402 15904
rect 50430 15852 50436 15904
rect 50488 15852 50494 15904
rect 51350 15852 51356 15904
rect 51408 15852 51414 15904
rect 55674 15852 55680 15904
rect 55732 15892 55738 15904
rect 56244 15901 56272 16000
rect 56505 15997 56517 16000
rect 56551 15997 56563 16031
rect 56505 15991 56563 15997
rect 56689 16031 56747 16037
rect 56689 15997 56701 16031
rect 56735 16028 56747 16031
rect 57054 16028 57060 16040
rect 56735 16000 57060 16028
rect 56735 15997 56747 16000
rect 56689 15991 56747 15997
rect 57054 15988 57060 16000
rect 57112 16028 57118 16040
rect 57885 16031 57943 16037
rect 57885 16028 57897 16031
rect 57112 16000 57897 16028
rect 57112 15988 57118 16000
rect 57885 15997 57897 16000
rect 57931 15997 57943 16031
rect 57885 15991 57943 15997
rect 56229 15895 56287 15901
rect 56229 15892 56241 15895
rect 55732 15864 56241 15892
rect 55732 15852 55738 15864
rect 56229 15861 56241 15864
rect 56275 15861 56287 15895
rect 56229 15855 56287 15861
rect 1104 15802 58880 15824
rect 1104 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 22616 15802
rect 22668 15750 22680 15802
rect 22732 15750 22744 15802
rect 22796 15750 22808 15802
rect 22860 15750 22872 15802
rect 22924 15750 37060 15802
rect 37112 15750 37124 15802
rect 37176 15750 37188 15802
rect 37240 15750 37252 15802
rect 37304 15750 37316 15802
rect 37368 15750 51504 15802
rect 51556 15750 51568 15802
rect 51620 15750 51632 15802
rect 51684 15750 51696 15802
rect 51748 15750 51760 15802
rect 51812 15750 58880 15802
rect 1104 15728 58880 15750
rect 4154 15688 4160 15700
rect 3896 15660 4160 15688
rect 3896 15561 3924 15660
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 6917 15691 6975 15697
rect 4540 15660 6132 15688
rect 4540 15629 4568 15660
rect 4525 15623 4583 15629
rect 4525 15589 4537 15623
rect 4571 15589 4583 15623
rect 4525 15583 4583 15589
rect 6104 15564 6132 15660
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 7834 15688 7840 15700
rect 6963 15660 7840 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 54018 15688 54024 15700
rect 8536 15660 54024 15688
rect 8536 15648 8542 15660
rect 54018 15648 54024 15660
rect 54076 15648 54082 15700
rect 6454 15620 6460 15632
rect 6380 15592 6460 15620
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 4062 15512 4068 15564
rect 4120 15512 4126 15564
rect 4890 15512 4896 15564
rect 4948 15561 4954 15564
rect 4948 15555 4976 15561
rect 4964 15521 4976 15555
rect 4948 15515 4976 15521
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15552 5135 15555
rect 5258 15552 5264 15564
rect 5123 15524 5264 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 4948 15512 4954 15515
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 6086 15512 6092 15564
rect 6144 15512 6150 15564
rect 6380 15561 6408 15592
rect 6454 15580 6460 15592
rect 6512 15620 6518 15632
rect 6730 15620 6736 15632
rect 6512 15592 6736 15620
rect 6512 15580 6518 15592
rect 6730 15580 6736 15592
rect 6788 15620 6794 15632
rect 10137 15623 10195 15629
rect 6788 15592 8248 15620
rect 6788 15580 6794 15592
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15521 6423 15555
rect 7006 15552 7012 15564
rect 6365 15515 6423 15521
rect 6472 15524 7012 15552
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2682 15484 2688 15496
rect 2096 15456 2688 15484
rect 2096 15444 2102 15456
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 4798 15444 4804 15496
rect 4856 15444 4862 15496
rect 6472 15493 6500 15524
rect 7006 15512 7012 15524
rect 7064 15552 7070 15564
rect 7064 15524 7420 15552
rect 7064 15512 7070 15524
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 5644 15456 6469 15484
rect 2130 15376 2136 15428
rect 2188 15416 2194 15428
rect 2286 15419 2344 15425
rect 2286 15416 2298 15419
rect 2188 15388 2298 15416
rect 2188 15376 2194 15388
rect 2286 15385 2298 15388
rect 2332 15385 2344 15419
rect 2286 15379 2344 15385
rect 3421 15351 3479 15357
rect 3421 15317 3433 15351
rect 3467 15348 3479 15351
rect 4338 15348 4344 15360
rect 3467 15320 4344 15348
rect 3467 15317 3479 15320
rect 3421 15311 3479 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 5644 15348 5672 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 7392 15493 7420 15524
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8220 15552 8248 15592
rect 10137 15589 10149 15623
rect 10183 15620 10195 15623
rect 10410 15620 10416 15632
rect 10183 15592 10416 15620
rect 10183 15589 10195 15592
rect 10137 15583 10195 15589
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 13170 15620 13176 15632
rect 12406 15592 13176 15620
rect 12406 15552 12434 15592
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 24121 15623 24179 15629
rect 24121 15589 24133 15623
rect 24167 15620 24179 15623
rect 27433 15623 27491 15629
rect 24167 15592 24440 15620
rect 24167 15589 24179 15592
rect 24121 15583 24179 15589
rect 7708 15524 8156 15552
rect 8220 15524 12434 15552
rect 7708 15512 7714 15524
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 5721 15419 5779 15425
rect 5721 15385 5733 15419
rect 5767 15416 5779 15419
rect 7098 15416 7104 15428
rect 5767 15388 7104 15416
rect 5767 15385 5779 15388
rect 5721 15379 5779 15385
rect 7098 15376 7104 15388
rect 7156 15376 7162 15428
rect 7190 15376 7196 15428
rect 7248 15376 7254 15428
rect 4488 15320 5672 15348
rect 4488 15308 4494 15320
rect 6086 15308 6092 15360
rect 6144 15348 6150 15360
rect 6914 15348 6920 15360
rect 6144 15320 6920 15348
rect 6144 15308 6150 15320
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7009 15351 7067 15357
rect 7009 15317 7021 15351
rect 7055 15348 7067 15351
rect 7208 15348 7236 15376
rect 8128 15360 8156 15524
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16724 15524 16773 15552
rect 16724 15512 16730 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 16761 15515 16819 15521
rect 18417 15555 18475 15561
rect 18417 15521 18429 15555
rect 18463 15552 18475 15555
rect 18506 15552 18512 15564
rect 18463 15524 18512 15552
rect 18463 15521 18475 15524
rect 18417 15515 18475 15521
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 24412 15561 24440 15592
rect 27433 15589 27445 15623
rect 27479 15620 27491 15623
rect 27614 15620 27620 15632
rect 27479 15592 27620 15620
rect 27479 15589 27491 15592
rect 27433 15583 27491 15589
rect 27614 15580 27620 15592
rect 27672 15580 27678 15632
rect 27706 15580 27712 15632
rect 27764 15580 27770 15632
rect 30101 15623 30159 15629
rect 30101 15589 30113 15623
rect 30147 15620 30159 15623
rect 30374 15620 30380 15632
rect 30147 15592 30380 15620
rect 30147 15589 30159 15592
rect 30101 15583 30159 15589
rect 30374 15580 30380 15592
rect 30432 15580 30438 15632
rect 30742 15580 30748 15632
rect 30800 15580 30806 15632
rect 30834 15580 30840 15632
rect 30892 15620 30898 15632
rect 30929 15623 30987 15629
rect 30929 15620 30941 15623
rect 30892 15592 30941 15620
rect 30892 15580 30898 15592
rect 30929 15589 30941 15592
rect 30975 15589 30987 15623
rect 31938 15620 31944 15632
rect 30929 15583 30987 15589
rect 31726 15592 31944 15620
rect 22741 15555 22799 15561
rect 22741 15552 22753 15555
rect 22520 15524 22753 15552
rect 22520 15512 22526 15524
rect 22741 15521 22753 15524
rect 22787 15521 22799 15555
rect 22741 15515 22799 15521
rect 24397 15555 24455 15561
rect 24397 15521 24409 15555
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 26053 15555 26111 15561
rect 26053 15552 26065 15555
rect 24912 15524 26065 15552
rect 24912 15512 24918 15524
rect 26053 15521 26065 15524
rect 26099 15521 26111 15555
rect 27724 15552 27752 15580
rect 28077 15555 28135 15561
rect 28077 15552 28089 15555
rect 27724 15524 28089 15552
rect 26053 15515 26111 15521
rect 28077 15521 28089 15524
rect 28123 15521 28135 15555
rect 28077 15515 28135 15521
rect 28718 15512 28724 15564
rect 28776 15512 28782 15564
rect 30653 15555 30711 15561
rect 30653 15521 30665 15555
rect 30699 15521 30711 15555
rect 30760 15552 30788 15580
rect 31481 15555 31539 15561
rect 31481 15552 31493 15555
rect 30760 15524 31493 15552
rect 30653 15515 30711 15521
rect 31481 15521 31493 15524
rect 31527 15521 31539 15555
rect 31481 15515 31539 15521
rect 9674 15444 9680 15496
rect 9732 15444 9738 15496
rect 12526 15444 12532 15496
rect 12584 15444 12590 15496
rect 12894 15444 12900 15496
rect 12952 15444 12958 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15484 18199 15487
rect 19058 15484 19064 15496
rect 18187 15456 19064 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 30466 15444 30472 15496
rect 30524 15444 30530 15496
rect 30668 15484 30696 15515
rect 30742 15484 30748 15496
rect 30668 15456 30748 15484
rect 30742 15444 30748 15456
rect 30800 15484 30806 15496
rect 31726 15484 31754 15592
rect 31938 15580 31944 15592
rect 31996 15580 32002 15632
rect 42334 15580 42340 15632
rect 42392 15580 42398 15632
rect 43165 15623 43223 15629
rect 43165 15589 43177 15623
rect 43211 15589 43223 15623
rect 43165 15583 43223 15589
rect 41969 15555 42027 15561
rect 41969 15521 41981 15555
rect 42015 15552 42027 15555
rect 42150 15552 42156 15564
rect 42015 15524 42156 15552
rect 42015 15521 42027 15524
rect 41969 15515 42027 15521
rect 42150 15512 42156 15524
rect 42208 15552 42214 15564
rect 42610 15552 42616 15564
rect 42208 15524 42616 15552
rect 42208 15512 42214 15524
rect 42610 15512 42616 15524
rect 42668 15512 42674 15564
rect 43180 15552 43208 15583
rect 43254 15580 43260 15632
rect 43312 15580 43318 15632
rect 44269 15623 44327 15629
rect 44269 15589 44281 15623
rect 44315 15620 44327 15623
rect 44818 15620 44824 15632
rect 44315 15592 44824 15620
rect 44315 15589 44327 15592
rect 44269 15583 44327 15589
rect 44818 15580 44824 15592
rect 44876 15580 44882 15632
rect 48130 15620 48136 15632
rect 47688 15592 48136 15620
rect 43809 15555 43867 15561
rect 43809 15552 43821 15555
rect 43180 15524 43821 15552
rect 43809 15521 43821 15524
rect 43855 15521 43867 15555
rect 43809 15515 43867 15521
rect 44174 15512 44180 15564
rect 44232 15552 44238 15564
rect 44545 15555 44603 15561
rect 44545 15552 44557 15555
rect 44232 15524 44557 15552
rect 44232 15512 44238 15524
rect 44545 15521 44557 15524
rect 44591 15552 44603 15555
rect 47578 15552 47584 15564
rect 44591 15524 47584 15552
rect 44591 15521 44603 15524
rect 44545 15515 44603 15521
rect 47578 15512 47584 15524
rect 47636 15552 47642 15564
rect 47688 15552 47716 15592
rect 48130 15580 48136 15592
rect 48188 15580 48194 15632
rect 48593 15623 48651 15629
rect 48593 15589 48605 15623
rect 48639 15620 48651 15623
rect 52365 15623 52423 15629
rect 48639 15592 49280 15620
rect 48639 15589 48651 15592
rect 48593 15583 48651 15589
rect 47636 15524 47716 15552
rect 47765 15555 47823 15561
rect 47636 15512 47642 15524
rect 47765 15521 47777 15555
rect 47811 15552 47823 15555
rect 48038 15552 48044 15564
rect 47811 15524 48044 15552
rect 47811 15521 47823 15524
rect 47765 15515 47823 15521
rect 48038 15512 48044 15524
rect 48096 15512 48102 15564
rect 49252 15561 49280 15592
rect 50080 15592 52316 15620
rect 49237 15555 49295 15561
rect 49237 15521 49249 15555
rect 49283 15521 49295 15555
rect 49237 15515 49295 15521
rect 30800 15456 31754 15484
rect 37553 15487 37611 15493
rect 30800 15444 30806 15456
rect 37553 15453 37565 15487
rect 37599 15484 37611 15487
rect 37826 15484 37832 15496
rect 37599 15456 37832 15484
rect 37599 15453 37611 15456
rect 37553 15447 37611 15453
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 18233 15419 18291 15425
rect 18233 15385 18245 15419
rect 18279 15416 18291 15419
rect 18322 15416 18328 15428
rect 18279 15388 18328 15416
rect 18279 15385 18291 15388
rect 18233 15379 18291 15385
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 20438 15416 20444 15428
rect 19168 15388 20444 15416
rect 19168 15360 19196 15388
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 23008 15419 23066 15425
rect 23008 15385 23020 15419
rect 23054 15416 23066 15419
rect 23198 15416 23204 15428
rect 23054 15388 23204 15416
rect 23054 15385 23066 15388
rect 23008 15379 23066 15385
rect 23198 15376 23204 15388
rect 23256 15376 23262 15428
rect 26320 15419 26378 15425
rect 26320 15385 26332 15419
rect 26366 15416 26378 15419
rect 27525 15419 27583 15425
rect 27525 15416 27537 15419
rect 26366 15388 27537 15416
rect 26366 15385 26378 15388
rect 26320 15379 26378 15385
rect 27525 15385 27537 15388
rect 27571 15385 27583 15419
rect 27525 15379 27583 15385
rect 30561 15419 30619 15425
rect 30561 15385 30573 15419
rect 30607 15416 30619 15419
rect 31202 15416 31208 15428
rect 30607 15388 31208 15416
rect 30607 15385 30619 15388
rect 30561 15379 30619 15385
rect 31202 15376 31208 15388
rect 31260 15376 31266 15428
rect 42628 15416 42656 15512
rect 42797 15487 42855 15493
rect 42797 15453 42809 15487
rect 42843 15484 42855 15487
rect 44634 15484 44640 15496
rect 42843 15456 44640 15484
rect 42843 15453 42855 15456
rect 42797 15447 42855 15453
rect 44634 15444 44640 15456
rect 44692 15444 44698 15496
rect 48222 15444 48228 15496
rect 48280 15444 48286 15496
rect 50080 15428 50108 15592
rect 50985 15555 51043 15561
rect 50985 15521 50997 15555
rect 51031 15552 51043 15555
rect 51031 15524 51212 15552
rect 51031 15521 51043 15524
rect 50985 15515 51043 15521
rect 50246 15444 50252 15496
rect 50304 15484 50310 15496
rect 51077 15487 51135 15493
rect 51077 15484 51089 15487
rect 50304 15456 51089 15484
rect 50304 15444 50310 15456
rect 51077 15453 51089 15456
rect 51123 15453 51135 15487
rect 51077 15447 51135 15453
rect 48133 15419 48191 15425
rect 42628 15388 48084 15416
rect 7055 15320 7236 15348
rect 7055 15317 7067 15320
rect 7009 15311 7067 15317
rect 7466 15308 7472 15360
rect 7524 15308 7530 15360
rect 8110 15308 8116 15360
rect 8168 15308 8174 15360
rect 9122 15308 9128 15360
rect 9180 15308 9186 15360
rect 11974 15308 11980 15360
rect 12032 15308 12038 15360
rect 13446 15308 13452 15360
rect 13504 15308 13510 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 15105 15351 15163 15357
rect 15105 15348 15117 15351
rect 15068 15320 15117 15348
rect 15068 15308 15074 15320
rect 15105 15317 15117 15320
rect 15151 15317 15163 15351
rect 15105 15311 15163 15317
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17405 15351 17463 15357
rect 17405 15348 17417 15351
rect 17276 15320 17417 15348
rect 17276 15308 17282 15320
rect 17405 15317 17417 15320
rect 17451 15317 17463 15351
rect 17405 15311 17463 15317
rect 17773 15351 17831 15357
rect 17773 15317 17785 15351
rect 17819 15348 17831 15351
rect 17954 15348 17960 15360
rect 17819 15320 17960 15348
rect 17819 15317 17831 15320
rect 17773 15311 17831 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18969 15351 19027 15357
rect 18969 15317 18981 15351
rect 19015 15348 19027 15351
rect 19150 15348 19156 15360
rect 19015 15320 19156 15348
rect 19015 15317 19027 15320
rect 18969 15311 19027 15317
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19610 15348 19616 15360
rect 19567 15320 19616 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19610 15308 19616 15320
rect 19668 15348 19674 15360
rect 20346 15348 20352 15360
rect 19668 15320 20352 15348
rect 19668 15308 19674 15320
rect 20346 15308 20352 15320
rect 20404 15348 20410 15360
rect 20898 15348 20904 15360
rect 20404 15320 20904 15348
rect 20404 15308 20410 15320
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 25038 15308 25044 15360
rect 25096 15308 25102 15360
rect 29270 15308 29276 15360
rect 29328 15348 29334 15360
rect 29365 15351 29423 15357
rect 29365 15348 29377 15351
rect 29328 15320 29377 15348
rect 29328 15308 29334 15320
rect 29365 15317 29377 15320
rect 29411 15317 29423 15351
rect 29365 15311 29423 15317
rect 37921 15351 37979 15357
rect 37921 15317 37933 15351
rect 37967 15348 37979 15351
rect 38286 15348 38292 15360
rect 37967 15320 38292 15348
rect 37967 15317 37979 15320
rect 37921 15311 37979 15317
rect 38286 15308 38292 15320
rect 38344 15308 38350 15360
rect 42705 15351 42763 15357
rect 42705 15317 42717 15351
rect 42751 15348 42763 15351
rect 42794 15348 42800 15360
rect 42751 15320 42800 15348
rect 42751 15317 42763 15320
rect 42705 15311 42763 15317
rect 42794 15308 42800 15320
rect 42852 15308 42858 15360
rect 48056 15348 48084 15388
rect 48133 15385 48145 15419
rect 48179 15416 48191 15419
rect 49602 15416 49608 15428
rect 48179 15388 49608 15416
rect 48179 15385 48191 15388
rect 48133 15379 48191 15385
rect 49602 15376 49608 15388
rect 49660 15376 49666 15428
rect 49697 15419 49755 15425
rect 49697 15385 49709 15419
rect 49743 15416 49755 15419
rect 50062 15416 50068 15428
rect 49743 15388 50068 15416
rect 49743 15385 49755 15388
rect 49697 15379 49755 15385
rect 50062 15376 50068 15388
rect 50120 15376 50126 15428
rect 51184 15416 51212 15524
rect 51258 15512 51264 15564
rect 51316 15552 51322 15564
rect 51721 15555 51779 15561
rect 51721 15552 51733 15555
rect 51316 15524 51733 15552
rect 51316 15512 51322 15524
rect 51721 15521 51733 15524
rect 51767 15552 51779 15555
rect 51902 15552 51908 15564
rect 51767 15524 51908 15552
rect 51767 15521 51779 15524
rect 51721 15515 51779 15521
rect 51902 15512 51908 15524
rect 51960 15512 51966 15564
rect 51997 15487 52055 15493
rect 51997 15453 52009 15487
rect 52043 15484 52055 15487
rect 52086 15484 52092 15496
rect 52043 15456 52092 15484
rect 52043 15453 52055 15456
rect 51997 15447 52055 15453
rect 52086 15444 52092 15456
rect 52144 15444 52150 15496
rect 52288 15484 52316 15592
rect 52365 15589 52377 15623
rect 52411 15620 52423 15623
rect 57241 15623 57299 15629
rect 52411 15592 53052 15620
rect 52411 15589 52423 15592
rect 52365 15583 52423 15589
rect 53024 15561 53052 15592
rect 57241 15589 57253 15623
rect 57287 15620 57299 15623
rect 57287 15592 57928 15620
rect 57287 15589 57299 15592
rect 57241 15583 57299 15589
rect 53009 15555 53067 15561
rect 53009 15521 53021 15555
rect 53055 15521 53067 15555
rect 56321 15555 56379 15561
rect 56321 15552 56333 15555
rect 53009 15515 53067 15521
rect 54036 15524 56333 15552
rect 53466 15484 53472 15496
rect 52288 15456 53472 15484
rect 53466 15444 53472 15456
rect 53524 15484 53530 15496
rect 54036 15484 54064 15524
rect 56321 15521 56333 15524
rect 56367 15552 56379 15555
rect 56597 15555 56655 15561
rect 56597 15552 56609 15555
rect 56367 15524 56609 15552
rect 56367 15521 56379 15524
rect 56321 15515 56379 15521
rect 56597 15521 56609 15524
rect 56643 15552 56655 15555
rect 57146 15552 57152 15564
rect 56643 15524 57152 15552
rect 56643 15521 56655 15524
rect 56597 15515 56655 15521
rect 57146 15512 57152 15524
rect 57204 15512 57210 15564
rect 57900 15561 57928 15592
rect 57885 15555 57943 15561
rect 57885 15521 57897 15555
rect 57931 15521 57943 15555
rect 57885 15515 57943 15521
rect 53524 15456 54064 15484
rect 53524 15444 53530 15456
rect 54110 15444 54116 15496
rect 54168 15444 54174 15496
rect 54846 15444 54852 15496
rect 54904 15444 54910 15496
rect 55214 15444 55220 15496
rect 55272 15484 55278 15496
rect 55309 15487 55367 15493
rect 55309 15484 55321 15487
rect 55272 15456 55321 15484
rect 55272 15444 55278 15456
rect 55309 15453 55321 15456
rect 55355 15453 55367 15487
rect 55309 15447 55367 15453
rect 55030 15416 55036 15428
rect 50632 15388 55036 15416
rect 48590 15348 48596 15360
rect 48056 15320 48596 15348
rect 48590 15308 48596 15320
rect 48648 15308 48654 15360
rect 48682 15308 48688 15360
rect 48740 15308 48746 15360
rect 49878 15308 49884 15360
rect 49936 15348 49942 15360
rect 50632 15357 50660 15388
rect 55030 15376 55036 15388
rect 55088 15376 55094 15428
rect 55122 15376 55128 15428
rect 55180 15416 55186 15428
rect 55180 15388 56916 15416
rect 55180 15376 55186 15388
rect 56888 15360 56916 15388
rect 50617 15351 50675 15357
rect 50617 15348 50629 15351
rect 49936 15320 50629 15348
rect 49936 15308 49942 15320
rect 50617 15317 50629 15320
rect 50663 15317 50675 15351
rect 50617 15311 50675 15317
rect 51169 15351 51227 15357
rect 51169 15317 51181 15351
rect 51215 15348 51227 15351
rect 51258 15348 51264 15360
rect 51215 15320 51264 15348
rect 51215 15317 51227 15320
rect 51169 15311 51227 15317
rect 51258 15308 51264 15320
rect 51316 15308 51322 15360
rect 51537 15351 51595 15357
rect 51537 15317 51549 15351
rect 51583 15348 51595 15351
rect 51810 15348 51816 15360
rect 51583 15320 51816 15348
rect 51583 15317 51595 15320
rect 51537 15311 51595 15317
rect 51810 15308 51816 15320
rect 51868 15308 51874 15360
rect 51905 15351 51963 15357
rect 51905 15317 51917 15351
rect 51951 15348 51963 15351
rect 52178 15348 52184 15360
rect 51951 15320 52184 15348
rect 51951 15317 51963 15320
rect 51905 15311 51963 15317
rect 52178 15308 52184 15320
rect 52236 15308 52242 15360
rect 52454 15308 52460 15360
rect 52512 15308 52518 15360
rect 53374 15308 53380 15360
rect 53432 15348 53438 15360
rect 53561 15351 53619 15357
rect 53561 15348 53573 15351
rect 53432 15320 53573 15348
rect 53432 15308 53438 15320
rect 53561 15317 53573 15320
rect 53607 15317 53619 15351
rect 53561 15311 53619 15317
rect 54294 15308 54300 15360
rect 54352 15308 54358 15360
rect 55953 15351 56011 15357
rect 55953 15317 55965 15351
rect 55999 15348 56011 15351
rect 56226 15348 56232 15360
rect 55999 15320 56232 15348
rect 55999 15317 56011 15320
rect 55953 15311 56011 15317
rect 56226 15308 56232 15320
rect 56284 15308 56290 15360
rect 56778 15308 56784 15360
rect 56836 15308 56842 15360
rect 56870 15308 56876 15360
rect 56928 15308 56934 15360
rect 57330 15308 57336 15360
rect 57388 15308 57394 15360
rect 1104 15258 59040 15280
rect 1104 15206 15394 15258
rect 15446 15206 15458 15258
rect 15510 15206 15522 15258
rect 15574 15206 15586 15258
rect 15638 15206 15650 15258
rect 15702 15206 29838 15258
rect 29890 15206 29902 15258
rect 29954 15206 29966 15258
rect 30018 15206 30030 15258
rect 30082 15206 30094 15258
rect 30146 15206 44282 15258
rect 44334 15206 44346 15258
rect 44398 15206 44410 15258
rect 44462 15206 44474 15258
rect 44526 15206 44538 15258
rect 44590 15206 58726 15258
rect 58778 15206 58790 15258
rect 58842 15206 58854 15258
rect 58906 15206 58918 15258
rect 58970 15206 58982 15258
rect 59034 15206 59040 15258
rect 1104 15184 59040 15206
rect 2130 15104 2136 15156
rect 2188 15104 2194 15156
rect 4249 15147 4307 15153
rect 4249 15113 4261 15147
rect 4295 15144 4307 15147
rect 5074 15144 5080 15156
rect 4295 15116 5080 15144
rect 4295 15113 4307 15116
rect 4249 15107 4307 15113
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 5350 15104 5356 15156
rect 5408 15104 5414 15156
rect 6730 15104 6736 15156
rect 6788 15104 6794 15156
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7834 15144 7840 15156
rect 7524 15116 7840 15144
rect 7524 15104 7530 15116
rect 7834 15104 7840 15116
rect 7892 15144 7898 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7892 15116 7941 15144
rect 7892 15104 7898 15116
rect 7929 15113 7941 15116
rect 7975 15113 7987 15147
rect 7929 15107 7987 15113
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 9180 15116 9229 15144
rect 9180 15104 9186 15116
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 12161 15147 12219 15153
rect 12161 15113 12173 15147
rect 12207 15144 12219 15147
rect 12526 15144 12532 15156
rect 12207 15116 12532 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 14642 15144 14648 15156
rect 14148 15116 14648 15144
rect 14148 15104 14154 15116
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 14752 15116 17540 15144
rect 2682 15036 2688 15088
rect 2740 15076 2746 15088
rect 3136 15079 3194 15085
rect 2740 15048 2912 15076
rect 2740 15036 2746 15048
rect 2884 15017 2912 15048
rect 3136 15045 3148 15079
rect 3182 15076 3194 15079
rect 3418 15076 3424 15088
rect 3182 15048 3424 15076
rect 3182 15045 3194 15048
rect 3136 15039 3194 15045
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 8110 15076 8116 15088
rect 7392 15048 8116 15076
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 4338 14968 4344 15020
rect 4396 14968 4402 15020
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 15008 6239 15011
rect 7190 15008 7196 15020
rect 6227 14980 7196 15008
rect 6227 14977 6239 14980
rect 6181 14971 6239 14977
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 2774 14900 2780 14952
rect 2832 14900 2838 14952
rect 7006 14900 7012 14952
rect 7064 14900 7070 14952
rect 7392 14949 7420 15048
rect 8110 15036 8116 15048
rect 8168 15036 8174 15088
rect 8478 15036 8484 15088
rect 8536 15036 8542 15088
rect 12069 15079 12127 15085
rect 12069 15045 12081 15079
rect 12115 15076 12127 15079
rect 12434 15076 12440 15088
rect 12115 15048 12440 15076
rect 12115 15045 12127 15048
rect 12069 15039 12127 15045
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12621 15079 12679 15085
rect 12621 15045 12633 15079
rect 12667 15076 12679 15079
rect 13924 15076 13952 15104
rect 12667 15048 13952 15076
rect 12667 15045 12679 15048
rect 12621 15039 12679 15045
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7524 14980 7849 15008
rect 7524 14968 7530 14980
rect 7837 14977 7849 14980
rect 7883 15008 7895 15011
rect 8496 15008 8524 15036
rect 12529 15011 12587 15017
rect 7883 14980 8524 15008
rect 9048 14980 10456 15008
rect 7883 14977 7895 14980
rect 7837 14971 7895 14977
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 9048 14949 9076 14980
rect 10428 14952 10456 14980
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 13446 15008 13452 15020
rect 12575 14980 13452 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 8481 14943 8539 14949
rect 8481 14940 8493 14943
rect 7616 14912 8493 14940
rect 7616 14900 7622 14912
rect 8481 14909 8493 14912
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9125 14903 9183 14909
rect 9600 14912 9873 14940
rect 7024 14872 7052 14900
rect 9140 14872 9168 14903
rect 9214 14872 9220 14884
rect 7024 14844 9220 14872
rect 9214 14832 9220 14844
rect 9272 14832 9278 14884
rect 9600 14881 9628 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 10962 14940 10968 14952
rect 10468 14912 10968 14940
rect 10468 14900 10474 14912
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 11256 14912 12817 14940
rect 9585 14875 9643 14881
rect 9585 14841 9597 14875
rect 9631 14841 9643 14875
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 9585 14835 9643 14841
rect 10336 14844 10793 14872
rect 10336 14816 10364 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 11256 14816 11284 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 12434 14832 12440 14884
rect 12492 14832 12498 14884
rect 12820 14872 12848 14903
rect 13170 14900 13176 14952
rect 13228 14900 13234 14952
rect 14752 14940 14780 15116
rect 17512 15085 17540 15116
rect 17586 15104 17592 15156
rect 17644 15104 17650 15156
rect 18969 15147 19027 15153
rect 18969 15113 18981 15147
rect 19015 15144 19027 15147
rect 19058 15144 19064 15156
rect 19015 15116 19064 15144
rect 19015 15113 19027 15116
rect 18969 15107 19027 15113
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 23753 15147 23811 15153
rect 23753 15113 23765 15147
rect 23799 15144 23811 15147
rect 25038 15144 25044 15156
rect 23799 15116 25044 15144
rect 23799 15113 23811 15116
rect 23753 15107 23811 15113
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 25682 15104 25688 15156
rect 25740 15104 25746 15156
rect 29362 15104 29368 15156
rect 29420 15104 29426 15156
rect 30098 15104 30104 15156
rect 30156 15144 30162 15156
rect 32306 15144 32312 15156
rect 30156 15116 32312 15144
rect 30156 15104 30162 15116
rect 32306 15104 32312 15116
rect 32364 15144 32370 15156
rect 36722 15144 36728 15156
rect 32364 15116 36728 15144
rect 32364 15104 32370 15116
rect 36722 15104 36728 15116
rect 36780 15104 36786 15156
rect 37550 15104 37556 15156
rect 37608 15104 37614 15156
rect 42978 15104 42984 15156
rect 43036 15144 43042 15156
rect 43625 15147 43683 15153
rect 43625 15144 43637 15147
rect 43036 15116 43637 15144
rect 43036 15104 43042 15116
rect 43625 15113 43637 15116
rect 43671 15144 43683 15147
rect 44082 15144 44088 15156
rect 43671 15116 44088 15144
rect 43671 15113 43683 15116
rect 43625 15107 43683 15113
rect 44082 15104 44088 15116
rect 44140 15104 44146 15156
rect 49602 15104 49608 15156
rect 49660 15144 49666 15156
rect 49697 15147 49755 15153
rect 49697 15144 49709 15147
rect 49660 15116 49709 15144
rect 49660 15104 49666 15116
rect 49697 15113 49709 15116
rect 49743 15113 49755 15147
rect 49697 15107 49755 15113
rect 50614 15104 50620 15156
rect 50672 15104 50678 15156
rect 50706 15104 50712 15156
rect 50764 15104 50770 15156
rect 52178 15144 52184 15156
rect 51092 15116 52184 15144
rect 17497 15079 17555 15085
rect 17497 15045 17509 15079
rect 17543 15076 17555 15079
rect 17543 15048 18552 15076
rect 17543 15045 17555 15048
rect 17497 15039 17555 15045
rect 18524 15020 18552 15048
rect 23842 15036 23848 15088
rect 23900 15036 23906 15088
rect 24210 15036 24216 15088
rect 24268 15076 24274 15088
rect 24489 15079 24547 15085
rect 24489 15076 24501 15079
rect 24268 15048 24501 15076
rect 24268 15036 24274 15048
rect 24489 15045 24501 15048
rect 24535 15076 24547 15079
rect 25700 15076 25728 15104
rect 24535 15048 25728 15076
rect 24535 15045 24547 15048
rect 24489 15039 24547 15045
rect 30466 15036 30472 15088
rect 30524 15076 30530 15088
rect 31478 15076 31484 15088
rect 30524 15048 31484 15076
rect 30524 15036 30530 15048
rect 31478 15036 31484 15048
rect 31536 15076 31542 15088
rect 35989 15079 36047 15085
rect 31536 15048 31754 15076
rect 31536 15036 31542 15048
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 14884 14980 15148 15008
rect 14884 14968 14890 14980
rect 15120 14949 15148 14980
rect 15194 14968 15200 15020
rect 15252 14968 15258 15020
rect 15286 14968 15292 15020
rect 15344 14968 15350 15020
rect 15387 14980 17816 15008
rect 13280 14912 14780 14940
rect 15105 14943 15163 14949
rect 13280 14872 13308 14912
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15387 14940 15415 14980
rect 17788 14952 17816 14980
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18012 14980 18153 15008
rect 18012 14968 18018 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18414 14968 18420 15020
rect 18472 14968 18478 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 23201 15011 23259 15017
rect 23201 15008 23213 15011
rect 18564 14980 23213 15008
rect 18564 14968 18570 14980
rect 23201 14977 23213 14980
rect 23247 15008 23259 15011
rect 28442 15008 28448 15020
rect 23247 14980 28448 15008
rect 23247 14977 23259 14980
rect 23201 14971 23259 14977
rect 15151 14912 15415 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15746 14900 15752 14952
rect 15804 14900 15810 14952
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 21450 14940 21456 14952
rect 17828 14912 21456 14940
rect 17828 14900 17834 14912
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 23952 14949 23980 14980
rect 28442 14968 28448 14980
rect 28500 14968 28506 15020
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28684 14980 28733 15008
rect 28684 14968 28690 14980
rect 28721 14977 28733 14980
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 30190 14968 30196 15020
rect 30248 14968 30254 15020
rect 23937 14943 23995 14949
rect 23937 14909 23949 14943
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 12820 14844 13308 14872
rect 13740 14844 14780 14872
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 4982 14804 4988 14816
rect 4856 14776 4988 14804
rect 4856 14764 4862 14776
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5534 14764 5540 14816
rect 5592 14764 5598 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 8018 14804 8024 14816
rect 6972 14776 8024 14804
rect 6972 14764 6978 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 9858 14804 9864 14816
rect 8168 14776 9864 14804
rect 8168 14764 8174 14776
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 11238 14764 11244 14816
rect 11296 14764 11302 14816
rect 12452 14804 12480 14832
rect 13740 14804 13768 14844
rect 12452 14776 13768 14804
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 14752 14804 14780 14844
rect 14918 14832 14924 14884
rect 14976 14872 14982 14884
rect 15194 14872 15200 14884
rect 14976 14844 15200 14872
rect 14976 14832 14982 14844
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15654 14832 15660 14884
rect 15712 14832 15718 14884
rect 18046 14872 18052 14884
rect 15764 14844 18052 14872
rect 15764 14804 15792 14844
rect 18046 14832 18052 14844
rect 18104 14872 18110 14884
rect 19242 14872 19248 14884
rect 18104 14844 19248 14872
rect 18104 14832 18110 14844
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 14752 14776 15792 14804
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16393 14807 16451 14813
rect 16393 14804 16405 14807
rect 15896 14776 16405 14804
rect 15896 14764 15902 14776
rect 16393 14773 16405 14776
rect 16439 14773 16451 14807
rect 16393 14767 16451 14773
rect 23382 14764 23388 14816
rect 23440 14764 23446 14816
rect 31478 14764 31484 14816
rect 31536 14764 31542 14816
rect 31726 14804 31754 15048
rect 35989 15045 36001 15079
rect 36035 15076 36047 15079
rect 36538 15076 36544 15088
rect 36035 15048 36544 15076
rect 36035 15045 36047 15048
rect 35989 15039 36047 15045
rect 36538 15036 36544 15048
rect 36596 15076 36602 15088
rect 37568 15076 37596 15104
rect 36596 15048 37596 15076
rect 47848 15079 47906 15085
rect 36596 15036 36602 15048
rect 47848 15045 47860 15079
rect 47894 15076 47906 15079
rect 48682 15076 48688 15088
rect 47894 15048 48688 15076
rect 47894 15045 47906 15048
rect 47848 15039 47906 15045
rect 48682 15036 48688 15048
rect 48740 15036 48746 15088
rect 51092 15076 51120 15116
rect 52178 15104 52184 15116
rect 52236 15104 52242 15156
rect 53653 15147 53711 15153
rect 53653 15113 53665 15147
rect 53699 15144 53711 15147
rect 54110 15144 54116 15156
rect 53699 15116 54116 15144
rect 53699 15113 53711 15116
rect 53653 15107 53711 15113
rect 54110 15104 54116 15116
rect 54168 15104 54174 15156
rect 54481 15147 54539 15153
rect 54481 15113 54493 15147
rect 54527 15144 54539 15147
rect 54846 15144 54852 15156
rect 54527 15116 54852 15144
rect 54527 15113 54539 15116
rect 54481 15107 54539 15113
rect 54846 15104 54852 15116
rect 54904 15104 54910 15156
rect 55030 15104 55036 15156
rect 55088 15144 55094 15156
rect 57790 15144 57796 15156
rect 55088 15116 57796 15144
rect 55088 15104 55094 15116
rect 57790 15104 57796 15116
rect 57848 15104 57854 15156
rect 51046 15048 51120 15076
rect 51844 15079 51902 15085
rect 43070 14968 43076 15020
rect 43128 14968 43134 15020
rect 47581 15011 47639 15017
rect 47581 14977 47593 15011
rect 47627 15008 47639 15011
rect 47670 15008 47676 15020
rect 47627 14980 47676 15008
rect 47627 14977 47639 14980
rect 47581 14971 47639 14977
rect 47670 14968 47676 14980
rect 47728 14968 47734 15020
rect 48406 14968 48412 15020
rect 48464 15008 48470 15020
rect 49326 15008 49332 15020
rect 48464 14980 49332 15008
rect 48464 14968 48470 14980
rect 49326 14968 49332 14980
rect 49384 15008 49390 15020
rect 50249 15011 50307 15017
rect 50249 15008 50261 15011
rect 49384 14980 50261 15008
rect 49384 14968 49390 14980
rect 50249 14977 50261 14980
rect 50295 15008 50307 15011
rect 51046 15008 51074 15048
rect 51844 15045 51856 15079
rect 51890 15076 51902 15079
rect 52454 15076 52460 15088
rect 51890 15048 52460 15076
rect 51890 15045 51902 15048
rect 51844 15039 51902 15045
rect 52454 15036 52460 15048
rect 52512 15036 52518 15088
rect 54202 15036 54208 15088
rect 54260 15036 54266 15088
rect 54941 15079 54999 15085
rect 54941 15045 54953 15079
rect 54987 15076 54999 15079
rect 56226 15076 56232 15088
rect 54987 15048 56232 15076
rect 54987 15045 54999 15048
rect 54941 15039 54999 15045
rect 56226 15036 56232 15048
rect 56284 15036 56290 15088
rect 56588 15079 56646 15085
rect 56588 15045 56600 15079
rect 56634 15076 56646 15079
rect 57330 15076 57336 15088
rect 56634 15048 57336 15076
rect 56634 15045 56646 15048
rect 56588 15039 56646 15045
rect 57330 15036 57336 15048
rect 57388 15036 57394 15088
rect 50295 14980 51074 15008
rect 52089 15011 52147 15017
rect 50295 14977 50307 14980
rect 50249 14971 50307 14977
rect 52089 14977 52101 15011
rect 52135 15008 52147 15011
rect 52362 15008 52368 15020
rect 52135 14980 52368 15008
rect 52135 14977 52147 14980
rect 52089 14971 52147 14977
rect 52362 14968 52368 14980
rect 52420 14968 52426 15020
rect 54021 15011 54079 15017
rect 54021 14977 54033 15011
rect 54067 14977 54079 15011
rect 54021 14971 54079 14977
rect 54113 15011 54171 15017
rect 54113 14977 54125 15011
rect 54159 15008 54171 15011
rect 54220 15008 54248 15036
rect 54849 15011 54907 15017
rect 54849 15008 54861 15011
rect 54159 14980 54861 15008
rect 54159 14977 54171 14980
rect 54113 14971 54171 14977
rect 54849 14977 54861 14980
rect 54895 15008 54907 15011
rect 55122 15008 55128 15020
rect 54895 14980 55128 15008
rect 54895 14977 54907 14980
rect 54849 14971 54907 14977
rect 35618 14940 35624 14952
rect 33244 14912 35624 14940
rect 33134 14872 33140 14884
rect 32784 14844 33140 14872
rect 32784 14816 32812 14844
rect 33134 14832 33140 14844
rect 33192 14832 33198 14884
rect 33244 14816 33272 14912
rect 35618 14900 35624 14912
rect 35676 14900 35682 14952
rect 35986 14900 35992 14952
rect 36044 14940 36050 14952
rect 37277 14943 37335 14949
rect 37277 14940 37289 14943
rect 36044 14912 37289 14940
rect 36044 14900 36050 14912
rect 37277 14909 37289 14912
rect 37323 14909 37335 14943
rect 37277 14903 37335 14909
rect 43346 14900 43352 14952
rect 43404 14940 43410 14952
rect 43717 14943 43775 14949
rect 43717 14940 43729 14943
rect 43404 14912 43729 14940
rect 43404 14900 43410 14912
rect 43717 14909 43729 14912
rect 43763 14909 43775 14943
rect 43717 14903 43775 14909
rect 49053 14943 49111 14949
rect 49053 14909 49065 14943
rect 49099 14909 49111 14943
rect 49053 14903 49111 14909
rect 36265 14875 36323 14881
rect 36265 14872 36277 14875
rect 33612 14844 36277 14872
rect 33612 14816 33640 14844
rect 36265 14841 36277 14844
rect 36311 14841 36323 14875
rect 38102 14872 38108 14884
rect 36265 14835 36323 14841
rect 37752 14844 38108 14872
rect 37752 14816 37780 14844
rect 38102 14832 38108 14844
rect 38160 14832 38166 14884
rect 48961 14875 49019 14881
rect 48961 14841 48973 14875
rect 49007 14872 49019 14875
rect 49068 14872 49096 14903
rect 50062 14900 50068 14952
rect 50120 14900 50126 14952
rect 50157 14943 50215 14949
rect 50157 14909 50169 14943
rect 50203 14940 50215 14943
rect 50890 14940 50896 14952
rect 50203 14912 50896 14940
rect 50203 14909 50215 14912
rect 50157 14903 50215 14909
rect 50890 14900 50896 14912
rect 50948 14900 50954 14952
rect 49007 14844 49096 14872
rect 49007 14841 49019 14844
rect 48961 14835 49019 14841
rect 49602 14832 49608 14884
rect 49660 14872 49666 14884
rect 51074 14872 51080 14884
rect 49660 14844 51080 14872
rect 49660 14832 49666 14844
rect 51074 14832 51080 14844
rect 51132 14832 51138 14884
rect 52086 14832 52092 14884
rect 52144 14872 52150 14884
rect 52362 14872 52368 14884
rect 52144 14844 52368 14872
rect 52144 14832 52150 14844
rect 52362 14832 52368 14844
rect 52420 14832 52426 14884
rect 54036 14872 54064 14971
rect 55122 14968 55128 14980
rect 55180 14968 55186 15020
rect 56134 14968 56140 15020
rect 56192 15008 56198 15020
rect 56321 15011 56379 15017
rect 56321 15008 56333 15011
rect 56192 14980 56333 15008
rect 56192 14968 56198 14980
rect 56321 14977 56333 14980
rect 56367 14977 56379 15011
rect 56321 14971 56379 14977
rect 57606 14968 57612 15020
rect 57664 15008 57670 15020
rect 57885 15011 57943 15017
rect 57885 15008 57897 15011
rect 57664 14980 57897 15008
rect 57664 14968 57670 14980
rect 57885 14977 57897 14980
rect 57931 14977 57943 15011
rect 57885 14971 57943 14977
rect 54202 14900 54208 14952
rect 54260 14900 54266 14952
rect 55030 14900 55036 14952
rect 55088 14900 55094 14952
rect 55306 14900 55312 14952
rect 55364 14900 55370 14952
rect 55953 14875 56011 14881
rect 55953 14872 55965 14875
rect 54036 14844 55965 14872
rect 55953 14841 55965 14844
rect 55999 14872 56011 14875
rect 56042 14872 56048 14884
rect 55999 14844 56048 14872
rect 55999 14841 56011 14844
rect 55953 14835 56011 14841
rect 56042 14832 56048 14844
rect 56100 14832 56106 14884
rect 32401 14807 32459 14813
rect 32401 14804 32413 14807
rect 31726 14776 32413 14804
rect 32401 14773 32413 14776
rect 32447 14804 32459 14807
rect 32766 14804 32772 14816
rect 32447 14776 32772 14804
rect 32447 14773 32459 14776
rect 32401 14767 32459 14773
rect 32766 14764 32772 14776
rect 32824 14764 32830 14816
rect 33045 14807 33103 14813
rect 33045 14773 33057 14807
rect 33091 14804 33103 14807
rect 33226 14804 33232 14816
rect 33091 14776 33232 14804
rect 33091 14773 33103 14776
rect 33045 14767 33103 14773
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 33594 14764 33600 14816
rect 33652 14764 33658 14816
rect 36817 14807 36875 14813
rect 36817 14773 36829 14807
rect 36863 14804 36875 14807
rect 37734 14804 37740 14816
rect 36863 14776 37740 14804
rect 36863 14773 36875 14776
rect 36817 14767 36875 14773
rect 37734 14764 37740 14776
rect 37792 14764 37798 14816
rect 37921 14807 37979 14813
rect 37921 14773 37933 14807
rect 37967 14804 37979 14807
rect 38194 14804 38200 14816
rect 37967 14776 38200 14804
rect 37967 14773 37979 14776
rect 37921 14767 37979 14773
rect 38194 14764 38200 14776
rect 38252 14764 38258 14816
rect 41782 14764 41788 14816
rect 41840 14804 41846 14816
rect 42426 14804 42432 14816
rect 41840 14776 42432 14804
rect 41840 14764 41846 14776
rect 42426 14764 42432 14776
rect 42484 14764 42490 14816
rect 43806 14764 43812 14816
rect 43864 14804 43870 14816
rect 44361 14807 44419 14813
rect 44361 14804 44373 14807
rect 43864 14776 44373 14804
rect 43864 14764 43870 14776
rect 44361 14773 44373 14776
rect 44407 14773 44419 14807
rect 44361 14767 44419 14773
rect 45002 14764 45008 14816
rect 45060 14764 45066 14816
rect 45370 14764 45376 14816
rect 45428 14764 45434 14816
rect 49510 14764 49516 14816
rect 49568 14804 49574 14816
rect 53561 14807 53619 14813
rect 53561 14804 53573 14807
rect 49568 14776 53573 14804
rect 49568 14764 49574 14776
rect 53561 14773 53573 14776
rect 53607 14804 53619 14807
rect 53834 14804 53840 14816
rect 53607 14776 53840 14804
rect 53607 14773 53619 14776
rect 53561 14767 53619 14773
rect 53834 14764 53840 14776
rect 53892 14804 53898 14816
rect 54202 14804 54208 14816
rect 53892 14776 54208 14804
rect 53892 14764 53898 14776
rect 54202 14764 54208 14776
rect 54260 14764 54266 14816
rect 57698 14764 57704 14816
rect 57756 14764 57762 14816
rect 58526 14764 58532 14816
rect 58584 14764 58590 14816
rect 1104 14714 58880 14736
rect 1104 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 22616 14714
rect 22668 14662 22680 14714
rect 22732 14662 22744 14714
rect 22796 14662 22808 14714
rect 22860 14662 22872 14714
rect 22924 14662 37060 14714
rect 37112 14662 37124 14714
rect 37176 14662 37188 14714
rect 37240 14662 37252 14714
rect 37304 14662 37316 14714
rect 37368 14662 51504 14714
rect 51556 14662 51568 14714
rect 51620 14662 51632 14714
rect 51684 14662 51696 14714
rect 51748 14662 51760 14714
rect 51812 14662 58880 14714
rect 1104 14640 58880 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 2832 14572 3801 14600
rect 2832 14560 2838 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 5350 14560 5356 14612
rect 5408 14600 5414 14612
rect 6825 14603 6883 14609
rect 5408 14572 6776 14600
rect 5408 14560 5414 14572
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 4304 14436 4353 14464
rect 4304 14424 4310 14436
rect 4341 14433 4353 14436
rect 4387 14464 4399 14467
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 4387 14436 4813 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 4801 14433 4813 14436
rect 4847 14433 4859 14467
rect 6748 14464 6776 14572
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7558 14600 7564 14612
rect 6871 14572 7564 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8941 14603 8999 14609
rect 8076 14572 8156 14600
rect 8076 14560 8082 14572
rect 8128 14541 8156 14572
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9674 14600 9680 14612
rect 8987 14572 9680 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10502 14560 10508 14612
rect 10560 14560 10566 14612
rect 12434 14560 12440 14612
rect 12492 14560 12498 14612
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 13170 14600 13176 14612
rect 12943 14572 13176 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 15286 14600 15292 14612
rect 14139 14572 15292 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 23198 14560 23204 14612
rect 23256 14560 23262 14612
rect 23382 14560 23388 14612
rect 23440 14560 23446 14612
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 24210 14600 24216 14612
rect 23624 14572 24216 14600
rect 23624 14560 23630 14572
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 29730 14600 29736 14612
rect 26108 14572 29736 14600
rect 26108 14560 26114 14572
rect 29730 14560 29736 14572
rect 29788 14560 29794 14612
rect 30098 14560 30104 14612
rect 30156 14560 30162 14612
rect 35253 14603 35311 14609
rect 35253 14569 35265 14603
rect 35299 14600 35311 14603
rect 35526 14600 35532 14612
rect 35299 14572 35532 14600
rect 35299 14569 35311 14572
rect 35253 14563 35311 14569
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 37734 14600 37740 14612
rect 37200 14572 37740 14600
rect 8113 14535 8171 14541
rect 8113 14501 8125 14535
rect 8159 14532 8171 14535
rect 8754 14532 8760 14544
rect 8159 14504 8760 14532
rect 8159 14501 8171 14504
rect 8113 14495 8171 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 9214 14492 9220 14544
rect 9272 14492 9278 14544
rect 7190 14464 7196 14476
rect 6748 14436 7196 14464
rect 4801 14427 4859 14433
rect 7190 14424 7196 14436
rect 7248 14464 7254 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7248 14436 7573 14464
rect 7248 14424 7254 14436
rect 7561 14433 7573 14436
rect 7607 14464 7619 14467
rect 8018 14464 8024 14476
rect 7607 14436 8024 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9122 14464 9128 14476
rect 8619 14436 9128 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4982 14396 4988 14408
rect 4203 14368 4988 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5994 14396 6000 14408
rect 5491 14368 6000 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 7742 14405 7748 14408
rect 7720 14399 7748 14405
rect 7720 14365 7732 14399
rect 7720 14359 7748 14365
rect 7742 14356 7748 14359
rect 7800 14356 7806 14408
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 8846 14396 8852 14408
rect 8803 14368 8852 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 4430 14328 4436 14340
rect 4295 14300 4436 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 4430 14288 4436 14300
rect 4488 14288 4494 14340
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 5690 14331 5748 14337
rect 5690 14328 5702 14331
rect 5592 14300 5702 14328
rect 5592 14288 5598 14300
rect 5690 14297 5702 14300
rect 5736 14297 5748 14331
rect 9232 14328 9260 14492
rect 10520 14464 10548 14560
rect 12452 14532 12480 14560
rect 12452 14504 13584 14532
rect 10244 14436 10548 14464
rect 10065 14399 10123 14405
rect 10065 14365 10077 14399
rect 10111 14396 10123 14399
rect 10244 14396 10272 14436
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 11054 14464 11060 14476
rect 10652 14436 11060 14464
rect 10652 14424 10658 14436
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 13556 14473 13584 14504
rect 15194 14492 15200 14544
rect 15252 14492 15258 14544
rect 17957 14535 18015 14541
rect 17957 14501 17969 14535
rect 18003 14532 18015 14535
rect 18690 14532 18696 14544
rect 18003 14504 18696 14532
rect 18003 14501 18015 14504
rect 17957 14495 18015 14501
rect 18690 14492 18696 14504
rect 18748 14532 18754 14544
rect 22922 14532 22928 14544
rect 18748 14504 22928 14532
rect 18748 14492 18754 14504
rect 22922 14492 22928 14504
rect 22980 14492 22986 14544
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14433 13599 14467
rect 13814 14464 13820 14476
rect 13541 14427 13599 14433
rect 13740 14436 13820 14464
rect 10111 14368 10272 14396
rect 10111 14365 10123 14368
rect 10065 14359 10123 14365
rect 10318 14356 10324 14408
rect 10376 14396 10382 14408
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 10376 14368 11529 14396
rect 10376 14356 10382 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 13740 14396 13768 14436
rect 13814 14424 13820 14436
rect 13872 14464 13878 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 13872 14436 15025 14464
rect 13872 14424 13878 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15212 14464 15240 14492
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15212 14436 15301 14464
rect 15013 14427 15071 14433
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16114 14464 16120 14476
rect 15795 14436 16120 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 16114 14424 16120 14436
rect 16172 14464 16178 14476
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16172 14436 16405 14464
rect 16172 14424 16178 14436
rect 16393 14433 16405 14436
rect 16439 14433 16451 14467
rect 16393 14427 16451 14433
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19852 14436 20085 14464
rect 19852 14424 19858 14436
rect 20073 14433 20085 14436
rect 20119 14464 20131 14467
rect 23400 14464 23428 14560
rect 26068 14532 26096 14560
rect 29549 14535 29607 14541
rect 29549 14532 29561 14535
rect 23860 14504 26096 14532
rect 29380 14504 29561 14532
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 20119 14436 23143 14464
rect 23400 14436 23765 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 13495 14368 13768 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 13906 14356 13912 14408
rect 13964 14356 13970 14408
rect 14734 14356 14740 14408
rect 14792 14356 14798 14408
rect 14826 14356 14832 14408
rect 14884 14405 14890 14408
rect 14884 14399 14933 14405
rect 14884 14365 14887 14399
rect 14921 14365 14933 14399
rect 14884 14359 14933 14365
rect 14884 14356 14890 14359
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15896 14368 15945 14396
rect 15896 14356 15902 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 16942 14356 16948 14408
rect 17000 14356 17006 14408
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 19760 14368 20269 14396
rect 19760 14356 19766 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 21450 14356 21456 14408
rect 21508 14356 21514 14408
rect 23115 14396 23143 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23860 14396 23888 14504
rect 24946 14424 24952 14476
rect 25004 14424 25010 14476
rect 29380 14473 29408 14504
rect 29549 14501 29561 14504
rect 29595 14501 29607 14535
rect 29549 14495 29607 14501
rect 30116 14473 30144 14560
rect 32953 14535 33011 14541
rect 32953 14501 32965 14535
rect 32999 14532 33011 14535
rect 32999 14504 34376 14532
rect 32999 14501 33011 14504
rect 32953 14495 33011 14501
rect 26145 14467 26203 14473
rect 26145 14433 26157 14467
rect 26191 14433 26203 14467
rect 26145 14427 26203 14433
rect 29365 14467 29423 14473
rect 29365 14433 29377 14467
rect 29411 14433 29423 14467
rect 29365 14427 29423 14433
rect 30101 14467 30159 14473
rect 30101 14433 30113 14467
rect 30147 14433 30159 14467
rect 31941 14467 31999 14473
rect 31941 14464 31953 14467
rect 30101 14427 30159 14433
rect 30208 14436 31953 14464
rect 23115 14368 23888 14396
rect 25958 14356 25964 14408
rect 26016 14356 26022 14408
rect 10781 14331 10839 14337
rect 10781 14328 10793 14331
rect 9232 14300 10793 14328
rect 5690 14291 5748 14297
rect 10781 14297 10793 14300
rect 10827 14297 10839 14331
rect 10781 14291 10839 14297
rect 11784 14331 11842 14337
rect 11784 14297 11796 14331
rect 11830 14328 11842 14331
rect 12434 14328 12440 14340
rect 11830 14300 12440 14328
rect 11830 14297 11842 14300
rect 11784 14291 11842 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13924 14328 13952 14356
rect 13403 14300 13952 14328
rect 19061 14331 19119 14337
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 19061 14297 19073 14331
rect 19107 14328 19119 14331
rect 19334 14328 19340 14340
rect 19107 14300 19340 14328
rect 19107 14297 19119 14300
rect 19061 14291 19119 14297
rect 19334 14288 19340 14300
rect 19392 14328 19398 14340
rect 21468 14328 21496 14356
rect 25409 14331 25467 14337
rect 25409 14328 25421 14331
rect 19392 14300 20116 14328
rect 21468 14300 25421 14328
rect 19392 14288 19398 14300
rect 20088 14272 20116 14300
rect 25409 14297 25421 14300
rect 25455 14328 25467 14331
rect 26160 14328 26188 14427
rect 26418 14356 26424 14408
rect 26476 14396 26482 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26476 14368 26985 14396
rect 26476 14356 26482 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 29730 14356 29736 14408
rect 29788 14396 29794 14408
rect 30208 14396 30236 14436
rect 31941 14433 31953 14436
rect 31987 14433 31999 14467
rect 31941 14427 31999 14433
rect 32309 14467 32367 14473
rect 32309 14433 32321 14467
rect 32355 14433 32367 14467
rect 32309 14427 32367 14433
rect 29788 14368 30236 14396
rect 29788 14356 29794 14368
rect 30282 14356 30288 14408
rect 30340 14396 30346 14408
rect 30926 14396 30932 14408
rect 30340 14368 30932 14396
rect 30340 14356 30346 14368
rect 30926 14356 30932 14368
rect 30984 14356 30990 14408
rect 31202 14356 31208 14408
rect 31260 14356 31266 14408
rect 25455 14300 26188 14328
rect 29917 14331 29975 14337
rect 25455 14297 25467 14300
rect 25409 14291 25467 14297
rect 29917 14297 29929 14331
rect 29963 14328 29975 14331
rect 31018 14328 31024 14340
rect 29963 14300 31024 14328
rect 29963 14297 29975 14300
rect 29917 14291 29975 14297
rect 31018 14288 31024 14300
rect 31076 14328 31082 14340
rect 31389 14331 31447 14337
rect 31389 14328 31401 14331
rect 31076 14300 31401 14328
rect 31076 14288 31082 14300
rect 31389 14297 31401 14300
rect 31435 14297 31447 14331
rect 32324 14328 32352 14427
rect 32398 14424 32404 14476
rect 32456 14464 32462 14476
rect 34348 14473 34376 14504
rect 33045 14467 33103 14473
rect 33045 14464 33057 14467
rect 32456 14436 33057 14464
rect 32456 14424 32462 14436
rect 33045 14433 33057 14436
rect 33091 14433 33103 14467
rect 33045 14427 33103 14433
rect 34333 14467 34391 14473
rect 34333 14433 34345 14467
rect 34379 14433 34391 14467
rect 35544 14464 35572 14560
rect 37200 14532 37228 14572
rect 37734 14560 37740 14572
rect 37792 14560 37798 14612
rect 38749 14603 38807 14609
rect 38749 14569 38761 14603
rect 38795 14600 38807 14603
rect 39022 14600 39028 14612
rect 38795 14572 39028 14600
rect 38795 14569 38807 14572
rect 38749 14563 38807 14569
rect 39022 14560 39028 14572
rect 39080 14560 39086 14612
rect 39117 14603 39175 14609
rect 39117 14569 39129 14603
rect 39163 14600 39175 14603
rect 39390 14600 39396 14612
rect 39163 14572 39396 14600
rect 39163 14569 39175 14572
rect 39117 14563 39175 14569
rect 39390 14560 39396 14572
rect 39448 14600 39454 14612
rect 44729 14603 44787 14609
rect 44729 14600 44741 14603
rect 39448 14572 44741 14600
rect 39448 14560 39454 14572
rect 44729 14569 44741 14572
rect 44775 14569 44787 14603
rect 44729 14563 44787 14569
rect 50157 14603 50215 14609
rect 50157 14569 50169 14603
rect 50203 14600 50215 14603
rect 51258 14600 51264 14612
rect 50203 14572 51264 14600
rect 50203 14569 50215 14572
rect 50157 14563 50215 14569
rect 37108 14504 37228 14532
rect 37645 14535 37703 14541
rect 37108 14473 37136 14504
rect 37645 14501 37657 14535
rect 37691 14532 37703 14535
rect 37691 14504 38332 14532
rect 37691 14501 37703 14504
rect 37645 14495 37703 14501
rect 38304 14473 38332 14504
rect 40034 14492 40040 14544
rect 40092 14492 40098 14544
rect 41877 14535 41935 14541
rect 41877 14501 41889 14535
rect 41923 14501 41935 14535
rect 41877 14495 41935 14501
rect 35897 14467 35955 14473
rect 35897 14464 35909 14467
rect 35544 14436 35909 14464
rect 34333 14427 34391 14433
rect 35897 14433 35909 14436
rect 35943 14433 35955 14467
rect 37093 14467 37151 14473
rect 35897 14427 35955 14433
rect 36648 14436 37044 14464
rect 32585 14399 32643 14405
rect 32585 14365 32597 14399
rect 32631 14396 32643 14399
rect 32674 14396 32680 14408
rect 32631 14368 32680 14396
rect 32631 14365 32643 14368
rect 32585 14359 32643 14365
rect 32674 14356 32680 14368
rect 32732 14356 32738 14408
rect 35805 14399 35863 14405
rect 35805 14365 35817 14399
rect 35851 14396 35863 14399
rect 36648 14396 36676 14436
rect 35851 14368 36676 14396
rect 35851 14365 35863 14368
rect 35805 14359 35863 14365
rect 36722 14356 36728 14408
rect 36780 14356 36786 14408
rect 37016 14396 37044 14436
rect 37093 14433 37105 14467
rect 37139 14433 37151 14467
rect 37093 14427 37151 14433
rect 38289 14467 38347 14473
rect 38289 14433 38301 14467
rect 38335 14433 38347 14467
rect 38289 14427 38347 14433
rect 38746 14424 38752 14476
rect 38804 14464 38810 14476
rect 39114 14464 39120 14476
rect 38804 14436 39120 14464
rect 38804 14424 38810 14436
rect 39114 14424 39120 14436
rect 39172 14424 39178 14476
rect 41785 14467 41843 14473
rect 41785 14433 41797 14467
rect 41831 14464 41843 14467
rect 41892 14464 41920 14495
rect 41831 14436 41920 14464
rect 41831 14433 41843 14436
rect 41785 14427 41843 14433
rect 42426 14424 42432 14476
rect 42484 14424 42490 14476
rect 42702 14424 42708 14476
rect 42760 14464 42766 14476
rect 43257 14467 43315 14473
rect 43257 14464 43269 14467
rect 42760 14436 43269 14464
rect 42760 14424 42766 14436
rect 43257 14433 43269 14436
rect 43303 14433 43315 14467
rect 43898 14464 43904 14476
rect 43257 14427 43315 14433
rect 43456 14436 43904 14464
rect 37274 14396 37280 14408
rect 37016 14368 37280 14396
rect 37274 14356 37280 14368
rect 37332 14396 37338 14408
rect 37458 14396 37464 14408
rect 37332 14368 37464 14396
rect 37332 14356 37338 14368
rect 37458 14356 37464 14368
rect 37516 14396 37522 14408
rect 38470 14396 38476 14408
rect 37516 14368 38476 14396
rect 37516 14356 37522 14368
rect 38470 14356 38476 14368
rect 38528 14356 38534 14408
rect 40218 14356 40224 14408
rect 40276 14356 40282 14408
rect 42245 14399 42303 14405
rect 42245 14365 42257 14399
rect 42291 14396 42303 14399
rect 43456 14396 43484 14436
rect 43898 14424 43904 14436
rect 43956 14464 43962 14476
rect 44177 14467 44235 14473
rect 44177 14464 44189 14467
rect 43956 14436 44189 14464
rect 43956 14424 43962 14436
rect 44177 14433 44189 14436
rect 44223 14433 44235 14467
rect 44744 14464 44772 14563
rect 51258 14560 51264 14572
rect 51316 14560 51322 14612
rect 54481 14603 54539 14609
rect 51368 14572 54064 14600
rect 51368 14541 51396 14572
rect 51353 14535 51411 14541
rect 45112 14504 47440 14532
rect 45112 14473 45140 14504
rect 45097 14467 45155 14473
rect 45097 14464 45109 14467
rect 44744 14436 45109 14464
rect 44177 14427 44235 14433
rect 45097 14433 45109 14436
rect 45143 14433 45155 14467
rect 45097 14427 45155 14433
rect 45278 14424 45284 14476
rect 45336 14424 45342 14476
rect 47412 14464 47440 14504
rect 51353 14501 51365 14535
rect 51399 14501 51411 14535
rect 54036 14532 54064 14572
rect 54481 14569 54493 14603
rect 54527 14600 54539 14603
rect 55306 14600 55312 14612
rect 54527 14572 55312 14600
rect 54527 14569 54539 14572
rect 54481 14563 54539 14569
rect 55306 14560 55312 14572
rect 55364 14560 55370 14612
rect 55600 14572 56456 14600
rect 54938 14532 54944 14544
rect 54036 14504 54944 14532
rect 51353 14495 51411 14501
rect 47412 14436 47532 14464
rect 42291 14368 43484 14396
rect 42291 14365 42303 14368
rect 42245 14359 42303 14365
rect 43530 14356 43536 14408
rect 43588 14356 43594 14408
rect 47397 14399 47455 14405
rect 47397 14396 47409 14399
rect 47320 14368 47409 14396
rect 33226 14328 33232 14340
rect 32324 14300 33232 14328
rect 31389 14291 31447 14297
rect 33226 14288 33232 14300
rect 33284 14288 33290 14340
rect 35713 14331 35771 14337
rect 35713 14297 35725 14331
rect 35759 14328 35771 14331
rect 36630 14328 36636 14340
rect 35759 14300 36636 14328
rect 35759 14297 35771 14300
rect 35713 14291 35771 14297
rect 36630 14288 36636 14300
rect 36688 14288 36694 14340
rect 37642 14288 37648 14340
rect 37700 14328 37706 14340
rect 40770 14328 40776 14340
rect 37700 14300 40776 14328
rect 37700 14288 37706 14300
rect 40770 14288 40776 14300
rect 40828 14288 40834 14340
rect 42337 14331 42395 14337
rect 42337 14297 42349 14331
rect 42383 14328 42395 14331
rect 42794 14328 42800 14340
rect 42383 14300 42800 14328
rect 42383 14297 42395 14300
rect 42337 14291 42395 14297
rect 42794 14288 42800 14300
rect 42852 14328 42858 14340
rect 43165 14331 43223 14337
rect 42852 14300 43116 14328
rect 42852 14288 42858 14300
rect 6914 14220 6920 14272
rect 6972 14220 6978 14272
rect 10410 14220 10416 14272
rect 10468 14220 10474 14272
rect 10870 14220 10876 14272
rect 10928 14220 10934 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 12526 14260 12532 14272
rect 11020 14232 12532 14260
rect 11020 14220 11026 14232
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 12986 14220 12992 14272
rect 13044 14220 13050 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14826 14260 14832 14272
rect 13504 14232 14832 14260
rect 13504 14220 13510 14232
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 20070 14220 20076 14272
rect 20128 14220 20134 14272
rect 20162 14220 20168 14272
rect 20220 14220 20226 14272
rect 20625 14263 20683 14269
rect 20625 14229 20637 14263
rect 20671 14260 20683 14263
rect 21174 14260 21180 14272
rect 20671 14232 21180 14260
rect 20671 14229 20683 14232
rect 20625 14223 20683 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21358 14220 21364 14272
rect 21416 14220 21422 14272
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 23658 14260 23664 14272
rect 22980 14232 23664 14260
rect 22980 14220 22986 14232
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25590 14220 25596 14272
rect 25648 14220 25654 14272
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 26053 14263 26111 14269
rect 26053 14260 26065 14263
rect 25740 14232 26065 14260
rect 25740 14220 25746 14232
rect 26053 14229 26065 14232
rect 26099 14229 26111 14263
rect 26053 14223 26111 14229
rect 26142 14220 26148 14272
rect 26200 14260 26206 14272
rect 26421 14263 26479 14269
rect 26421 14260 26433 14263
rect 26200 14232 26433 14260
rect 26200 14220 26206 14232
rect 26421 14229 26433 14232
rect 26467 14229 26479 14263
rect 26421 14223 26479 14229
rect 28718 14220 28724 14272
rect 28776 14220 28782 14272
rect 30009 14263 30067 14269
rect 30009 14229 30021 14263
rect 30055 14260 30067 14263
rect 30282 14260 30288 14272
rect 30055 14232 30288 14260
rect 30055 14229 30067 14232
rect 30009 14223 30067 14229
rect 30282 14220 30288 14232
rect 30340 14220 30346 14272
rect 30650 14220 30656 14272
rect 30708 14220 30714 14272
rect 32490 14220 32496 14272
rect 32548 14220 32554 14272
rect 33502 14220 33508 14272
rect 33560 14260 33566 14272
rect 33689 14263 33747 14269
rect 33689 14260 33701 14263
rect 33560 14232 33701 14260
rect 33560 14220 33566 14232
rect 33689 14229 33701 14232
rect 33735 14229 33747 14263
rect 33689 14223 33747 14229
rect 33778 14220 33784 14272
rect 33836 14220 33842 14272
rect 35342 14220 35348 14272
rect 35400 14220 35406 14272
rect 35894 14220 35900 14272
rect 35952 14260 35958 14272
rect 36173 14263 36231 14269
rect 36173 14260 36185 14263
rect 35952 14232 36185 14260
rect 35952 14220 35958 14232
rect 36173 14229 36185 14232
rect 36219 14229 36231 14263
rect 36173 14223 36231 14229
rect 37185 14263 37243 14269
rect 37185 14229 37197 14263
rect 37231 14260 37243 14263
rect 37366 14260 37372 14272
rect 37231 14232 37372 14260
rect 37231 14229 37243 14232
rect 37185 14223 37243 14229
rect 37366 14220 37372 14232
rect 37424 14220 37430 14272
rect 37737 14263 37795 14269
rect 37737 14229 37749 14263
rect 37783 14260 37795 14263
rect 37918 14260 37924 14272
rect 37783 14232 37924 14260
rect 37783 14229 37795 14232
rect 37737 14223 37795 14229
rect 37918 14220 37924 14232
rect 37976 14220 37982 14272
rect 38286 14220 38292 14272
rect 38344 14260 38350 14272
rect 38654 14260 38660 14272
rect 38344 14232 38660 14260
rect 38344 14220 38350 14232
rect 38654 14220 38660 14232
rect 38712 14220 38718 14272
rect 40862 14220 40868 14272
rect 40920 14220 40926 14272
rect 41138 14220 41144 14272
rect 41196 14220 41202 14272
rect 42705 14263 42763 14269
rect 42705 14229 42717 14263
rect 42751 14260 42763 14263
rect 42886 14260 42892 14272
rect 42751 14232 42892 14260
rect 42751 14229 42763 14232
rect 42705 14223 42763 14229
rect 42886 14220 42892 14232
rect 42944 14220 42950 14272
rect 43088 14269 43116 14300
rect 43165 14297 43177 14331
rect 43211 14328 43223 14331
rect 43806 14328 43812 14340
rect 43211 14300 43812 14328
rect 43211 14297 43223 14300
rect 43165 14291 43223 14297
rect 43806 14288 43812 14300
rect 43864 14288 43870 14340
rect 47320 14272 47348 14368
rect 47397 14365 47409 14368
rect 47443 14365 47455 14399
rect 47504 14396 47532 14436
rect 49326 14424 49332 14476
rect 49384 14424 49390 14476
rect 49510 14424 49516 14476
rect 49568 14424 49574 14476
rect 49694 14464 49700 14476
rect 49620 14436 49700 14464
rect 49237 14399 49295 14405
rect 47504 14368 49188 14396
rect 47397 14359 47455 14365
rect 47664 14331 47722 14337
rect 47664 14297 47676 14331
rect 47710 14328 47722 14331
rect 48314 14328 48320 14340
rect 47710 14300 48320 14328
rect 47710 14297 47722 14300
rect 47664 14291 47722 14297
rect 48314 14288 48320 14300
rect 48372 14288 48378 14340
rect 49160 14328 49188 14368
rect 49237 14365 49249 14399
rect 49283 14396 49295 14399
rect 49620 14396 49648 14436
rect 49694 14424 49700 14436
rect 49752 14464 49758 14476
rect 50939 14467 50997 14473
rect 50939 14464 50951 14467
rect 49752 14436 50951 14464
rect 49752 14424 49758 14436
rect 50939 14433 50951 14436
rect 50985 14433 50997 14467
rect 50939 14427 50997 14433
rect 51074 14424 51080 14476
rect 51132 14424 51138 14476
rect 51258 14424 51264 14476
rect 51316 14464 51322 14476
rect 51368 14464 51396 14495
rect 54938 14492 54944 14504
rect 54996 14532 55002 14544
rect 55600 14532 55628 14572
rect 54996 14504 55628 14532
rect 54996 14492 55002 14504
rect 51316 14436 51396 14464
rect 51813 14467 51871 14473
rect 51316 14424 51322 14436
rect 51813 14433 51825 14467
rect 51859 14464 51871 14467
rect 52362 14464 52368 14476
rect 51859 14436 52368 14464
rect 51859 14433 51871 14436
rect 51813 14427 51871 14433
rect 52362 14424 52368 14436
rect 52420 14424 52426 14476
rect 55582 14424 55588 14476
rect 55640 14464 55646 14476
rect 55953 14467 56011 14473
rect 55953 14464 55965 14467
rect 55640 14436 55965 14464
rect 55640 14424 55646 14436
rect 55953 14433 55965 14436
rect 55999 14433 56011 14467
rect 55953 14427 56011 14433
rect 56042 14424 56048 14476
rect 56100 14473 56106 14476
rect 56100 14467 56149 14473
rect 56100 14433 56103 14467
rect 56137 14433 56149 14467
rect 56100 14427 56149 14433
rect 56100 14424 56106 14427
rect 56226 14424 56232 14476
rect 56284 14424 56290 14476
rect 56428 14464 56456 14572
rect 56502 14560 56508 14612
rect 56560 14600 56566 14612
rect 56560 14572 57744 14600
rect 56560 14560 56566 14572
rect 56505 14467 56563 14473
rect 56505 14464 56517 14467
rect 56428 14436 56517 14464
rect 56505 14433 56517 14436
rect 56551 14433 56563 14467
rect 56505 14427 56563 14433
rect 56778 14424 56784 14476
rect 56836 14464 56842 14476
rect 57716 14473 57744 14572
rect 57149 14467 57207 14473
rect 57149 14464 57161 14467
rect 56836 14436 57161 14464
rect 56836 14424 56842 14436
rect 57149 14433 57161 14436
rect 57195 14433 57207 14467
rect 57149 14427 57207 14433
rect 57701 14467 57759 14473
rect 57701 14433 57713 14467
rect 57747 14433 57759 14467
rect 57701 14427 57759 14433
rect 49878 14396 49884 14408
rect 49283 14368 49648 14396
rect 49804 14368 49884 14396
rect 49283 14365 49295 14368
rect 49237 14359 49295 14365
rect 49804 14328 49832 14368
rect 49878 14356 49884 14368
rect 49936 14356 49942 14408
rect 50798 14356 50804 14408
rect 50856 14356 50862 14408
rect 51994 14356 52000 14408
rect 52052 14356 52058 14408
rect 53374 14405 53380 14408
rect 53101 14399 53159 14405
rect 53101 14396 53113 14399
rect 53024 14368 53113 14396
rect 49160 14300 49832 14328
rect 53024 14272 53052 14368
rect 53101 14365 53113 14368
rect 53147 14365 53159 14399
rect 53368 14396 53380 14405
rect 53335 14368 53380 14396
rect 53101 14359 53159 14365
rect 53368 14359 53380 14368
rect 53374 14356 53380 14359
rect 53432 14356 53438 14408
rect 56962 14356 56968 14408
rect 57020 14356 57026 14408
rect 57164 14396 57192 14427
rect 57790 14424 57796 14476
rect 57848 14464 57854 14476
rect 58253 14467 58311 14473
rect 58253 14464 58265 14467
rect 57848 14436 58265 14464
rect 57848 14424 57854 14436
rect 58253 14433 58265 14436
rect 58299 14433 58311 14467
rect 58253 14427 58311 14433
rect 57882 14396 57888 14408
rect 57164 14368 57888 14396
rect 57882 14356 57888 14368
rect 57940 14356 57946 14408
rect 57609 14331 57667 14337
rect 57609 14328 57621 14331
rect 56980 14300 57621 14328
rect 43073 14263 43131 14269
rect 43073 14229 43085 14263
rect 43119 14260 43131 14263
rect 43438 14260 43444 14272
rect 43119 14232 43444 14260
rect 43119 14229 43131 14232
rect 43073 14223 43131 14229
rect 43438 14220 43444 14232
rect 43496 14220 43502 14272
rect 45373 14263 45431 14269
rect 45373 14229 45385 14263
rect 45419 14260 45431 14263
rect 45462 14260 45468 14272
rect 45419 14232 45468 14260
rect 45419 14229 45431 14232
rect 45373 14223 45431 14229
rect 45462 14220 45468 14232
rect 45520 14220 45526 14272
rect 45738 14220 45744 14272
rect 45796 14220 45802 14272
rect 47302 14220 47308 14272
rect 47360 14220 47366 14272
rect 48774 14220 48780 14272
rect 48832 14220 48838 14272
rect 48866 14220 48872 14272
rect 48924 14220 48930 14272
rect 49970 14220 49976 14272
rect 50028 14260 50034 14272
rect 53006 14260 53012 14272
rect 50028 14232 53012 14260
rect 50028 14220 50034 14232
rect 53006 14220 53012 14232
rect 53064 14220 53070 14272
rect 54849 14263 54907 14269
rect 54849 14229 54861 14263
rect 54895 14260 54907 14263
rect 55030 14260 55036 14272
rect 54895 14232 55036 14260
rect 54895 14229 54907 14232
rect 54849 14223 54907 14229
rect 55030 14220 55036 14232
rect 55088 14220 55094 14272
rect 55309 14263 55367 14269
rect 55309 14229 55321 14263
rect 55355 14260 55367 14263
rect 56980 14260 57008 14300
rect 57609 14297 57621 14300
rect 57655 14297 57667 14331
rect 57609 14291 57667 14297
rect 55355 14232 57008 14260
rect 55355 14229 55367 14232
rect 55309 14223 55367 14229
rect 57238 14220 57244 14272
rect 57296 14220 57302 14272
rect 1104 14170 59040 14192
rect 1104 14118 15394 14170
rect 15446 14118 15458 14170
rect 15510 14118 15522 14170
rect 15574 14118 15586 14170
rect 15638 14118 15650 14170
rect 15702 14118 29838 14170
rect 29890 14118 29902 14170
rect 29954 14118 29966 14170
rect 30018 14118 30030 14170
rect 30082 14118 30094 14170
rect 30146 14118 44282 14170
rect 44334 14118 44346 14170
rect 44398 14118 44410 14170
rect 44462 14118 44474 14170
rect 44526 14118 44538 14170
rect 44590 14118 58726 14170
rect 58778 14118 58790 14170
rect 58842 14118 58854 14170
rect 58906 14118 58918 14170
rect 58970 14118 58982 14170
rect 59034 14118 59040 14170
rect 1104 14096 59040 14118
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7285 14059 7343 14065
rect 7285 14056 7297 14059
rect 6972 14028 7297 14056
rect 6972 14016 6978 14028
rect 7285 14025 7297 14028
rect 7331 14025 7343 14059
rect 7285 14019 7343 14025
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8662 14056 8668 14068
rect 8067 14028 8668 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 7156 13960 7389 13988
rect 7156 13948 7162 13960
rect 7377 13957 7389 13960
rect 7423 13957 7435 13991
rect 7377 13951 7435 13957
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7282 13852 7288 13864
rect 7156 13824 7288 13852
rect 7156 13812 7162 13824
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7834 13852 7840 13864
rect 7607 13824 7840 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 8036 13852 8064 14019
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 12894 14016 12900 14068
rect 12952 14016 12958 14068
rect 14826 14056 14832 14068
rect 13372 14028 14832 14056
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 8297 13991 8355 13997
rect 8297 13988 8309 13991
rect 8168 13960 8309 13988
rect 8168 13948 8174 13960
rect 8297 13957 8309 13960
rect 8343 13988 8355 13991
rect 9490 13988 9496 14000
rect 8343 13960 9496 13988
rect 8343 13957 8355 13960
rect 8297 13951 8355 13957
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 9616 13991 9674 13997
rect 9616 13957 9628 13991
rect 9662 13988 9674 13991
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 9662 13960 10057 13988
rect 9662 13957 9674 13960
rect 9616 13951 9674 13957
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10045 13951 10103 13957
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 11333 13991 11391 13997
rect 11333 13988 11345 13991
rect 11112 13960 11345 13988
rect 11112 13948 11118 13960
rect 11333 13957 11345 13960
rect 11379 13988 11391 13991
rect 11784 13991 11842 13997
rect 11379 13960 11652 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 10336 13892 11529 13920
rect 10336 13864 10364 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11624 13920 11652 13960
rect 11784 13957 11796 13991
rect 11830 13988 11842 13991
rect 11974 13988 11980 14000
rect 11830 13960 11980 13988
rect 11830 13957 11842 13960
rect 11784 13951 11842 13957
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 12342 13920 12348 13932
rect 11624 13892 12348 13920
rect 11517 13883 11575 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 13372 13864 13400 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 14921 14059 14979 14065
rect 14921 14025 14933 14059
rect 14967 14056 14979 14059
rect 15746 14056 15752 14068
rect 14967 14028 15752 14056
rect 14967 14025 14979 14028
rect 14921 14019 14979 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 16485 14059 16543 14065
rect 16485 14025 16497 14059
rect 16531 14056 16543 14059
rect 16942 14056 16948 14068
rect 16531 14028 16948 14056
rect 16531 14025 16543 14028
rect 16485 14019 16543 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 13630 13948 13636 14000
rect 13688 13988 13694 14000
rect 13688 13960 15148 13988
rect 13688 13948 13694 13960
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13648 13920 13676 13948
rect 15120 13932 15148 13960
rect 13814 13929 13820 13932
rect 13587 13892 13676 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13808 13883 13820 13929
rect 13814 13880 13820 13883
rect 13872 13880 13878 13932
rect 15102 13880 15108 13932
rect 15160 13880 15166 13932
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15361 13923 15419 13929
rect 15361 13920 15373 13923
rect 15252 13892 15373 13920
rect 15252 13880 15258 13892
rect 15361 13889 15373 13892
rect 15407 13889 15419 13923
rect 15361 13883 15419 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13920 18015 13923
rect 18064 13920 18092 14019
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18417 14059 18475 14065
rect 18417 14025 18429 14059
rect 18463 14056 18475 14059
rect 19334 14056 19340 14068
rect 18463 14028 19340 14056
rect 18463 14025 18475 14028
rect 18417 14019 18475 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 20806 14016 20812 14068
rect 20864 14016 20870 14068
rect 23109 14059 23167 14065
rect 23109 14025 23121 14059
rect 23155 14025 23167 14059
rect 23109 14019 23167 14025
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 23523 14028 24593 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 24581 14025 24593 14028
rect 24627 14056 24639 14059
rect 25406 14056 25412 14068
rect 24627 14028 25412 14056
rect 24627 14025 24639 14028
rect 24581 14019 24639 14025
rect 18340 13988 18368 14016
rect 18509 13991 18567 13997
rect 18509 13988 18521 13991
rect 18340 13960 18521 13988
rect 18509 13957 18521 13960
rect 18555 13988 18567 13991
rect 18782 13988 18788 14000
rect 18555 13960 18788 13988
rect 18555 13957 18567 13960
rect 18509 13951 18567 13957
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 18003 13892 18092 13920
rect 19429 13923 19487 13929
rect 18003 13889 18015 13892
rect 17957 13883 18015 13889
rect 19429 13889 19441 13923
rect 19475 13920 19487 13923
rect 19518 13920 19524 13932
rect 19475 13892 19524 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19702 13929 19708 13932
rect 19696 13883 19708 13929
rect 19702 13880 19708 13883
rect 19760 13880 19766 13932
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13920 23075 13923
rect 23124 13920 23152 14019
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 26142 14016 26148 14068
rect 26200 14056 26206 14068
rect 26237 14059 26295 14065
rect 26237 14056 26249 14059
rect 26200 14028 26249 14056
rect 26200 14016 26206 14028
rect 26237 14025 26249 14028
rect 26283 14025 26295 14059
rect 26237 14019 26295 14025
rect 26605 14059 26663 14065
rect 26605 14025 26617 14059
rect 26651 14025 26663 14059
rect 26605 14019 26663 14025
rect 23566 13988 23572 14000
rect 23063 13892 23152 13920
rect 23400 13960 23572 13988
rect 23063 13889 23075 13892
rect 23017 13883 23075 13889
rect 7892 13824 8064 13852
rect 9861 13855 9919 13861
rect 7892 13812 7898 13824
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10318 13852 10324 13864
rect 9907 13824 10324 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 10468 13824 10609 13852
rect 10468 13812 10474 13824
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 18690 13812 18696 13864
rect 18748 13812 18754 13864
rect 21450 13812 21456 13864
rect 21508 13812 21514 13864
rect 23400 13852 23428 13960
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 24302 13988 24308 14000
rect 23900 13960 24308 13988
rect 23900 13948 23906 13960
rect 24302 13948 24308 13960
rect 24360 13988 24366 14000
rect 24360 13960 25544 13988
rect 24360 13948 24366 13960
rect 21560 13824 23428 13852
rect 23492 13892 23796 13920
rect 19150 13784 19156 13796
rect 17880 13756 19156 13784
rect 17880 13728 17908 13756
rect 19150 13744 19156 13756
rect 19208 13784 19214 13796
rect 21560 13784 21588 13824
rect 19208 13756 19472 13784
rect 19208 13744 19214 13756
rect 6822 13676 6828 13728
rect 6880 13676 6886 13728
rect 6914 13676 6920 13728
rect 6972 13676 6978 13728
rect 8481 13719 8539 13725
rect 8481 13685 8493 13719
rect 8527 13716 8539 13719
rect 8846 13716 8852 13728
rect 8527 13688 8852 13716
rect 8527 13685 8539 13688
rect 8481 13679 8539 13685
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 13262 13716 13268 13728
rect 12308 13688 13268 13716
rect 12308 13676 12314 13688
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 17313 13719 17371 13725
rect 17313 13685 17325 13719
rect 17359 13716 17371 13719
rect 17402 13716 17408 13728
rect 17359 13688 17408 13716
rect 17359 13685 17371 13688
rect 17313 13679 17371 13685
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17862 13676 17868 13728
rect 17920 13676 17926 13728
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 19058 13716 19064 13728
rect 18012 13688 19064 13716
rect 18012 13676 18018 13688
rect 19058 13676 19064 13688
rect 19116 13676 19122 13728
rect 19444 13716 19472 13756
rect 20456 13756 21588 13784
rect 20456 13728 20484 13756
rect 21910 13744 21916 13796
rect 21968 13784 21974 13796
rect 23492 13784 23520 13892
rect 23569 13855 23627 13861
rect 23569 13821 23581 13855
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 21968 13756 23520 13784
rect 21968 13744 21974 13756
rect 20438 13716 20444 13728
rect 19444 13688 20444 13716
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 20898 13676 20904 13728
rect 20956 13676 20962 13728
rect 22373 13719 22431 13725
rect 22373 13685 22385 13719
rect 22419 13716 22431 13719
rect 22462 13716 22468 13728
rect 22419 13688 22468 13716
rect 22419 13685 22431 13688
rect 22373 13679 22431 13685
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 23584 13716 23612 13815
rect 23658 13812 23664 13864
rect 23716 13812 23722 13864
rect 23768 13784 23796 13892
rect 23934 13812 23940 13864
rect 23992 13812 23998 13864
rect 25130 13812 25136 13864
rect 25188 13812 25194 13864
rect 25516 13852 25544 13960
rect 25608 13920 25636 14016
rect 25685 13923 25743 13929
rect 25685 13920 25697 13923
rect 25608 13892 25697 13920
rect 25685 13889 25697 13892
rect 25731 13889 25743 13923
rect 25866 13920 25872 13932
rect 25685 13883 25743 13889
rect 25792 13892 25872 13920
rect 25792 13852 25820 13892
rect 25866 13880 25872 13892
rect 25924 13920 25930 13932
rect 26620 13920 26648 14019
rect 29730 14016 29736 14068
rect 29788 14056 29794 14068
rect 29825 14059 29883 14065
rect 29825 14056 29837 14059
rect 29788 14028 29837 14056
rect 29788 14016 29794 14028
rect 29825 14025 29837 14028
rect 29871 14025 29883 14059
rect 30650 14056 30656 14068
rect 29825 14019 29883 14025
rect 30116 14028 30656 14056
rect 28718 13997 28724 14000
rect 28712 13988 28724 13997
rect 28679 13960 28724 13988
rect 28712 13951 28724 13960
rect 28718 13948 28724 13951
rect 28776 13948 28782 14000
rect 30116 13929 30144 14028
rect 30650 14016 30656 14028
rect 30708 14016 30714 14068
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 31941 14059 31999 14065
rect 30892 14028 31800 14056
rect 30892 14016 30898 14028
rect 31772 13988 31800 14028
rect 31941 14025 31953 14059
rect 31987 14056 31999 14059
rect 32490 14056 32496 14068
rect 31987 14028 32496 14056
rect 31987 14025 31999 14028
rect 31941 14019 31999 14025
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 33410 14056 33416 14068
rect 32600 14028 33416 14056
rect 32122 13988 32128 14000
rect 31772 13960 32128 13988
rect 32122 13948 32128 13960
rect 32180 13988 32186 14000
rect 32600 13988 32628 14028
rect 33410 14016 33416 14028
rect 33468 14016 33474 14068
rect 33502 14016 33508 14068
rect 33560 14016 33566 14068
rect 33594 14016 33600 14068
rect 33652 14016 33658 14068
rect 35894 14016 35900 14068
rect 35952 14016 35958 14068
rect 35986 14016 35992 14068
rect 36044 14016 36050 14068
rect 36081 14059 36139 14065
rect 36081 14025 36093 14059
rect 36127 14056 36139 14059
rect 36722 14056 36728 14068
rect 36127 14028 36728 14056
rect 36127 14025 36139 14028
rect 36081 14019 36139 14025
rect 36722 14016 36728 14028
rect 36780 14016 36786 14068
rect 38194 14056 38200 14068
rect 37476 14028 38200 14056
rect 32180 13960 32628 13988
rect 33260 13991 33318 13997
rect 32180 13948 32186 13960
rect 33260 13957 33272 13991
rect 33306 13988 33318 13991
rect 33520 13988 33548 14016
rect 33306 13960 33548 13988
rect 33306 13957 33318 13960
rect 33260 13951 33318 13957
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 25924 13892 26188 13920
rect 26620 13892 27169 13920
rect 25924 13880 25930 13892
rect 26160 13861 26188 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 30101 13923 30159 13929
rect 30101 13889 30113 13923
rect 30147 13889 30159 13923
rect 30101 13883 30159 13889
rect 30285 13923 30343 13929
rect 30285 13889 30297 13923
rect 30331 13889 30343 13923
rect 30285 13883 30343 13889
rect 25516 13824 25820 13852
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13821 26019 13855
rect 25961 13815 26019 13821
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 27246 13852 27252 13864
rect 26191 13824 27252 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 24949 13787 25007 13793
rect 24949 13784 24961 13787
rect 23768 13756 24961 13784
rect 24949 13753 24961 13756
rect 24995 13784 25007 13787
rect 25976 13784 26004 13815
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 28445 13855 28503 13861
rect 28445 13852 28457 13855
rect 28092 13824 28457 13852
rect 24995 13756 26004 13784
rect 24995 13753 25007 13756
rect 24949 13747 25007 13753
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 27614 13784 27620 13796
rect 26292 13756 27620 13784
rect 26292 13744 26298 13756
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 28092 13728 28120 13824
rect 28445 13821 28457 13824
rect 28491 13821 28503 13855
rect 30300 13852 30328 13883
rect 31018 13880 31024 13932
rect 31076 13880 31082 13932
rect 33505 13923 33563 13929
rect 32140 13892 33456 13920
rect 30834 13852 30840 13864
rect 30300 13824 30840 13852
rect 28445 13815 28503 13821
rect 30834 13812 30840 13824
rect 30892 13812 30898 13864
rect 31110 13812 31116 13864
rect 31168 13861 31174 13864
rect 31168 13855 31196 13861
rect 31184 13821 31196 13855
rect 31168 13815 31196 13821
rect 31297 13855 31355 13861
rect 31297 13821 31309 13855
rect 31343 13852 31355 13855
rect 32030 13852 32036 13864
rect 31343 13824 32036 13852
rect 31343 13821 31355 13824
rect 31297 13815 31355 13821
rect 31168 13812 31174 13815
rect 32030 13812 32036 13824
rect 32088 13812 32094 13864
rect 30466 13744 30472 13796
rect 30524 13784 30530 13796
rect 32140 13793 32168 13892
rect 33428 13852 33456 13892
rect 33505 13889 33517 13923
rect 33551 13920 33563 13923
rect 33612 13920 33640 14016
rect 34876 13991 34934 13997
rect 34876 13957 34888 13991
rect 34922 13988 34934 13991
rect 35912 13988 35940 14016
rect 34922 13960 35940 13988
rect 36541 13991 36599 13997
rect 34922 13957 34934 13960
rect 34876 13951 34934 13957
rect 36541 13957 36553 13991
rect 36587 13988 36599 13991
rect 37476 13988 37504 14028
rect 38194 14016 38200 14028
rect 38252 14016 38258 14068
rect 38930 14016 38936 14068
rect 38988 14056 38994 14068
rect 39485 14059 39543 14065
rect 39485 14056 39497 14059
rect 38988 14028 39497 14056
rect 38988 14016 38994 14028
rect 39485 14025 39497 14028
rect 39531 14025 39543 14059
rect 39485 14019 39543 14025
rect 39945 14059 40003 14065
rect 39945 14025 39957 14059
rect 39991 14056 40003 14059
rect 40218 14056 40224 14068
rect 39991 14028 40224 14056
rect 39991 14025 40003 14028
rect 39945 14019 40003 14025
rect 40218 14016 40224 14028
rect 40276 14016 40282 14068
rect 40405 14059 40463 14065
rect 40405 14025 40417 14059
rect 40451 14056 40463 14059
rect 40862 14056 40868 14068
rect 40451 14028 40868 14056
rect 40451 14025 40463 14028
rect 40405 14019 40463 14025
rect 40862 14016 40868 14028
rect 40920 14016 40926 14068
rect 42245 14059 42303 14065
rect 42245 14025 42257 14059
rect 42291 14056 42303 14059
rect 43530 14056 43536 14068
rect 42291 14028 43536 14056
rect 42291 14025 42303 14028
rect 42245 14019 42303 14025
rect 43530 14016 43536 14028
rect 43588 14016 43594 14068
rect 43622 14016 43628 14068
rect 43680 14056 43686 14068
rect 45002 14056 45008 14068
rect 43680 14028 45008 14056
rect 43680 14016 43686 14028
rect 45002 14016 45008 14028
rect 45060 14016 45066 14068
rect 45462 14016 45468 14068
rect 45520 14016 45526 14068
rect 45738 14016 45744 14068
rect 45796 14016 45802 14068
rect 46661 14059 46719 14065
rect 46661 14025 46673 14059
rect 46707 14056 46719 14059
rect 47026 14056 47032 14068
rect 46707 14028 47032 14056
rect 46707 14025 46719 14028
rect 46661 14019 46719 14025
rect 47026 14016 47032 14028
rect 47084 14016 47090 14068
rect 48314 14016 48320 14068
rect 48372 14016 48378 14068
rect 49329 14059 49387 14065
rect 49329 14025 49341 14059
rect 49375 14056 49387 14059
rect 49510 14056 49516 14068
rect 49375 14028 49516 14056
rect 49375 14025 49387 14028
rect 49329 14019 49387 14025
rect 49510 14016 49516 14028
rect 49568 14016 49574 14068
rect 50801 14059 50859 14065
rect 50801 14025 50813 14059
rect 50847 14025 50859 14059
rect 50801 14019 50859 14025
rect 36587 13960 37504 13988
rect 36587 13957 36599 13960
rect 36541 13951 36599 13957
rect 40034 13948 40040 14000
rect 40092 13988 40098 14000
rect 41138 13997 41144 14000
rect 41121 13991 41144 13997
rect 40092 13960 40724 13988
rect 40092 13948 40098 13960
rect 34606 13920 34612 13932
rect 33551 13892 34612 13920
rect 33551 13889 33563 13892
rect 33505 13883 33563 13889
rect 34606 13880 34612 13892
rect 34664 13880 34670 13932
rect 36449 13923 36507 13929
rect 36449 13889 36461 13923
rect 36495 13920 36507 13923
rect 37182 13920 37188 13932
rect 36495 13892 37188 13920
rect 36495 13889 36507 13892
rect 36449 13883 36507 13889
rect 37182 13880 37188 13892
rect 37240 13880 37246 13932
rect 37277 13923 37335 13929
rect 37277 13889 37289 13923
rect 37323 13920 37335 13923
rect 37366 13920 37372 13932
rect 37323 13892 37372 13920
rect 37323 13889 37335 13892
rect 37277 13883 37335 13889
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 37642 13880 37648 13932
rect 37700 13880 37706 13932
rect 38194 13880 38200 13932
rect 38252 13880 38258 13932
rect 38473 13923 38531 13929
rect 38473 13889 38485 13923
rect 38519 13889 38531 13923
rect 38473 13883 38531 13889
rect 39117 13923 39175 13929
rect 39117 13889 39129 13923
rect 39163 13920 39175 13923
rect 39577 13923 39635 13929
rect 39577 13920 39589 13923
rect 39163 13892 39589 13920
rect 39163 13889 39175 13892
rect 39117 13883 39175 13889
rect 39577 13889 39589 13892
rect 39623 13889 39635 13923
rect 39577 13883 39635 13889
rect 34149 13855 34207 13861
rect 34149 13852 34161 13855
rect 33428 13824 34161 13852
rect 34149 13821 34161 13824
rect 34195 13821 34207 13855
rect 34149 13815 34207 13821
rect 36538 13812 36544 13864
rect 36596 13852 36602 13864
rect 36633 13855 36691 13861
rect 36633 13852 36645 13855
rect 36596 13824 36645 13852
rect 36596 13812 36602 13824
rect 36633 13821 36645 13824
rect 36679 13821 36691 13855
rect 36633 13815 36691 13821
rect 36722 13812 36728 13864
rect 36780 13852 36786 13864
rect 37461 13855 37519 13861
rect 36780 13824 37412 13852
rect 36780 13812 36786 13824
rect 30745 13787 30803 13793
rect 30745 13784 30757 13787
rect 30524 13756 30757 13784
rect 30524 13744 30530 13756
rect 30745 13753 30757 13756
rect 30791 13753 30803 13787
rect 30745 13747 30803 13753
rect 32125 13787 32183 13793
rect 32125 13753 32137 13787
rect 32171 13753 32183 13787
rect 37384 13784 37412 13824
rect 37461 13821 37473 13855
rect 37507 13852 37519 13855
rect 37660 13852 37688 13880
rect 38335 13855 38393 13861
rect 38335 13852 38347 13855
rect 37507 13824 37688 13852
rect 37752 13824 38347 13852
rect 37507 13821 37519 13824
rect 37461 13815 37519 13821
rect 37752 13784 37780 13824
rect 38335 13821 38347 13824
rect 38381 13821 38393 13855
rect 38488 13852 38516 13883
rect 38654 13852 38660 13864
rect 38488 13824 38660 13852
rect 38335 13815 38393 13821
rect 38654 13812 38660 13824
rect 38712 13812 38718 13864
rect 39390 13812 39396 13864
rect 39448 13812 39454 13864
rect 39758 13812 39764 13864
rect 39816 13812 39822 13864
rect 40494 13812 40500 13864
rect 40552 13812 40558 13864
rect 40696 13861 40724 13960
rect 41121 13957 41133 13991
rect 41121 13951 41144 13957
rect 41138 13948 41144 13951
rect 41196 13948 41202 14000
rect 44729 13991 44787 13997
rect 44729 13957 44741 13991
rect 44775 13988 44787 13991
rect 45480 13988 45508 14016
rect 44775 13960 45508 13988
rect 45756 13988 45784 14016
rect 45756 13960 46612 13988
rect 44775 13957 44787 13960
rect 44729 13951 44787 13957
rect 43806 13880 43812 13932
rect 43864 13880 43870 13932
rect 43898 13880 43904 13932
rect 43956 13929 43962 13932
rect 43956 13923 43984 13929
rect 43972 13889 43984 13923
rect 43956 13883 43984 13889
rect 43956 13880 43962 13883
rect 44082 13880 44088 13932
rect 44140 13880 44146 13932
rect 45281 13923 45339 13929
rect 45281 13889 45293 13923
rect 45327 13920 45339 13923
rect 45370 13920 45376 13932
rect 45327 13892 45376 13920
rect 45327 13889 45339 13892
rect 45281 13883 45339 13889
rect 45370 13880 45376 13892
rect 45428 13880 45434 13932
rect 45548 13923 45606 13929
rect 45548 13889 45560 13923
rect 45594 13920 45606 13923
rect 45830 13920 45836 13932
rect 45594 13892 45836 13920
rect 45594 13889 45606 13892
rect 45548 13883 45606 13889
rect 45830 13880 45836 13892
rect 45888 13880 45894 13932
rect 46584 13920 46612 13960
rect 47302 13948 47308 14000
rect 47360 13988 47366 14000
rect 49970 13988 49976 14000
rect 47360 13960 49976 13988
rect 47360 13948 47366 13960
rect 47397 13923 47455 13929
rect 47397 13920 47409 13923
rect 46584 13892 47409 13920
rect 47397 13889 47409 13892
rect 47443 13889 47455 13923
rect 47397 13883 47455 13889
rect 48866 13880 48872 13932
rect 48924 13880 48930 13932
rect 49436 13929 49464 13960
rect 49970 13948 49976 13960
rect 50028 13948 50034 14000
rect 50430 13948 50436 14000
rect 50488 13948 50494 14000
rect 49421 13923 49479 13929
rect 49421 13889 49433 13923
rect 49467 13889 49479 13923
rect 49421 13883 49479 13889
rect 49688 13923 49746 13929
rect 49688 13889 49700 13923
rect 49734 13920 49746 13923
rect 50448 13920 50476 13948
rect 49734 13892 50476 13920
rect 50816 13920 50844 14019
rect 50890 14016 50896 14068
rect 50948 14056 50954 14068
rect 51537 14059 51595 14065
rect 51537 14056 51549 14059
rect 50948 14028 51549 14056
rect 50948 14016 50954 14028
rect 51537 14025 51549 14028
rect 51583 14056 51595 14059
rect 51994 14056 52000 14068
rect 51583 14028 52000 14056
rect 51583 14025 51595 14028
rect 51537 14019 51595 14025
rect 51994 14016 52000 14028
rect 52052 14016 52058 14068
rect 54481 14059 54539 14065
rect 54481 14025 54493 14059
rect 54527 14056 54539 14059
rect 55214 14056 55220 14068
rect 54527 14028 55220 14056
rect 54527 14025 54539 14028
rect 54481 14019 54539 14025
rect 55214 14016 55220 14028
rect 55272 14016 55278 14068
rect 56045 14059 56103 14065
rect 56045 14025 56057 14059
rect 56091 14056 56103 14059
rect 57517 14059 57575 14065
rect 56091 14028 56272 14056
rect 56091 14025 56103 14028
rect 56045 14019 56103 14025
rect 56244 13988 56272 14028
rect 57517 14025 57529 14059
rect 57563 14056 57575 14059
rect 58434 14056 58440 14068
rect 57563 14028 58440 14056
rect 57563 14025 57575 14028
rect 57517 14019 57575 14025
rect 58434 14016 58440 14028
rect 58492 14016 58498 14068
rect 56382 13991 56440 13997
rect 56382 13988 56394 13991
rect 56244 13960 56394 13988
rect 56382 13957 56394 13960
rect 56428 13957 56440 13991
rect 56382 13951 56440 13957
rect 57698 13948 57704 14000
rect 57756 13948 57762 14000
rect 57882 13948 57888 14000
rect 57940 13948 57946 14000
rect 50893 13923 50951 13929
rect 50893 13920 50905 13923
rect 50816 13892 50905 13920
rect 49734 13889 49746 13892
rect 49688 13883 49746 13889
rect 50893 13889 50905 13892
rect 50939 13889 50951 13923
rect 50893 13883 50951 13889
rect 51902 13880 51908 13932
rect 51960 13920 51966 13932
rect 52181 13923 52239 13929
rect 52181 13920 52193 13923
rect 51960 13892 52193 13920
rect 51960 13880 51966 13892
rect 52181 13889 52193 13892
rect 52227 13889 52239 13923
rect 52181 13883 52239 13889
rect 53368 13923 53426 13929
rect 53368 13889 53380 13923
rect 53414 13920 53426 13923
rect 54294 13920 54300 13932
rect 53414 13892 54300 13920
rect 53414 13889 53426 13892
rect 53368 13883 53426 13889
rect 54294 13880 54300 13892
rect 54352 13880 54358 13932
rect 54938 13880 54944 13932
rect 54996 13880 55002 13932
rect 57716 13920 57744 13948
rect 58437 13923 58495 13929
rect 58437 13920 58449 13923
rect 57716 13892 58449 13920
rect 58437 13889 58449 13892
rect 58483 13889 58495 13923
rect 58437 13883 58495 13889
rect 40681 13855 40739 13861
rect 40681 13821 40693 13855
rect 40727 13821 40739 13855
rect 40681 13815 40739 13821
rect 40865 13855 40923 13861
rect 40865 13821 40877 13855
rect 40911 13821 40923 13855
rect 40865 13815 40923 13821
rect 32125 13747 32183 13753
rect 33520 13756 33732 13784
rect 23842 13716 23848 13728
rect 23584 13688 23848 13716
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 27706 13676 27712 13728
rect 27764 13716 27770 13728
rect 27801 13719 27859 13725
rect 27801 13716 27813 13719
rect 27764 13688 27813 13716
rect 27764 13676 27770 13688
rect 27801 13685 27813 13688
rect 27847 13685 27859 13719
rect 27801 13679 27859 13685
rect 28074 13676 28080 13728
rect 28132 13676 28138 13728
rect 29914 13676 29920 13728
rect 29972 13716 29978 13728
rect 33520 13716 33548 13756
rect 29972 13688 33548 13716
rect 29972 13676 29978 13688
rect 33594 13676 33600 13728
rect 33652 13676 33658 13728
rect 33704 13716 33732 13756
rect 35912 13756 36124 13784
rect 37384 13756 37780 13784
rect 35912 13716 35940 13756
rect 33704 13688 35940 13716
rect 36096 13716 36124 13756
rect 37826 13744 37832 13796
rect 37884 13784 37890 13796
rect 37921 13787 37979 13793
rect 37921 13784 37933 13787
rect 37884 13756 37933 13784
rect 37884 13744 37890 13756
rect 37921 13753 37933 13756
rect 37967 13753 37979 13787
rect 39776 13784 39804 13812
rect 40880 13784 40908 13815
rect 42702 13812 42708 13864
rect 42760 13812 42766 13864
rect 42889 13855 42947 13861
rect 42889 13821 42901 13855
rect 42935 13852 42947 13855
rect 42978 13852 42984 13864
rect 42935 13824 42984 13852
rect 42935 13821 42947 13824
rect 42889 13815 42947 13821
rect 42978 13812 42984 13824
rect 43036 13812 43042 13864
rect 43073 13855 43131 13861
rect 43073 13821 43085 13855
rect 43119 13852 43131 13855
rect 45002 13852 45008 13864
rect 43119 13824 45008 13852
rect 43119 13821 43131 13824
rect 43073 13815 43131 13821
rect 45002 13812 45008 13824
rect 45060 13812 45066 13864
rect 51074 13812 51080 13864
rect 51132 13852 51138 13864
rect 51629 13855 51687 13861
rect 51629 13852 51641 13855
rect 51132 13824 51641 13852
rect 51132 13812 51138 13824
rect 51629 13821 51641 13824
rect 51675 13821 51687 13855
rect 51629 13815 51687 13821
rect 51994 13812 52000 13864
rect 52052 13852 52058 13864
rect 52270 13852 52276 13864
rect 52052 13824 52276 13852
rect 52052 13812 52058 13824
rect 52270 13812 52276 13824
rect 52328 13812 52334 13864
rect 53006 13812 53012 13864
rect 53064 13852 53070 13864
rect 53101 13855 53159 13861
rect 53101 13852 53113 13855
rect 53064 13824 53113 13852
rect 53064 13812 53070 13824
rect 53101 13821 53113 13824
rect 53147 13821 53159 13855
rect 53101 13815 53159 13821
rect 39776 13756 40908 13784
rect 37921 13747 37979 13753
rect 39942 13716 39948 13728
rect 36096 13688 39948 13716
rect 39942 13676 39948 13688
rect 40000 13676 40006 13728
rect 40034 13676 40040 13728
rect 40092 13676 40098 13728
rect 40880 13716 40908 13756
rect 43533 13787 43591 13793
rect 43533 13753 43545 13787
rect 43579 13784 43591 13787
rect 43622 13784 43628 13796
rect 43579 13756 43628 13784
rect 43579 13753 43591 13756
rect 43533 13747 43591 13753
rect 43622 13744 43628 13756
rect 43680 13744 43686 13796
rect 41598 13716 41604 13728
rect 40880 13688 41604 13716
rect 41598 13676 41604 13688
rect 41656 13676 41662 13728
rect 44082 13676 44088 13728
rect 44140 13716 44146 13728
rect 45005 13719 45063 13725
rect 45005 13716 45017 13719
rect 44140 13688 45017 13716
rect 44140 13676 44146 13688
rect 45005 13685 45017 13688
rect 45051 13716 45063 13719
rect 46566 13716 46572 13728
rect 45051 13688 46572 13716
rect 45051 13685 45063 13688
rect 45005 13679 45063 13685
rect 46566 13676 46572 13688
rect 46624 13676 46630 13728
rect 46750 13676 46756 13728
rect 46808 13676 46814 13728
rect 50430 13676 50436 13728
rect 50488 13716 50494 13728
rect 51258 13716 51264 13728
rect 50488 13688 51264 13716
rect 50488 13676 50494 13688
rect 51258 13676 51264 13688
rect 51316 13676 51322 13728
rect 53009 13719 53067 13725
rect 53009 13685 53021 13719
rect 53055 13716 53067 13719
rect 53116 13716 53144 13815
rect 55490 13812 55496 13864
rect 55548 13812 55554 13864
rect 56134 13812 56140 13864
rect 56192 13812 56198 13864
rect 56152 13716 56180 13812
rect 53055 13688 56180 13716
rect 53055 13685 53067 13688
rect 53009 13679 53067 13685
rect 1104 13626 58880 13648
rect 1104 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 22616 13626
rect 22668 13574 22680 13626
rect 22732 13574 22744 13626
rect 22796 13574 22808 13626
rect 22860 13574 22872 13626
rect 22924 13574 37060 13626
rect 37112 13574 37124 13626
rect 37176 13574 37188 13626
rect 37240 13574 37252 13626
rect 37304 13574 37316 13626
rect 37368 13574 51504 13626
rect 51556 13574 51568 13626
rect 51620 13574 51632 13626
rect 51684 13574 51696 13626
rect 51748 13574 51760 13626
rect 51812 13574 58880 13626
rect 1104 13552 58880 13574
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10870 13512 10876 13524
rect 10091 13484 10876 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13320 13484 18368 13512
rect 13320 13472 13326 13484
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 15657 13447 15715 13453
rect 15657 13413 15669 13447
rect 15703 13444 15715 13447
rect 17034 13444 17040 13456
rect 15703 13416 17040 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 7392 13376 7420 13407
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7392 13348 7481 13376
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 8904 13348 9413 13376
rect 8904 13336 8910 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 10686 13336 10692 13388
rect 10744 13336 10750 13388
rect 12986 13336 12992 13388
rect 13044 13336 13050 13388
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13376 13967 13379
rect 14737 13379 14795 13385
rect 14737 13376 14749 13379
rect 13955 13348 14749 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 14737 13345 14749 13348
rect 14783 13376 14795 13379
rect 14918 13376 14924 13388
rect 14783 13348 14924 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 3510 13268 3516 13320
rect 3568 13268 3574 13320
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 3936 13280 4261 13308
rect 3936 13268 3942 13280
rect 4249 13277 4261 13280
rect 4295 13308 4307 13311
rect 5994 13308 6000 13320
rect 4295 13280 6000 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5994 13268 6000 13280
rect 6052 13308 6058 13320
rect 6822 13308 6828 13320
rect 6052 13280 6828 13308
rect 6052 13268 6058 13280
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 13924 13308 13952 13339
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 16408 13385 16436 13416
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 16080 13348 16221 13376
rect 16080 13336 16086 13348
rect 16209 13345 16221 13348
rect 16255 13345 16267 13379
rect 16209 13339 16267 13345
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 16439 13348 16473 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 17310 13336 17316 13388
rect 17368 13336 17374 13388
rect 18340 13376 18368 13484
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18564 13484 18705 13512
rect 18564 13472 18570 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18693 13475 18751 13481
rect 19245 13515 19303 13521
rect 19245 13481 19257 13515
rect 19291 13512 19303 13515
rect 20162 13512 20168 13524
rect 19291 13484 20168 13512
rect 19291 13481 19303 13484
rect 19245 13475 19303 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 21177 13515 21235 13521
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 21450 13512 21456 13524
rect 21223 13484 21456 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 23845 13515 23903 13521
rect 22066 13484 23428 13512
rect 22066 13444 22094 13484
rect 20364 13416 22094 13444
rect 20364 13376 20392 13416
rect 22462 13404 22468 13456
rect 22520 13404 22526 13456
rect 23400 13444 23428 13484
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 23934 13512 23940 13524
rect 23891 13484 23940 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24780 13484 25636 13512
rect 24780 13444 24808 13484
rect 23400 13416 24808 13444
rect 25608 13444 25636 13484
rect 26418 13472 26424 13524
rect 26476 13472 26482 13524
rect 29914 13512 29920 13524
rect 26896 13484 29920 13512
rect 26896 13444 26924 13484
rect 29914 13472 29920 13484
rect 29972 13472 29978 13524
rect 30374 13472 30380 13524
rect 30432 13512 30438 13524
rect 31478 13512 31484 13524
rect 30432 13484 31484 13512
rect 30432 13472 30438 13484
rect 31478 13472 31484 13484
rect 31536 13512 31542 13524
rect 31536 13484 39896 13512
rect 31536 13472 31542 13484
rect 25608 13416 26924 13444
rect 31021 13447 31079 13453
rect 31021 13413 31033 13447
rect 31067 13444 31079 13447
rect 31202 13444 31208 13456
rect 31067 13416 31208 13444
rect 31067 13413 31079 13416
rect 31021 13407 31079 13413
rect 31202 13404 31208 13416
rect 31260 13404 31266 13456
rect 32398 13404 32404 13456
rect 32456 13444 32462 13456
rect 32493 13447 32551 13453
rect 32493 13444 32505 13447
rect 32456 13416 32505 13444
rect 32456 13404 32462 13416
rect 32493 13413 32505 13416
rect 32539 13413 32551 13447
rect 32493 13407 32551 13413
rect 33965 13447 34023 13453
rect 33965 13413 33977 13447
rect 34011 13444 34023 13447
rect 34514 13444 34520 13456
rect 34011 13416 34520 13444
rect 34011 13413 34023 13416
rect 33965 13407 34023 13413
rect 34514 13404 34520 13416
rect 34572 13404 34578 13456
rect 18340 13348 20392 13376
rect 20438 13336 20444 13388
rect 20496 13336 20502 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 21821 13379 21879 13385
rect 20772 13348 21680 13376
rect 20772 13336 20778 13348
rect 12400 13280 13952 13308
rect 14553 13311 14611 13317
rect 12400 13268 12406 13280
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 15838 13308 15844 13320
rect 14599 13280 15844 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 16114 13268 16120 13320
rect 16172 13268 16178 13320
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17569 13311 17627 13317
rect 17569 13308 17581 13311
rect 17460 13280 17581 13308
rect 17460 13268 17466 13280
rect 17569 13277 17581 13280
rect 17615 13277 17627 13311
rect 17569 13271 17627 13277
rect 19058 13268 19064 13320
rect 19116 13268 19122 13320
rect 19886 13268 19892 13320
rect 19944 13268 19950 13320
rect 20070 13317 20076 13320
rect 20048 13311 20076 13317
rect 20048 13277 20060 13311
rect 20048 13271 20076 13277
rect 20070 13268 20076 13271
rect 20128 13268 20134 13320
rect 20162 13268 20168 13320
rect 20220 13268 20226 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 6264 13243 6322 13249
rect 6264 13209 6276 13243
rect 6310 13240 6322 13243
rect 6454 13240 6460 13252
rect 6310 13212 6460 13240
rect 6310 13209 6322 13212
rect 6264 13203 6322 13209
rect 6454 13200 6460 13212
rect 6512 13200 6518 13252
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 9217 13243 9275 13249
rect 9217 13240 9229 13243
rect 8812 13212 9229 13240
rect 8812 13200 8818 13212
rect 9217 13209 9229 13212
rect 9263 13240 9275 13243
rect 9263 13212 10916 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 10888 13184 10916 13212
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 13964 13212 14473 13240
rect 13964 13200 13970 13212
rect 14461 13209 14473 13212
rect 14507 13209 14519 13243
rect 14461 13203 14519 13209
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 15197 13243 15255 13249
rect 15197 13240 15209 13243
rect 15160 13212 15209 13240
rect 15160 13200 15166 13212
rect 15197 13209 15209 13212
rect 15243 13240 15255 13243
rect 15243 13212 16804 13240
rect 15243 13209 15255 13212
rect 15197 13203 15255 13209
rect 16776 13184 16804 13212
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 18414 13240 18420 13252
rect 17092 13212 18420 13240
rect 17092 13200 17098 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 19076 13240 19104 13268
rect 20916 13240 20944 13271
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21358 13308 21364 13320
rect 21140 13280 21364 13308
rect 21140 13268 21146 13280
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21652 13317 21680 13348
rect 21821 13345 21833 13379
rect 21867 13376 21879 13379
rect 21867 13348 21956 13376
rect 21867 13345 21879 13348
rect 21821 13339 21879 13345
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 21450 13240 21456 13252
rect 19076 13212 19334 13240
rect 20916 13212 21456 13240
rect 2958 13132 2964 13184
rect 3016 13132 3022 13184
rect 8110 13132 8116 13184
rect 8168 13132 8174 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 13630 13172 13636 13184
rect 13495 13144 13636 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14366 13172 14372 13184
rect 14139 13144 14372 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 16022 13172 16028 13184
rect 15896 13144 16028 13172
rect 15896 13132 15902 13144
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16758 13132 16764 13184
rect 16816 13132 16822 13184
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17862 13172 17868 13184
rect 17276 13144 17868 13172
rect 17276 13132 17282 13144
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 19058 13132 19064 13184
rect 19116 13132 19122 13184
rect 19306 13172 19334 13212
rect 21450 13200 21456 13212
rect 21508 13200 21514 13252
rect 21928 13184 21956 13348
rect 22370 13336 22376 13388
rect 22428 13336 22434 13388
rect 22480 13376 22508 13404
rect 24213 13379 24271 13385
rect 22480 13348 22600 13376
rect 22388 13308 22416 13336
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22388 13280 22477 13308
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22572 13308 22600 13348
rect 24213 13345 24225 13379
rect 24259 13376 24271 13379
rect 24762 13376 24768 13388
rect 24259 13348 24768 13376
rect 24259 13345 24271 13348
rect 24213 13339 24271 13345
rect 24762 13336 24768 13348
rect 24820 13376 24826 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 24820 13348 25145 13376
rect 24820 13336 24826 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 25409 13379 25467 13385
rect 25409 13345 25421 13379
rect 25455 13376 25467 13379
rect 25590 13376 25596 13388
rect 25455 13348 25596 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 25590 13336 25596 13348
rect 25648 13336 25654 13388
rect 25685 13379 25743 13385
rect 25685 13345 25697 13379
rect 25731 13376 25743 13379
rect 25774 13376 25780 13388
rect 25731 13348 25780 13376
rect 25731 13345 25743 13348
rect 25685 13339 25743 13345
rect 25774 13336 25780 13348
rect 25832 13336 25838 13388
rect 26142 13336 26148 13388
rect 26200 13336 26206 13388
rect 31941 13379 31999 13385
rect 31941 13345 31953 13379
rect 31987 13376 31999 13379
rect 31987 13348 32720 13376
rect 31987 13345 31999 13348
rect 31941 13339 31999 13345
rect 25314 13317 25320 13320
rect 22721 13311 22779 13317
rect 22721 13308 22733 13311
rect 22572 13280 22733 13308
rect 22465 13271 22523 13277
rect 22721 13277 22733 13280
rect 22767 13277 22779 13311
rect 22721 13271 22779 13277
rect 25292 13311 25320 13317
rect 25292 13277 25304 13311
rect 25292 13271 25320 13277
rect 25314 13268 25320 13271
rect 25372 13268 25378 13320
rect 26234 13268 26240 13320
rect 26292 13308 26298 13320
rect 26329 13311 26387 13317
rect 26329 13308 26341 13311
rect 26292 13280 26341 13308
rect 26292 13268 26298 13280
rect 26329 13277 26341 13280
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 27798 13268 27804 13320
rect 27856 13308 27862 13320
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 27856 13280 27997 13308
rect 27856 13268 27862 13280
rect 27985 13277 27997 13280
rect 28031 13308 28043 13311
rect 28074 13308 28080 13320
rect 28031 13280 28080 13308
rect 28031 13277 28043 13280
rect 27985 13271 28043 13277
rect 28074 13268 28080 13280
rect 28132 13308 28138 13320
rect 29641 13311 29699 13317
rect 29641 13308 29653 13311
rect 28132 13280 29653 13308
rect 28132 13268 28138 13280
rect 29641 13277 29653 13280
rect 29687 13308 29699 13311
rect 29730 13308 29736 13320
rect 29687 13280 29736 13308
rect 29687 13277 29699 13280
rect 29641 13271 29699 13277
rect 29730 13268 29736 13280
rect 29788 13308 29794 13320
rect 31389 13311 31447 13317
rect 31389 13308 31401 13311
rect 29788 13280 31401 13308
rect 29788 13268 29794 13280
rect 31389 13277 31401 13280
rect 31435 13308 31447 13311
rect 32585 13311 32643 13317
rect 32585 13308 32597 13311
rect 31435 13280 32597 13308
rect 31435 13277 31447 13280
rect 31389 13271 31447 13277
rect 32585 13277 32597 13280
rect 32631 13277 32643 13311
rect 32692 13308 32720 13348
rect 34606 13336 34612 13388
rect 34664 13376 34670 13388
rect 34701 13379 34759 13385
rect 34701 13376 34713 13379
rect 34664 13348 34713 13376
rect 34664 13336 34670 13348
rect 34701 13345 34713 13348
rect 34747 13345 34759 13379
rect 34701 13339 34759 13345
rect 34716 13308 34744 13339
rect 39868 13320 39896 13484
rect 45830 13472 45836 13524
rect 45888 13472 45894 13524
rect 46661 13515 46719 13521
rect 46661 13512 46673 13515
rect 46023 13484 46673 13512
rect 43073 13447 43131 13453
rect 43073 13413 43085 13447
rect 43119 13444 43131 13447
rect 43346 13444 43352 13456
rect 43119 13416 43352 13444
rect 43119 13413 43131 13416
rect 43073 13407 43131 13413
rect 43346 13404 43352 13416
rect 43404 13404 43410 13456
rect 41598 13336 41604 13388
rect 41656 13376 41662 13388
rect 41693 13379 41751 13385
rect 41693 13376 41705 13379
rect 41656 13348 41705 13376
rect 41656 13336 41662 13348
rect 41693 13345 41705 13348
rect 41739 13345 41751 13379
rect 41693 13339 41751 13345
rect 45186 13336 45192 13388
rect 45244 13336 45250 13388
rect 46023 13376 46051 13484
rect 46661 13481 46673 13484
rect 46707 13481 46719 13515
rect 46661 13475 46719 13481
rect 49694 13472 49700 13524
rect 49752 13472 49758 13524
rect 55490 13472 55496 13524
rect 55548 13472 55554 13524
rect 55582 13472 55588 13524
rect 55640 13472 55646 13524
rect 56045 13515 56103 13521
rect 56045 13481 56057 13515
rect 56091 13512 56103 13515
rect 56134 13512 56140 13524
rect 56091 13484 56140 13512
rect 56091 13481 56103 13484
rect 56045 13475 56103 13481
rect 56134 13472 56140 13484
rect 56192 13472 56198 13524
rect 46198 13404 46204 13456
rect 46256 13444 46262 13456
rect 55508 13444 55536 13472
rect 56229 13447 56287 13453
rect 56229 13444 56241 13447
rect 46256 13416 51074 13444
rect 55508 13416 56241 13444
rect 46256 13404 46262 13416
rect 45480 13348 46051 13376
rect 35802 13308 35808 13320
rect 32692 13280 34376 13308
rect 34716 13280 35808 13308
rect 32585 13271 32643 13277
rect 27556 13243 27614 13249
rect 27556 13209 27568 13243
rect 27602 13240 27614 13243
rect 27706 13240 27712 13252
rect 27602 13212 27712 13240
rect 27602 13209 27614 13212
rect 27556 13203 27614 13209
rect 27706 13200 27712 13212
rect 27764 13200 27770 13252
rect 28252 13243 28310 13249
rect 28252 13209 28264 13243
rect 28298 13240 28310 13243
rect 28626 13240 28632 13252
rect 28298 13212 28632 13240
rect 28298 13209 28310 13212
rect 28252 13203 28310 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 29908 13243 29966 13249
rect 29908 13209 29920 13243
rect 29954 13240 29966 13243
rect 30466 13240 30472 13252
rect 29954 13212 30472 13240
rect 29954 13209 29966 13212
rect 29908 13203 29966 13209
rect 30466 13200 30472 13212
rect 30524 13200 30530 13252
rect 30926 13200 30932 13252
rect 30984 13240 30990 13252
rect 32033 13243 32091 13249
rect 32033 13240 32045 13243
rect 30984 13212 32045 13240
rect 30984 13200 30990 13212
rect 32033 13209 32045 13212
rect 32079 13240 32091 13243
rect 32600 13240 32628 13271
rect 32674 13240 32680 13252
rect 32079 13212 32260 13240
rect 32600 13212 32680 13240
rect 32079 13209 32091 13212
rect 32033 13203 32091 13209
rect 19886 13172 19892 13184
rect 19306 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 21542 13132 21548 13184
rect 21600 13132 21606 13184
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 22189 13175 22247 13181
rect 22189 13172 22201 13175
rect 21968 13144 22201 13172
rect 21968 13132 21974 13144
rect 22189 13141 22201 13144
rect 22235 13141 22247 13175
rect 22189 13135 22247 13141
rect 24489 13175 24547 13181
rect 24489 13141 24501 13175
rect 24535 13172 24547 13175
rect 25682 13172 25688 13184
rect 24535 13144 25688 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 25682 13132 25688 13144
rect 25740 13132 25746 13184
rect 29365 13175 29423 13181
rect 29365 13141 29377 13175
rect 29411 13172 29423 13175
rect 31018 13172 31024 13184
rect 29411 13144 31024 13172
rect 29411 13141 29423 13144
rect 29365 13135 29423 13141
rect 31018 13132 31024 13144
rect 31076 13132 31082 13184
rect 32122 13132 32128 13184
rect 32180 13132 32186 13184
rect 32232 13172 32260 13212
rect 32674 13200 32680 13212
rect 32732 13200 32738 13252
rect 32858 13249 32864 13252
rect 32852 13203 32864 13249
rect 32858 13200 32864 13203
rect 32916 13200 32922 13252
rect 34348 13184 34376 13280
rect 35802 13268 35808 13280
rect 35860 13308 35866 13320
rect 36357 13311 36415 13317
rect 36357 13308 36369 13311
rect 35860 13280 36369 13308
rect 35860 13268 35866 13280
rect 36357 13277 36369 13280
rect 36403 13308 36415 13311
rect 37921 13311 37979 13317
rect 37921 13308 37933 13311
rect 36403 13280 37933 13308
rect 36403 13277 36415 13280
rect 36357 13271 36415 13277
rect 37921 13277 37933 13280
rect 37967 13308 37979 13311
rect 39577 13311 39635 13317
rect 39577 13308 39589 13311
rect 37967 13280 39589 13308
rect 37967 13277 37979 13280
rect 37921 13271 37979 13277
rect 39577 13277 39589 13280
rect 39623 13308 39635 13311
rect 39758 13308 39764 13320
rect 39623 13280 39764 13308
rect 39623 13277 39635 13280
rect 39577 13271 39635 13277
rect 39758 13268 39764 13280
rect 39816 13268 39822 13320
rect 39850 13268 39856 13320
rect 39908 13268 39914 13320
rect 44545 13311 44603 13317
rect 44545 13277 44557 13311
rect 44591 13308 44603 13311
rect 44634 13308 44640 13320
rect 44591 13280 44640 13308
rect 44591 13277 44603 13280
rect 44545 13271 44603 13277
rect 44634 13268 44640 13280
rect 44692 13308 44698 13320
rect 45370 13308 45376 13320
rect 44692 13280 45376 13308
rect 44692 13268 44698 13280
rect 45370 13268 45376 13280
rect 45428 13268 45434 13320
rect 34968 13243 35026 13249
rect 34968 13209 34980 13243
rect 35014 13240 35026 13243
rect 35158 13240 35164 13252
rect 35014 13212 35164 13240
rect 35014 13209 35026 13212
rect 34968 13203 35026 13209
rect 35158 13200 35164 13212
rect 35216 13200 35222 13252
rect 35434 13200 35440 13252
rect 35492 13200 35498 13252
rect 36624 13243 36682 13249
rect 36624 13209 36636 13243
rect 36670 13240 36682 13243
rect 38188 13243 38246 13249
rect 36670 13212 37964 13240
rect 36670 13209 36682 13212
rect 36624 13203 36682 13209
rect 32950 13172 32956 13184
rect 32232 13144 32956 13172
rect 32950 13132 32956 13144
rect 33008 13132 33014 13184
rect 34330 13132 34336 13184
rect 34388 13172 34394 13184
rect 35452 13172 35480 13200
rect 37936 13184 37964 13212
rect 38188 13209 38200 13243
rect 38234 13240 38246 13243
rect 39390 13240 39396 13252
rect 38234 13212 39396 13240
rect 38234 13209 38246 13212
rect 38188 13203 38246 13209
rect 39390 13200 39396 13212
rect 39448 13200 39454 13252
rect 41960 13243 42018 13249
rect 41960 13209 41972 13243
rect 42006 13240 42018 13243
rect 42334 13240 42340 13252
rect 42006 13212 42340 13240
rect 42006 13209 42018 13212
rect 41960 13203 42018 13209
rect 42334 13200 42340 13212
rect 42392 13200 42398 13252
rect 44300 13243 44358 13249
rect 44300 13209 44312 13243
rect 44346 13240 44358 13243
rect 44726 13240 44732 13252
rect 44346 13212 44732 13240
rect 44346 13209 44358 13212
rect 44300 13203 44358 13209
rect 44726 13200 44732 13212
rect 44784 13200 44790 13252
rect 45002 13200 45008 13252
rect 45060 13240 45066 13252
rect 45480 13240 45508 13348
rect 46106 13336 46112 13388
rect 46164 13376 46170 13388
rect 46385 13379 46443 13385
rect 46385 13376 46397 13379
rect 46164 13348 46397 13376
rect 46164 13336 46170 13348
rect 46385 13345 46397 13348
rect 46431 13345 46443 13379
rect 46385 13339 46443 13345
rect 46566 13336 46572 13388
rect 46624 13376 46630 13388
rect 48130 13376 48136 13388
rect 46624 13348 48136 13376
rect 46624 13336 46630 13348
rect 48130 13336 48136 13348
rect 48188 13376 48194 13388
rect 48188 13348 48314 13376
rect 48188 13336 48194 13348
rect 46201 13311 46259 13317
rect 46201 13277 46213 13311
rect 46247 13308 46259 13311
rect 46750 13308 46756 13320
rect 46247 13280 46756 13308
rect 46247 13277 46259 13280
rect 46201 13271 46259 13277
rect 46750 13268 46756 13280
rect 46808 13268 46814 13320
rect 47210 13268 47216 13320
rect 47268 13268 47274 13320
rect 47949 13311 48007 13317
rect 47949 13277 47961 13311
rect 47995 13277 48007 13311
rect 48286 13308 48314 13348
rect 48774 13336 48780 13388
rect 48832 13376 48838 13388
rect 49053 13379 49111 13385
rect 49053 13376 49065 13379
rect 48832 13348 49065 13376
rect 48832 13336 48838 13348
rect 49053 13345 49065 13348
rect 49099 13345 49111 13379
rect 51046 13376 51074 13416
rect 56229 13413 56241 13416
rect 56275 13413 56287 13447
rect 56229 13407 56287 13413
rect 56686 13376 56692 13388
rect 51046 13348 56692 13376
rect 49053 13339 49111 13345
rect 56686 13336 56692 13348
rect 56744 13336 56750 13388
rect 56778 13336 56784 13388
rect 56836 13376 56842 13388
rect 57241 13379 57299 13385
rect 57241 13376 57253 13379
rect 56836 13348 57253 13376
rect 56836 13336 56842 13348
rect 57241 13345 57253 13348
rect 57287 13345 57299 13379
rect 57241 13339 57299 13345
rect 58434 13336 58440 13388
rect 58492 13336 58498 13388
rect 50709 13311 50767 13317
rect 50709 13308 50721 13311
rect 48286 13280 50721 13308
rect 47949 13271 48007 13277
rect 50709 13277 50721 13280
rect 50755 13308 50767 13311
rect 50798 13308 50804 13320
rect 50755 13280 50804 13308
rect 50755 13277 50767 13280
rect 50709 13271 50767 13277
rect 47964 13240 47992 13271
rect 50798 13268 50804 13280
rect 50856 13268 50862 13320
rect 56597 13311 56655 13317
rect 56597 13277 56609 13311
rect 56643 13308 56655 13311
rect 56962 13308 56968 13320
rect 56643 13280 56968 13308
rect 56643 13277 56655 13280
rect 56597 13271 56655 13277
rect 56962 13268 56968 13280
rect 57020 13308 57026 13320
rect 57885 13311 57943 13317
rect 57885 13308 57897 13311
rect 57020 13280 57897 13308
rect 57020 13268 57026 13280
rect 57885 13277 57897 13280
rect 57931 13277 57943 13311
rect 57885 13271 57943 13277
rect 45060 13212 45508 13240
rect 45756 13212 47992 13240
rect 45060 13200 45066 13212
rect 34388 13144 35480 13172
rect 34388 13132 34394 13144
rect 36078 13132 36084 13184
rect 36136 13132 36142 13184
rect 37734 13132 37740 13184
rect 37792 13132 37798 13184
rect 37918 13132 37924 13184
rect 37976 13132 37982 13184
rect 39298 13132 39304 13184
rect 39356 13132 39362 13184
rect 41325 13175 41383 13181
rect 41325 13141 41337 13175
rect 41371 13172 41383 13175
rect 42518 13172 42524 13184
rect 41371 13144 42524 13172
rect 41371 13141 41383 13144
rect 41325 13135 41383 13141
rect 42518 13132 42524 13144
rect 42576 13132 42582 13184
rect 43162 13132 43168 13184
rect 43220 13132 43226 13184
rect 45278 13132 45284 13184
rect 45336 13132 45342 13184
rect 45388 13181 45416 13212
rect 45756 13181 45784 13212
rect 45373 13175 45431 13181
rect 45373 13141 45385 13175
rect 45419 13141 45431 13175
rect 45373 13135 45431 13141
rect 45741 13175 45799 13181
rect 45741 13141 45753 13175
rect 45787 13141 45799 13175
rect 45741 13135 45799 13141
rect 46290 13132 46296 13184
rect 46348 13132 46354 13184
rect 47394 13132 47400 13184
rect 47452 13132 47458 13184
rect 50430 13132 50436 13184
rect 50488 13132 50494 13184
rect 56689 13175 56747 13181
rect 56689 13141 56701 13175
rect 56735 13172 56747 13175
rect 56870 13172 56876 13184
rect 56735 13144 56876 13172
rect 56735 13141 56747 13144
rect 56689 13135 56747 13141
rect 56870 13132 56876 13144
rect 56928 13172 56934 13184
rect 57514 13172 57520 13184
rect 56928 13144 57520 13172
rect 56928 13132 56934 13144
rect 57514 13132 57520 13144
rect 57572 13132 57578 13184
rect 1104 13082 59040 13104
rect 1104 13030 15394 13082
rect 15446 13030 15458 13082
rect 15510 13030 15522 13082
rect 15574 13030 15586 13082
rect 15638 13030 15650 13082
rect 15702 13030 29838 13082
rect 29890 13030 29902 13082
rect 29954 13030 29966 13082
rect 30018 13030 30030 13082
rect 30082 13030 30094 13082
rect 30146 13030 44282 13082
rect 44334 13030 44346 13082
rect 44398 13030 44410 13082
rect 44462 13030 44474 13082
rect 44526 13030 44538 13082
rect 44590 13030 58726 13082
rect 58778 13030 58790 13082
rect 58842 13030 58854 13082
rect 58906 13030 58918 13082
rect 58970 13030 58982 13082
rect 59034 13030 59040 13082
rect 1104 13008 59040 13030
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7742 12968 7748 12980
rect 6963 12940 7748 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 8110 12968 8116 12980
rect 7800 12940 8116 12968
rect 7800 12928 7806 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12768 12940 13093 12968
rect 12768 12928 12774 12940
rect 13081 12937 13093 12940
rect 13127 12968 13139 12971
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 13127 12940 13461 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13449 12937 13461 12940
rect 13495 12968 13507 12971
rect 13630 12968 13636 12980
rect 13495 12940 13636 12968
rect 13495 12937 13507 12940
rect 13449 12931 13507 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13722 12928 13728 12980
rect 13780 12928 13786 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13872 12940 14013 12968
rect 13872 12928 13878 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 18509 12971 18567 12977
rect 18509 12968 18521 12971
rect 14001 12931 14059 12937
rect 14099 12940 18521 12968
rect 2958 12909 2964 12912
rect 2952 12900 2964 12909
rect 2919 12872 2964 12900
rect 2952 12863 2964 12872
rect 2958 12860 2964 12863
rect 3016 12860 3022 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 7650 12900 7656 12912
rect 7064 12872 7656 12900
rect 7064 12860 7070 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 14099 12900 14127 12940
rect 18509 12937 18521 12940
rect 18555 12968 18567 12971
rect 20990 12968 20996 12980
rect 18555 12940 20996 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21450 12928 21456 12980
rect 21508 12968 21514 12980
rect 22094 12968 22100 12980
rect 21508 12940 22100 12968
rect 21508 12928 21514 12940
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 24213 12971 24271 12977
rect 24213 12937 24225 12971
rect 24259 12968 24271 12971
rect 25314 12968 25320 12980
rect 24259 12940 25320 12968
rect 24259 12937 24271 12940
rect 24213 12931 24271 12937
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 26292 12940 26985 12968
rect 26292 12928 26298 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 26973 12931 27031 12937
rect 27985 12971 28043 12977
rect 27985 12937 27997 12971
rect 28031 12968 28043 12971
rect 28994 12968 29000 12980
rect 28031 12940 29000 12968
rect 28031 12937 28043 12940
rect 27985 12931 28043 12937
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 30650 12928 30656 12980
rect 30708 12928 30714 12980
rect 30926 12928 30932 12980
rect 30984 12928 30990 12980
rect 31018 12928 31024 12980
rect 31076 12928 31082 12980
rect 32030 12928 32036 12980
rect 32088 12968 32094 12980
rect 32309 12971 32367 12977
rect 32309 12968 32321 12971
rect 32088 12940 32321 12968
rect 32088 12928 32094 12940
rect 32309 12937 32321 12940
rect 32355 12937 32367 12971
rect 32309 12931 32367 12937
rect 32858 12928 32864 12980
rect 32916 12928 32922 12980
rect 33229 12971 33287 12977
rect 33229 12937 33241 12971
rect 33275 12968 33287 12971
rect 33778 12968 33784 12980
rect 33275 12940 33784 12968
rect 33275 12937 33287 12940
rect 33229 12931 33287 12937
rect 33778 12928 33784 12940
rect 33836 12928 33842 12980
rect 33962 12928 33968 12980
rect 34020 12968 34026 12980
rect 34238 12968 34244 12980
rect 34020 12940 34244 12968
rect 34020 12928 34026 12940
rect 34238 12928 34244 12940
rect 34296 12928 34302 12980
rect 35158 12928 35164 12980
rect 35216 12928 35222 12980
rect 35802 12928 35808 12980
rect 35860 12968 35866 12980
rect 36909 12971 36967 12977
rect 36909 12968 36921 12971
rect 35860 12940 36921 12968
rect 35860 12928 35866 12940
rect 36909 12937 36921 12940
rect 36955 12968 36967 12971
rect 38473 12971 38531 12977
rect 38473 12968 38485 12971
rect 36955 12940 38485 12968
rect 36955 12937 36967 12940
rect 36909 12931 36967 12937
rect 38473 12937 38485 12940
rect 38519 12937 38531 12971
rect 38473 12931 38531 12937
rect 12636 12872 14127 12900
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 12636 12841 12664 12872
rect 14366 12860 14372 12912
rect 14424 12860 14430 12912
rect 15010 12860 15016 12912
rect 15068 12900 15074 12912
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 15068 12872 15117 12900
rect 15068 12860 15074 12872
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15105 12863 15163 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 15565 12903 15623 12909
rect 15565 12900 15577 12903
rect 15252 12872 15577 12900
rect 15252 12860 15258 12872
rect 15565 12869 15577 12872
rect 15611 12869 15623 12903
rect 15565 12863 15623 12869
rect 15746 12860 15752 12912
rect 15804 12860 15810 12912
rect 16776 12872 19104 12900
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 10284 12804 12633 12832
rect 10284 12792 10290 12804
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 13909 12835 13967 12841
rect 13909 12801 13921 12835
rect 13955 12801 13967 12835
rect 14384 12832 14412 12860
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 14384 12804 14565 12832
rect 13909 12795 13967 12801
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 15764 12832 15792 12860
rect 16776 12844 16804 12872
rect 19076 12844 19104 12872
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 30374 12900 30380 12912
rect 20036 12872 30380 12900
rect 20036 12860 20042 12872
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 30561 12903 30619 12909
rect 30561 12869 30573 12903
rect 30607 12900 30619 12903
rect 30944 12900 30972 12928
rect 30607 12872 30972 12900
rect 30607 12869 30619 12872
rect 30561 12863 30619 12869
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15764 12804 16129 12832
rect 14553 12795 14611 12801
rect 16117 12801 16129 12804
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12733 2743 12767
rect 2685 12727 2743 12733
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7374 12764 7380 12776
rect 7239 12736 7380 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 2700 12628 2728 12727
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12696 4123 12699
rect 4172 12696 4200 12727
rect 7374 12724 7380 12736
rect 7432 12764 7438 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7432 12736 7941 12764
rect 7432 12724 7438 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 13924 12764 13952 12795
rect 16758 12792 16764 12844
rect 16816 12792 16822 12844
rect 17028 12835 17086 12841
rect 17028 12801 17040 12835
rect 17074 12832 17086 12835
rect 17586 12832 17592 12844
rect 17074 12804 17592 12832
rect 17074 12801 17086 12804
rect 17028 12795 17086 12801
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19116 12804 20085 12832
rect 19116 12792 19122 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20340 12835 20398 12841
rect 20340 12801 20352 12835
rect 20386 12832 20398 12835
rect 20898 12832 20904 12844
rect 20386 12804 20904 12832
rect 20386 12801 20398 12804
rect 20340 12795 20398 12801
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 22370 12792 22376 12844
rect 22428 12792 22434 12844
rect 22640 12835 22698 12841
rect 22640 12801 22652 12835
rect 22686 12832 22698 12835
rect 23014 12832 23020 12844
rect 22686 12804 23020 12832
rect 22686 12801 22698 12804
rect 22640 12795 22698 12801
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 25676 12835 25734 12841
rect 25676 12801 25688 12835
rect 25722 12832 25734 12835
rect 26418 12832 26424 12844
rect 25722 12804 26424 12832
rect 25722 12801 25734 12804
rect 25676 12795 25734 12801
rect 26418 12792 26424 12804
rect 26476 12792 26482 12844
rect 27893 12835 27951 12841
rect 27893 12801 27905 12835
rect 27939 12801 27951 12835
rect 27893 12795 27951 12801
rect 14826 12764 14832 12776
rect 13924 12736 14832 12764
rect 7929 12727 7987 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15194 12724 15200 12776
rect 15252 12724 15258 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 4111 12668 4200 12696
rect 5353 12699 5411 12705
rect 4111 12665 4123 12668
rect 4065 12659 4123 12665
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 6822 12696 6828 12708
rect 5399 12668 6828 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 6822 12656 6828 12668
rect 6880 12696 6886 12708
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 6880 12668 7665 12696
rect 6880 12656 6886 12668
rect 7653 12665 7665 12668
rect 7699 12696 7711 12699
rect 7699 12668 8064 12696
rect 7699 12665 7711 12668
rect 7653 12659 7711 12665
rect 8036 12640 8064 12668
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14550 12696 14556 12708
rect 13964 12668 14556 12696
rect 13964 12656 13970 12668
rect 14550 12656 14556 12668
rect 14608 12696 14614 12708
rect 15304 12696 15332 12727
rect 23842 12724 23848 12776
rect 23900 12764 23906 12776
rect 24397 12767 24455 12773
rect 24397 12764 24409 12767
rect 23900 12736 24409 12764
rect 23900 12724 23906 12736
rect 24397 12733 24409 12736
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12733 24731 12767
rect 24673 12727 24731 12733
rect 14608 12668 15332 12696
rect 23753 12699 23811 12705
rect 14608 12656 14614 12668
rect 23753 12665 23765 12699
rect 23799 12696 23811 12699
rect 24688 12696 24716 12727
rect 25406 12724 25412 12776
rect 25464 12724 25470 12776
rect 27525 12767 27583 12773
rect 27525 12764 27537 12767
rect 26804 12736 27537 12764
rect 26804 12705 26832 12736
rect 27525 12733 27537 12736
rect 27571 12733 27583 12767
rect 27908 12764 27936 12795
rect 27982 12792 27988 12844
rect 28040 12832 28046 12844
rect 28169 12835 28227 12841
rect 28169 12832 28181 12835
rect 28040 12804 28181 12832
rect 28040 12792 28046 12804
rect 28169 12801 28181 12804
rect 28215 12801 28227 12835
rect 28169 12795 28227 12801
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12801 29423 12835
rect 29365 12795 29423 12801
rect 29457 12835 29515 12841
rect 29457 12801 29469 12835
rect 29503 12832 29515 12835
rect 30576 12832 30604 12863
rect 31036 12841 31064 12928
rect 33321 12903 33379 12909
rect 33321 12869 33333 12903
rect 33367 12900 33379 12903
rect 34974 12900 34980 12912
rect 33367 12872 34980 12900
rect 33367 12869 33379 12872
rect 33321 12863 33379 12869
rect 34974 12860 34980 12872
rect 35032 12860 35038 12912
rect 36078 12900 36084 12912
rect 36004 12872 36084 12900
rect 29503 12804 30604 12832
rect 31021 12835 31079 12841
rect 29503 12801 29515 12804
rect 29457 12795 29515 12801
rect 31021 12801 31033 12835
rect 31067 12801 31079 12835
rect 31021 12795 31079 12801
rect 29178 12764 29184 12776
rect 27908 12736 29184 12764
rect 27525 12727 27583 12733
rect 29178 12724 29184 12736
rect 29236 12724 29242 12776
rect 23799 12668 24716 12696
rect 26789 12699 26847 12705
rect 23799 12665 23811 12668
rect 23753 12659 23811 12665
rect 26789 12665 26801 12699
rect 26835 12665 26847 12699
rect 26789 12659 26847 12665
rect 26878 12656 26884 12708
rect 26936 12696 26942 12708
rect 28902 12696 28908 12708
rect 26936 12668 28908 12696
rect 26936 12656 26942 12668
rect 28902 12656 28908 12668
rect 28960 12656 28966 12708
rect 29380 12696 29408 12795
rect 35342 12792 35348 12844
rect 35400 12832 35406 12844
rect 36004 12841 36032 12872
rect 36078 12860 36084 12872
rect 36136 12860 36142 12912
rect 36630 12860 36636 12912
rect 36688 12860 36694 12912
rect 37550 12860 37556 12912
rect 37608 12860 37614 12912
rect 37734 12860 37740 12912
rect 37792 12860 37798 12912
rect 35713 12835 35771 12841
rect 35713 12832 35725 12835
rect 35400 12804 35725 12832
rect 35400 12792 35406 12804
rect 35713 12801 35725 12804
rect 35759 12801 35771 12835
rect 35713 12795 35771 12801
rect 35989 12835 36047 12841
rect 35989 12801 36001 12835
rect 36035 12801 36047 12835
rect 37752 12832 37780 12860
rect 38105 12835 38163 12841
rect 38105 12832 38117 12835
rect 37752 12804 38117 12832
rect 35989 12795 36047 12801
rect 38105 12801 38117 12804
rect 38151 12801 38163 12835
rect 38488 12832 38516 12931
rect 39850 12928 39856 12980
rect 39908 12968 39914 12980
rect 41417 12971 41475 12977
rect 41417 12968 41429 12971
rect 39908 12940 41429 12968
rect 39908 12928 39914 12940
rect 41417 12937 41429 12940
rect 41463 12937 41475 12971
rect 41417 12931 41475 12937
rect 41598 12928 41604 12980
rect 41656 12968 41662 12980
rect 42153 12971 42211 12977
rect 42153 12968 42165 12971
rect 41656 12940 42165 12968
rect 41656 12928 41662 12940
rect 42153 12937 42165 12940
rect 42199 12968 42211 12971
rect 42613 12971 42671 12977
rect 42613 12968 42625 12971
rect 42199 12940 42625 12968
rect 42199 12937 42211 12940
rect 42153 12931 42211 12937
rect 42613 12937 42625 12940
rect 42659 12937 42671 12971
rect 42613 12931 42671 12937
rect 42978 12928 42984 12980
rect 43036 12968 43042 12980
rect 43257 12971 43315 12977
rect 43257 12968 43269 12971
rect 43036 12940 43269 12968
rect 43036 12928 43042 12940
rect 43257 12937 43269 12940
rect 43303 12937 43315 12971
rect 43257 12931 43315 12937
rect 43349 12971 43407 12977
rect 43349 12937 43361 12971
rect 43395 12968 43407 12971
rect 43438 12968 43444 12980
rect 43395 12940 43444 12968
rect 43395 12937 43407 12940
rect 43349 12931 43407 12937
rect 43438 12928 43444 12940
rect 43496 12968 43502 12980
rect 45278 12968 45284 12980
rect 43496 12940 45284 12968
rect 43496 12928 43502 12940
rect 45278 12928 45284 12940
rect 45336 12928 45342 12980
rect 45370 12928 45376 12980
rect 45428 12928 45434 12980
rect 47121 12971 47179 12977
rect 47121 12937 47133 12971
rect 47167 12968 47179 12971
rect 47210 12968 47216 12980
rect 47167 12940 47216 12968
rect 47167 12937 47179 12940
rect 47121 12931 47179 12937
rect 47210 12928 47216 12940
rect 47268 12928 47274 12980
rect 47394 12928 47400 12980
rect 47452 12928 47458 12980
rect 49970 12928 49976 12980
rect 50028 12968 50034 12980
rect 50065 12971 50123 12977
rect 50065 12968 50077 12971
rect 50028 12940 50077 12968
rect 50028 12928 50034 12940
rect 50065 12937 50077 12940
rect 50111 12937 50123 12971
rect 50065 12931 50123 12937
rect 39200 12903 39258 12909
rect 39200 12869 39212 12903
rect 39246 12900 39258 12903
rect 40034 12900 40040 12912
rect 39246 12872 40040 12900
rect 39246 12869 39258 12872
rect 39200 12863 39258 12869
rect 40034 12860 40040 12872
rect 40092 12860 40098 12912
rect 40770 12860 40776 12912
rect 40828 12860 40834 12912
rect 42518 12860 42524 12912
rect 42576 12900 42582 12912
rect 43714 12900 43720 12912
rect 42576 12872 43720 12900
rect 42576 12860 42582 12872
rect 43714 12860 43720 12872
rect 43772 12900 43778 12912
rect 43901 12903 43959 12909
rect 43901 12900 43913 12903
rect 43772 12872 43913 12900
rect 43772 12860 43778 12872
rect 43901 12869 43913 12872
rect 43947 12869 43959 12903
rect 43901 12863 43959 12869
rect 38933 12835 38991 12841
rect 38933 12832 38945 12835
rect 38488 12804 38945 12832
rect 38105 12795 38163 12801
rect 38933 12801 38945 12804
rect 38979 12801 38991 12835
rect 41785 12835 41843 12841
rect 41785 12832 41797 12835
rect 38933 12795 38991 12801
rect 40972 12804 41797 12832
rect 40972 12776 41000 12804
rect 41785 12801 41797 12804
rect 41831 12832 41843 12835
rect 45186 12832 45192 12844
rect 41831 12804 45192 12832
rect 41831 12801 41843 12804
rect 41785 12795 41843 12801
rect 45186 12792 45192 12804
rect 45244 12792 45250 12844
rect 45388 12832 45416 12928
rect 46008 12903 46066 12909
rect 46008 12869 46020 12903
rect 46054 12900 46066 12903
rect 47412 12900 47440 12928
rect 46054 12872 47440 12900
rect 46054 12869 46066 12872
rect 46008 12863 46066 12869
rect 45741 12835 45799 12841
rect 45741 12832 45753 12835
rect 45388 12804 45753 12832
rect 45741 12801 45753 12804
rect 45787 12801 45799 12835
rect 50080 12832 50108 12931
rect 54938 12928 54944 12980
rect 54996 12968 55002 12980
rect 55033 12971 55091 12977
rect 55033 12968 55045 12971
rect 54996 12940 55045 12968
rect 54996 12928 55002 12940
rect 55033 12937 55045 12940
rect 55079 12968 55091 12971
rect 55122 12968 55128 12980
rect 55079 12940 55128 12968
rect 55079 12937 55091 12940
rect 55033 12931 55091 12937
rect 55122 12928 55128 12940
rect 55180 12928 55186 12980
rect 55493 12971 55551 12977
rect 55493 12937 55505 12971
rect 55539 12968 55551 12971
rect 55582 12968 55588 12980
rect 55539 12940 55588 12968
rect 55539 12937 55551 12940
rect 55493 12931 55551 12937
rect 55582 12928 55588 12940
rect 55640 12928 55646 12980
rect 58066 12860 58072 12912
rect 58124 12900 58130 12912
rect 58253 12903 58311 12909
rect 58253 12900 58265 12903
rect 58124 12872 58265 12900
rect 58124 12860 58130 12872
rect 58253 12869 58265 12872
rect 58299 12869 58311 12903
rect 58253 12863 58311 12869
rect 50522 12841 50528 12844
rect 50249 12835 50307 12841
rect 50249 12832 50261 12835
rect 50080 12804 50261 12832
rect 45741 12795 45799 12801
rect 50249 12801 50261 12804
rect 50295 12801 50307 12835
rect 50249 12795 50307 12801
rect 50516 12795 50528 12841
rect 50522 12792 50528 12795
rect 50580 12792 50586 12844
rect 56962 12792 56968 12844
rect 57020 12792 57026 12844
rect 58434 12792 58440 12844
rect 58492 12792 58498 12844
rect 29638 12724 29644 12776
rect 29696 12724 29702 12776
rect 30837 12767 30895 12773
rect 30837 12733 30849 12767
rect 30883 12764 30895 12767
rect 31294 12764 31300 12776
rect 30883 12736 31300 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 31294 12724 31300 12736
rect 31352 12724 31358 12776
rect 33505 12767 33563 12773
rect 33505 12733 33517 12767
rect 33551 12764 33563 12767
rect 33962 12764 33968 12776
rect 33551 12736 33968 12764
rect 33551 12733 33563 12736
rect 33505 12727 33563 12733
rect 33962 12724 33968 12736
rect 34020 12724 34026 12776
rect 40865 12767 40923 12773
rect 40865 12733 40877 12767
rect 40911 12733 40923 12767
rect 40865 12727 40923 12733
rect 31110 12696 31116 12708
rect 29380 12668 31116 12696
rect 31110 12656 31116 12668
rect 31168 12696 31174 12708
rect 31665 12699 31723 12705
rect 31665 12696 31677 12699
rect 31168 12668 31677 12696
rect 31168 12656 31174 12668
rect 31665 12665 31677 12668
rect 31711 12665 31723 12699
rect 40880 12696 40908 12727
rect 40954 12724 40960 12776
rect 41012 12724 41018 12776
rect 43070 12724 43076 12776
rect 43128 12724 43134 12776
rect 48314 12724 48320 12776
rect 48372 12724 48378 12776
rect 54662 12724 54668 12776
rect 54720 12724 54726 12776
rect 55953 12767 56011 12773
rect 55953 12733 55965 12767
rect 55999 12764 56011 12767
rect 55999 12736 56640 12764
rect 55999 12733 56011 12736
rect 55953 12727 56011 12733
rect 31665 12659 31723 12665
rect 39868 12668 40908 12696
rect 43088 12696 43116 12724
rect 50062 12696 50068 12708
rect 43088 12668 45140 12696
rect 2958 12628 2964 12640
rect 2700 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 4798 12588 4804 12640
rect 4856 12588 4862 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 7006 12628 7012 12640
rect 6595 12600 7012 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 8018 12588 8024 12640
rect 8076 12588 8082 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10318 12628 10324 12640
rect 10091 12600 10324 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 14734 12588 14740 12640
rect 14792 12588 14798 12640
rect 18138 12588 18144 12640
rect 18196 12588 18202 12640
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 21266 12628 21272 12640
rect 21140 12600 21272 12628
rect 21140 12588 21146 12600
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 23842 12588 23848 12640
rect 23900 12588 23906 12640
rect 28442 12588 28448 12640
rect 28500 12628 28506 12640
rect 28813 12631 28871 12637
rect 28813 12628 28825 12631
rect 28500 12600 28825 12628
rect 28500 12588 28506 12600
rect 28813 12597 28825 12600
rect 28859 12597 28871 12631
rect 28813 12591 28871 12597
rect 28994 12588 29000 12640
rect 29052 12588 29058 12640
rect 29730 12588 29736 12640
rect 29788 12628 29794 12640
rect 30009 12631 30067 12637
rect 30009 12628 30021 12631
rect 29788 12600 30021 12628
rect 29788 12588 29794 12600
rect 30009 12597 30021 12600
rect 30055 12597 30067 12631
rect 30009 12591 30067 12597
rect 30193 12631 30251 12637
rect 30193 12597 30205 12631
rect 30239 12628 30251 12631
rect 30650 12628 30656 12640
rect 30239 12600 30656 12628
rect 30239 12597 30251 12600
rect 30193 12591 30251 12597
rect 30650 12588 30656 12600
rect 30708 12588 30714 12640
rect 32674 12588 32680 12640
rect 32732 12588 32738 12640
rect 38470 12588 38476 12640
rect 38528 12628 38534 12640
rect 39868 12628 39896 12668
rect 38528 12600 39896 12628
rect 38528 12588 38534 12600
rect 40310 12588 40316 12640
rect 40368 12588 40374 12640
rect 40402 12588 40408 12640
rect 40460 12588 40466 12640
rect 42426 12588 42432 12640
rect 42484 12628 42490 12640
rect 42610 12628 42616 12640
rect 42484 12600 42616 12628
rect 42484 12588 42490 12600
rect 42610 12588 42616 12600
rect 42668 12588 42674 12640
rect 43717 12631 43775 12637
rect 43717 12597 43729 12631
rect 43763 12628 43775 12631
rect 44082 12628 44088 12640
rect 43763 12600 44088 12628
rect 43763 12597 43775 12600
rect 43717 12591 43775 12597
rect 44082 12588 44088 12600
rect 44140 12588 44146 12640
rect 45112 12628 45140 12668
rect 47688 12668 50068 12696
rect 47688 12628 47716 12668
rect 50062 12656 50068 12668
rect 50120 12656 50126 12708
rect 56612 12705 56640 12736
rect 57054 12724 57060 12776
rect 57112 12724 57118 12776
rect 57146 12724 57152 12776
rect 57204 12764 57210 12776
rect 57609 12767 57667 12773
rect 57609 12764 57621 12767
rect 57204 12736 57621 12764
rect 57204 12724 57210 12736
rect 57609 12733 57621 12736
rect 57655 12733 57667 12767
rect 57609 12727 57667 12733
rect 56597 12699 56655 12705
rect 56597 12665 56609 12699
rect 56643 12665 56655 12699
rect 56597 12659 56655 12665
rect 45112 12600 47716 12628
rect 47762 12588 47768 12640
rect 47820 12588 47826 12640
rect 51629 12631 51687 12637
rect 51629 12597 51641 12631
rect 51675 12628 51687 12631
rect 52270 12628 52276 12640
rect 51675 12600 52276 12628
rect 51675 12597 51687 12600
rect 51629 12591 51687 12597
rect 52270 12588 52276 12600
rect 52328 12588 52334 12640
rect 54110 12588 54116 12640
rect 54168 12588 54174 12640
rect 56505 12631 56563 12637
rect 56505 12597 56517 12631
rect 56551 12628 56563 12631
rect 56686 12628 56692 12640
rect 56551 12600 56692 12628
rect 56551 12597 56563 12600
rect 56505 12591 56563 12597
rect 56686 12588 56692 12600
rect 56744 12588 56750 12640
rect 1104 12538 58880 12560
rect 1104 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 22616 12538
rect 22668 12486 22680 12538
rect 22732 12486 22744 12538
rect 22796 12486 22808 12538
rect 22860 12486 22872 12538
rect 22924 12486 37060 12538
rect 37112 12486 37124 12538
rect 37176 12486 37188 12538
rect 37240 12486 37252 12538
rect 37304 12486 37316 12538
rect 37368 12486 51504 12538
rect 51556 12486 51568 12538
rect 51620 12486 51632 12538
rect 51684 12486 51696 12538
rect 51748 12486 51760 12538
rect 51812 12486 58880 12538
rect 1104 12464 58880 12486
rect 6454 12384 6460 12436
rect 6512 12384 6518 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 7616 12396 10609 12424
rect 7616 12384 7622 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 13906 12424 13912 12436
rect 10836 12396 13912 12424
rect 10836 12384 10842 12396
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 15841 12427 15899 12433
rect 14200 12396 15792 12424
rect 5169 12359 5227 12365
rect 5169 12325 5181 12359
rect 5215 12356 5227 12359
rect 5215 12328 5856 12356
rect 5215 12325 5227 12328
rect 5169 12319 5227 12325
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 5828 12297 5856 12328
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 10796 12356 10824 12384
rect 7800 12328 10824 12356
rect 7800 12316 7806 12328
rect 13538 12316 13544 12368
rect 13596 12356 13602 12368
rect 14200 12356 14228 12396
rect 13596 12328 14228 12356
rect 15764 12356 15792 12396
rect 15841 12393 15853 12427
rect 15887 12424 15899 12427
rect 15930 12424 15936 12436
rect 15887 12396 15936 12424
rect 15887 12393 15899 12396
rect 15841 12387 15899 12393
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 16758 12424 16764 12436
rect 16715 12396 16764 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17586 12384 17592 12436
rect 17644 12384 17650 12436
rect 18874 12424 18880 12436
rect 18156 12396 18880 12424
rect 18156 12356 18184 12396
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 19978 12424 19984 12436
rect 19843 12396 19984 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21082 12424 21088 12436
rect 21039 12396 21088 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21542 12384 21548 12436
rect 21600 12384 21606 12436
rect 23014 12384 23020 12436
rect 23072 12424 23078 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 23072 12396 23305 12424
rect 23072 12384 23078 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 23293 12387 23351 12393
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 24857 12427 24915 12433
rect 24857 12424 24869 12427
rect 23440 12396 24869 12424
rect 23440 12384 23446 12396
rect 24857 12393 24869 12396
rect 24903 12424 24915 12427
rect 24903 12396 25912 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 15764 12328 18184 12356
rect 18325 12359 18383 12365
rect 13596 12316 13602 12328
rect 18325 12325 18337 12359
rect 18371 12325 18383 12359
rect 21361 12359 21419 12365
rect 21361 12356 21373 12359
rect 18325 12319 18383 12325
rect 20548 12328 21373 12356
rect 5813 12291 5871 12297
rect 3016 12260 3832 12288
rect 3016 12248 3022 12260
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3804 12229 3832 12260
rect 5813 12257 5825 12291
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7116 12260 8125 12288
rect 3513 12223 3571 12229
rect 3513 12220 3525 12223
rect 3344 12192 3525 12220
rect 2716 12155 2774 12161
rect 2716 12121 2728 12155
rect 2762 12152 2774 12155
rect 2958 12152 2964 12164
rect 2762 12124 2964 12152
rect 2762 12121 2774 12124
rect 2716 12115 2774 12121
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 3344 12096 3372 12192
rect 3513 12189 3525 12192
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 3878 12220 3884 12232
rect 3835 12192 3884 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7116 12220 7144 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 9548 12260 10333 12288
rect 9548 12248 9554 12260
rect 10321 12257 10333 12260
rect 10367 12288 10379 12291
rect 10502 12288 10508 12300
rect 10367 12260 10508 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10502 12248 10508 12260
rect 10560 12288 10566 12300
rect 12158 12288 12164 12300
rect 10560 12260 12164 12288
rect 10560 12248 10566 12260
rect 12158 12248 12164 12260
rect 12216 12288 12222 12300
rect 14090 12288 14096 12300
rect 12216 12260 14096 12288
rect 12216 12248 12222 12260
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18340 12288 18368 12319
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 18279 12260 18368 12288
rect 18432 12260 18889 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 6696 12192 7144 12220
rect 7469 12223 7527 12229
rect 6696 12180 6702 12192
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 8018 12220 8024 12232
rect 7515 12192 8024 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 10778 12180 10784 12232
rect 10836 12180 10842 12232
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12308 12192 12725 12220
rect 12308 12180 12314 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13964 12192 14197 12220
rect 13964 12180 13970 12192
rect 14185 12189 14197 12192
rect 14231 12220 14243 12223
rect 14274 12220 14280 12232
rect 14231 12192 14280 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14452 12223 14510 12229
rect 14452 12189 14464 12223
rect 14498 12220 14510 12223
rect 14734 12220 14740 12232
rect 14498 12192 14740 12220
rect 14498 12189 14510 12192
rect 14452 12183 14510 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17310 12220 17316 12232
rect 17083 12192 17316 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 18432 12220 18460 12260
rect 18877 12257 18889 12260
rect 18923 12288 18935 12291
rect 20162 12288 20168 12300
rect 18923 12260 20168 12288
rect 18923 12257 18935 12260
rect 18877 12251 18935 12257
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 20548 12297 20576 12328
rect 21361 12325 21373 12328
rect 21407 12325 21419 12359
rect 21361 12319 21419 12325
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 18340 12192 18460 12220
rect 18693 12223 18751 12229
rect 4056 12155 4114 12161
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4246 12152 4252 12164
rect 4102 12124 4252 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 10244 12152 10272 12180
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10244 12124 10885 12152
rect 10873 12121 10885 12124
rect 10919 12152 10931 12155
rect 11422 12152 11428 12164
rect 10919 12124 11428 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 1578 12044 1584 12096
rect 1636 12044 1642 12096
rect 3050 12044 3056 12096
rect 3108 12044 3114 12096
rect 3326 12044 3332 12096
rect 3384 12044 3390 12096
rect 3418 12044 3424 12096
rect 3476 12044 3482 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5261 12087 5319 12093
rect 5261 12084 5273 12087
rect 5132 12056 5273 12084
rect 5132 12044 5138 12056
rect 5261 12053 5273 12056
rect 5307 12053 5319 12087
rect 5261 12047 5319 12053
rect 7558 12044 7564 12096
rect 7616 12044 7622 12096
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 8662 12084 8668 12096
rect 8619 12056 8668 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9766 12044 9772 12096
rect 9824 12044 9830 12096
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11020 12056 12173 12084
rect 11020 12044 11026 12056
rect 12161 12053 12173 12056
rect 12207 12084 12219 12087
rect 12710 12084 12716 12096
rect 12207 12056 12716 12084
rect 12207 12053 12219 12056
rect 12161 12047 12219 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13556 12084 13584 12115
rect 15746 12112 15752 12164
rect 15804 12112 15810 12164
rect 18340 12096 18368 12192
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 20070 12220 20076 12232
rect 18739 12192 20076 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 20824 12220 20852 12248
rect 20395 12192 20852 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 18840 12124 20300 12152
rect 18840 12112 18846 12124
rect 13906 12084 13912 12096
rect 13556 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 16114 12084 16120 12096
rect 15611 12056 16120 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 16448 12056 16865 12084
rect 16448 12044 16454 12056
rect 16853 12053 16865 12056
rect 16899 12053 16911 12087
rect 16853 12047 16911 12053
rect 18322 12044 18328 12096
rect 18380 12044 18386 12096
rect 19886 12044 19892 12096
rect 19944 12044 19950 12096
rect 20272 12093 20300 12124
rect 20898 12112 20904 12164
rect 20956 12112 20962 12164
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12084 20315 12087
rect 20714 12084 20720 12096
rect 20303 12056 20720 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 20714 12044 20720 12056
rect 20772 12084 20778 12096
rect 20990 12084 20996 12096
rect 20772 12056 20996 12084
rect 20772 12044 20778 12056
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 21376 12084 21404 12319
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21508 12328 25820 12356
rect 21508 12316 21514 12328
rect 22094 12248 22100 12300
rect 22152 12248 22158 12300
rect 23842 12248 23848 12300
rect 23900 12248 23906 12300
rect 25498 12288 25504 12300
rect 24504 12260 25504 12288
rect 24504 12096 24532 12260
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 25130 12180 25136 12232
rect 25188 12220 25194 12232
rect 25317 12223 25375 12229
rect 25317 12220 25329 12223
rect 25188 12192 25329 12220
rect 25188 12180 25194 12192
rect 25317 12189 25329 12192
rect 25363 12189 25375 12223
rect 25792 12220 25820 12328
rect 25884 12297 25912 12396
rect 26418 12384 26424 12436
rect 26476 12424 26482 12436
rect 26605 12427 26663 12433
rect 26605 12424 26617 12427
rect 26476 12396 26617 12424
rect 26476 12384 26482 12396
rect 26605 12393 26617 12396
rect 26651 12393 26663 12427
rect 26605 12387 26663 12393
rect 28626 12384 28632 12436
rect 28684 12384 28690 12436
rect 29178 12384 29184 12436
rect 29236 12424 29242 12436
rect 29454 12424 29460 12436
rect 29236 12396 29460 12424
rect 29236 12384 29242 12396
rect 29454 12384 29460 12396
rect 29512 12384 29518 12436
rect 29730 12384 29736 12436
rect 29788 12384 29794 12436
rect 30101 12427 30159 12433
rect 30101 12393 30113 12427
rect 30147 12424 30159 12427
rect 30282 12424 30288 12436
rect 30147 12396 30288 12424
rect 30147 12393 30159 12396
rect 30101 12387 30159 12393
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 40497 12427 40555 12433
rect 40497 12393 40509 12427
rect 40543 12424 40555 12427
rect 40770 12424 40776 12436
rect 40543 12396 40776 12424
rect 40543 12393 40555 12396
rect 40497 12387 40555 12393
rect 40770 12384 40776 12396
rect 40828 12384 40834 12436
rect 42334 12384 42340 12436
rect 42392 12384 42398 12436
rect 42978 12384 42984 12436
rect 43036 12424 43042 12436
rect 43073 12427 43131 12433
rect 43073 12424 43085 12427
rect 43036 12396 43085 12424
rect 43036 12384 43042 12396
rect 43073 12393 43085 12396
rect 43119 12393 43131 12427
rect 43073 12387 43131 12393
rect 44726 12384 44732 12436
rect 44784 12384 44790 12436
rect 45186 12384 45192 12436
rect 45244 12424 45250 12436
rect 45554 12424 45560 12436
rect 45244 12396 45560 12424
rect 45244 12384 45250 12396
rect 45554 12384 45560 12396
rect 45612 12384 45618 12436
rect 46017 12427 46075 12433
rect 46017 12393 46029 12427
rect 46063 12424 46075 12427
rect 46106 12424 46112 12436
rect 46063 12396 46112 12424
rect 46063 12393 46075 12396
rect 46017 12387 46075 12393
rect 46106 12384 46112 12396
rect 46164 12424 46170 12436
rect 46164 12396 49464 12424
rect 46164 12384 46170 12396
rect 45094 12356 45100 12368
rect 25976 12328 45100 12356
rect 25869 12291 25927 12297
rect 25869 12257 25881 12291
rect 25915 12257 25927 12291
rect 25869 12251 25927 12257
rect 25976 12220 26004 12328
rect 45094 12316 45100 12328
rect 45152 12316 45158 12368
rect 46474 12316 46480 12368
rect 46532 12356 46538 12368
rect 47029 12359 47087 12365
rect 47029 12356 47041 12359
rect 46532 12328 47041 12356
rect 46532 12316 46538 12328
rect 47029 12325 47041 12328
rect 47075 12325 47087 12359
rect 47029 12319 47087 12325
rect 48685 12359 48743 12365
rect 48685 12325 48697 12359
rect 48731 12356 48743 12359
rect 49436 12356 49464 12396
rect 50522 12384 50528 12436
rect 50580 12424 50586 12436
rect 50709 12427 50767 12433
rect 50709 12424 50721 12427
rect 50580 12396 50721 12424
rect 50580 12384 50586 12396
rect 50709 12393 50721 12396
rect 50755 12393 50767 12427
rect 50709 12387 50767 12393
rect 51994 12384 52000 12436
rect 52052 12384 52058 12436
rect 53834 12384 53840 12436
rect 53892 12424 53898 12436
rect 53929 12427 53987 12433
rect 53929 12424 53941 12427
rect 53892 12396 53941 12424
rect 53892 12384 53898 12396
rect 53929 12393 53941 12396
rect 53975 12393 53987 12427
rect 53929 12387 53987 12393
rect 54113 12427 54171 12433
rect 54113 12393 54125 12427
rect 54159 12424 54171 12427
rect 54662 12424 54668 12436
rect 54159 12396 54668 12424
rect 54159 12393 54171 12396
rect 54113 12387 54171 12393
rect 50617 12359 50675 12365
rect 50617 12356 50629 12359
rect 48731 12328 49372 12356
rect 49436 12328 50629 12356
rect 48731 12325 48743 12328
rect 48685 12319 48743 12325
rect 26053 12291 26111 12297
rect 26053 12257 26065 12291
rect 26099 12288 26111 12291
rect 26234 12288 26240 12300
rect 26099 12260 26240 12288
rect 26099 12257 26111 12260
rect 26053 12251 26111 12257
rect 26234 12248 26240 12260
rect 26292 12248 26298 12300
rect 29178 12248 29184 12300
rect 29236 12248 29242 12300
rect 30650 12248 30656 12300
rect 30708 12248 30714 12300
rect 39298 12248 39304 12300
rect 39356 12288 39362 12300
rect 39853 12291 39911 12297
rect 39853 12288 39865 12291
rect 39356 12260 39865 12288
rect 39356 12248 39362 12260
rect 39853 12257 39865 12260
rect 39899 12257 39911 12291
rect 39853 12251 39911 12257
rect 40402 12248 40408 12300
rect 40460 12288 40466 12300
rect 41141 12291 41199 12297
rect 41141 12288 41153 12291
rect 40460 12260 41153 12288
rect 40460 12248 40466 12260
rect 41141 12257 41153 12260
rect 41187 12257 41199 12291
rect 41141 12251 41199 12257
rect 42886 12248 42892 12300
rect 42944 12248 42950 12300
rect 43162 12248 43168 12300
rect 43220 12288 43226 12300
rect 43625 12291 43683 12297
rect 43625 12288 43637 12291
rect 43220 12260 43637 12288
rect 43220 12248 43226 12260
rect 43625 12257 43637 12260
rect 43671 12257 43683 12291
rect 43625 12251 43683 12257
rect 44082 12248 44088 12300
rect 44140 12248 44146 12300
rect 47302 12288 47308 12300
rect 46860 12260 47308 12288
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 25792 12192 26004 12220
rect 26528 12192 27169 12220
rect 25317 12183 25375 12189
rect 25866 12152 25872 12164
rect 24872 12124 25872 12152
rect 24872 12096 24900 12124
rect 25866 12112 25872 12124
rect 25924 12152 25930 12164
rect 25924 12124 26188 12152
rect 25924 12112 25930 12124
rect 23014 12084 23020 12096
rect 21376 12056 23020 12084
rect 23014 12044 23020 12056
rect 23072 12084 23078 12096
rect 23382 12084 23388 12096
rect 23072 12056 23388 12084
rect 23072 12044 23078 12056
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 24486 12044 24492 12096
rect 24544 12044 24550 12096
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 24946 12044 24952 12096
rect 25004 12044 25010 12096
rect 25222 12044 25228 12096
rect 25280 12084 25286 12096
rect 26160 12093 26188 12124
rect 26528 12093 26556 12192
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 27157 12183 27215 12189
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 28258 12220 28264 12232
rect 27672 12192 28264 12220
rect 27672 12180 27678 12192
rect 28258 12180 28264 12192
rect 28316 12220 28322 12232
rect 37461 12223 37519 12229
rect 37461 12220 37473 12223
rect 28316 12192 37473 12220
rect 28316 12180 28322 12192
rect 37461 12189 37473 12192
rect 37507 12220 37519 12223
rect 37642 12220 37648 12232
rect 37507 12192 37648 12220
rect 37507 12189 37519 12192
rect 37461 12183 37519 12189
rect 37642 12180 37648 12192
rect 37700 12180 37706 12232
rect 39390 12180 39396 12232
rect 39448 12220 39454 12232
rect 40589 12223 40647 12229
rect 40589 12220 40601 12223
rect 39448 12192 40601 12220
rect 39448 12180 39454 12192
rect 40589 12189 40601 12192
rect 40635 12189 40647 12223
rect 40589 12183 40647 12189
rect 44634 12180 44640 12232
rect 44692 12220 44698 12232
rect 45189 12223 45247 12229
rect 45189 12220 45201 12223
rect 44692 12192 45201 12220
rect 44692 12180 44698 12192
rect 45189 12189 45201 12192
rect 45235 12220 45247 12223
rect 46293 12223 46351 12229
rect 46293 12220 46305 12223
rect 45235 12192 46305 12220
rect 45235 12189 45247 12192
rect 45189 12183 45247 12189
rect 46293 12189 46305 12192
rect 46339 12220 46351 12223
rect 46750 12220 46756 12232
rect 46339 12192 46756 12220
rect 46339 12189 46351 12192
rect 46293 12183 46351 12189
rect 46750 12180 46756 12192
rect 46808 12220 46814 12232
rect 46860 12229 46888 12260
rect 47302 12248 47308 12260
rect 47360 12248 47366 12300
rect 49344 12297 49372 12328
rect 50617 12325 50629 12328
rect 50663 12356 50675 12359
rect 50663 12328 51074 12356
rect 50663 12325 50675 12328
rect 50617 12319 50675 12325
rect 49329 12291 49387 12297
rect 49329 12257 49341 12291
rect 49375 12257 49387 12291
rect 51046 12288 51074 12328
rect 51261 12291 51319 12297
rect 51261 12288 51273 12291
rect 51046 12260 51273 12288
rect 49329 12251 49387 12257
rect 51261 12257 51273 12260
rect 51307 12257 51319 12291
rect 53944 12288 53972 12387
rect 54662 12384 54668 12396
rect 54720 12384 54726 12436
rect 55306 12384 55312 12436
rect 55364 12424 55370 12436
rect 56594 12424 56600 12436
rect 55364 12396 56600 12424
rect 55364 12384 55370 12396
rect 56594 12384 56600 12396
rect 56652 12384 56658 12436
rect 57793 12359 57851 12365
rect 57793 12325 57805 12359
rect 57839 12356 57851 12359
rect 57839 12328 58480 12356
rect 57839 12325 57851 12328
rect 57793 12319 57851 12325
rect 58452 12297 58480 12328
rect 54665 12291 54723 12297
rect 54665 12288 54677 12291
rect 53944 12260 54677 12288
rect 51261 12251 51319 12257
rect 54665 12257 54677 12260
rect 54711 12257 54723 12291
rect 54665 12251 54723 12257
rect 58437 12291 58495 12297
rect 58437 12257 58449 12291
rect 58483 12257 58495 12291
rect 58437 12251 58495 12257
rect 46845 12223 46903 12229
rect 46845 12220 46857 12223
rect 46808 12192 46857 12220
rect 46808 12180 46814 12192
rect 46845 12189 46857 12192
rect 46891 12189 46903 12223
rect 46845 12183 46903 12189
rect 47210 12180 47216 12232
rect 47268 12180 47274 12232
rect 51074 12180 51080 12232
rect 51132 12180 51138 12232
rect 52362 12180 52368 12232
rect 52420 12220 52426 12232
rect 52641 12223 52699 12229
rect 52641 12220 52653 12223
rect 52420 12192 52653 12220
rect 52420 12180 52426 12192
rect 52641 12189 52653 12192
rect 52687 12189 52699 12223
rect 52641 12183 52699 12189
rect 55306 12180 55312 12232
rect 55364 12180 55370 12232
rect 56226 12180 56232 12232
rect 56284 12220 56290 12232
rect 56686 12229 56692 12232
rect 56413 12223 56471 12229
rect 56413 12220 56425 12223
rect 56284 12192 56425 12220
rect 56284 12180 56290 12192
rect 56413 12189 56425 12192
rect 56459 12189 56471 12223
rect 56413 12183 56471 12189
rect 56680 12183 56692 12229
rect 56686 12180 56692 12183
rect 56744 12180 56750 12232
rect 42610 12112 42616 12164
rect 42668 12152 42674 12164
rect 42668 12124 43208 12152
rect 42668 12112 42674 12124
rect 25409 12087 25467 12093
rect 25409 12084 25421 12087
rect 25280 12056 25421 12084
rect 25280 12044 25286 12056
rect 25409 12053 25421 12056
rect 25455 12053 25467 12087
rect 25409 12047 25467 12053
rect 26145 12087 26203 12093
rect 26145 12053 26157 12087
rect 26191 12053 26203 12087
rect 26145 12047 26203 12053
rect 26513 12087 26571 12093
rect 26513 12053 26525 12087
rect 26559 12053 26571 12087
rect 26513 12047 26571 12053
rect 27614 12044 27620 12096
rect 27672 12084 27678 12096
rect 27798 12084 27804 12096
rect 27672 12056 27804 12084
rect 27672 12044 27678 12056
rect 27798 12044 27804 12056
rect 27856 12044 27862 12096
rect 31110 12044 31116 12096
rect 31168 12044 31174 12096
rect 35989 12087 36047 12093
rect 35989 12053 36001 12087
rect 36035 12084 36047 12087
rect 36078 12084 36084 12096
rect 36035 12056 36084 12084
rect 36035 12053 36047 12056
rect 35989 12047 36047 12053
rect 36078 12044 36084 12056
rect 36136 12044 36142 12096
rect 36906 12044 36912 12096
rect 36964 12084 36970 12096
rect 37093 12087 37151 12093
rect 37093 12084 37105 12087
rect 36964 12056 37105 12084
rect 36964 12044 36970 12056
rect 37093 12053 37105 12056
rect 37139 12084 37151 12087
rect 38286 12084 38292 12096
rect 37139 12056 38292 12084
rect 37139 12053 37151 12056
rect 37093 12047 37151 12053
rect 38286 12044 38292 12056
rect 38344 12044 38350 12096
rect 41782 12044 41788 12096
rect 41840 12084 41846 12096
rect 42153 12087 42211 12093
rect 42153 12084 42165 12087
rect 41840 12056 42165 12084
rect 41840 12044 41846 12056
rect 42153 12053 42165 12056
rect 42199 12084 42211 12087
rect 43070 12084 43076 12096
rect 42199 12056 43076 12084
rect 42199 12053 42211 12056
rect 42153 12047 42211 12053
rect 43070 12044 43076 12056
rect 43128 12044 43134 12096
rect 43180 12084 43208 12124
rect 45554 12112 45560 12164
rect 45612 12152 45618 12164
rect 47572 12155 47630 12161
rect 45612 12124 47256 12152
rect 45612 12112 45618 12124
rect 46474 12084 46480 12096
rect 43180 12056 46480 12084
rect 46474 12044 46480 12056
rect 46532 12044 46538 12096
rect 47228 12084 47256 12124
rect 47572 12121 47584 12155
rect 47618 12152 47630 12155
rect 49050 12152 49056 12164
rect 47618 12124 49056 12152
rect 47618 12121 47630 12124
rect 47572 12115 47630 12121
rect 49050 12112 49056 12124
rect 49108 12112 49114 12164
rect 52086 12112 52092 12164
rect 52144 12112 52150 12164
rect 54481 12155 54539 12161
rect 54481 12121 54493 12155
rect 54527 12152 54539 12155
rect 55953 12155 56011 12161
rect 55953 12152 55965 12155
rect 54527 12124 55965 12152
rect 54527 12121 54539 12124
rect 54481 12115 54539 12121
rect 55953 12121 55965 12124
rect 55999 12152 56011 12155
rect 56134 12152 56140 12164
rect 55999 12124 56140 12152
rect 55999 12121 56011 12124
rect 55953 12115 56011 12121
rect 56134 12112 56140 12124
rect 56192 12112 56198 12164
rect 48590 12084 48596 12096
rect 47228 12056 48596 12084
rect 48590 12044 48596 12056
rect 48648 12044 48654 12096
rect 48774 12044 48780 12096
rect 48832 12044 48838 12096
rect 51169 12087 51227 12093
rect 51169 12053 51181 12087
rect 51215 12084 51227 12087
rect 51350 12084 51356 12096
rect 51215 12056 51356 12084
rect 51215 12053 51227 12056
rect 51169 12047 51227 12053
rect 51350 12044 51356 12056
rect 51408 12044 51414 12096
rect 52914 12044 52920 12096
rect 52972 12084 52978 12096
rect 53285 12087 53343 12093
rect 53285 12084 53297 12087
rect 52972 12056 53297 12084
rect 52972 12044 52978 12056
rect 53285 12053 53297 12056
rect 53331 12053 53343 12087
rect 53285 12047 53343 12053
rect 54573 12087 54631 12093
rect 54573 12053 54585 12087
rect 54619 12084 54631 12087
rect 54662 12084 54668 12096
rect 54619 12056 54668 12084
rect 54619 12053 54631 12056
rect 54573 12047 54631 12053
rect 54662 12044 54668 12056
rect 54720 12044 54726 12096
rect 57054 12044 57060 12096
rect 57112 12084 57118 12096
rect 57885 12087 57943 12093
rect 57885 12084 57897 12087
rect 57112 12056 57897 12084
rect 57112 12044 57118 12056
rect 57885 12053 57897 12056
rect 57931 12053 57943 12087
rect 57885 12047 57943 12053
rect 1104 11994 59040 12016
rect 1104 11942 15394 11994
rect 15446 11942 15458 11994
rect 15510 11942 15522 11994
rect 15574 11942 15586 11994
rect 15638 11942 15650 11994
rect 15702 11942 29838 11994
rect 29890 11942 29902 11994
rect 29954 11942 29966 11994
rect 30018 11942 30030 11994
rect 30082 11942 30094 11994
rect 30146 11942 44282 11994
rect 44334 11942 44346 11994
rect 44398 11942 44410 11994
rect 44462 11942 44474 11994
rect 44526 11942 44538 11994
rect 44590 11942 58726 11994
rect 58778 11942 58790 11994
rect 58842 11942 58854 11994
rect 58906 11942 58918 11994
rect 58970 11942 58982 11994
rect 59034 11942 59040 11994
rect 1104 11920 59040 11942
rect 1578 11840 1584 11892
rect 1636 11840 1642 11892
rect 2958 11840 2964 11892
rect 3016 11840 3022 11892
rect 3050 11840 3056 11892
rect 3108 11840 3114 11892
rect 3878 11840 3884 11892
rect 3936 11840 3942 11892
rect 4246 11840 4252 11892
rect 4304 11840 4310 11892
rect 11238 11880 11244 11892
rect 9048 11852 11244 11880
rect 1596 11744 1624 11840
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 1596 11716 2237 11744
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 3068 11744 3096 11840
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 9048 11812 9076 11852
rect 11238 11840 11244 11852
rect 11296 11880 11302 11892
rect 16482 11880 16488 11892
rect 11296 11852 16488 11880
rect 11296 11840 11302 11852
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 19797 11883 19855 11889
rect 19797 11880 19809 11883
rect 19760 11852 19809 11880
rect 19760 11840 19766 11852
rect 19797 11849 19809 11852
rect 19843 11849 19855 11883
rect 19797 11843 19855 11849
rect 23750 11840 23756 11892
rect 23808 11840 23814 11892
rect 24946 11840 24952 11892
rect 25004 11840 25010 11892
rect 28905 11883 28963 11889
rect 28905 11849 28917 11883
rect 28951 11880 28963 11883
rect 29730 11880 29736 11892
rect 28951 11852 29736 11880
rect 28951 11849 28963 11852
rect 28905 11843 28963 11849
rect 29730 11840 29736 11852
rect 29788 11840 29794 11892
rect 34882 11840 34888 11892
rect 34940 11880 34946 11892
rect 34977 11883 35035 11889
rect 34977 11880 34989 11883
rect 34940 11852 34989 11880
rect 34940 11840 34946 11852
rect 34977 11849 34989 11852
rect 35023 11849 35035 11883
rect 34977 11843 35035 11849
rect 38197 11883 38255 11889
rect 38197 11849 38209 11883
rect 38243 11880 38255 11883
rect 38562 11880 38568 11892
rect 38243 11852 38568 11880
rect 38243 11849 38255 11852
rect 38197 11843 38255 11849
rect 38562 11840 38568 11852
rect 38620 11840 38626 11892
rect 41417 11883 41475 11889
rect 41417 11849 41429 11883
rect 41463 11880 41475 11883
rect 41598 11880 41604 11892
rect 41463 11852 41604 11880
rect 41463 11849 41475 11852
rect 41417 11843 41475 11849
rect 41598 11840 41604 11852
rect 41656 11880 41662 11892
rect 43349 11883 43407 11889
rect 43349 11880 43361 11883
rect 41656 11852 43361 11880
rect 41656 11840 41662 11852
rect 43349 11849 43361 11852
rect 43395 11880 43407 11883
rect 44085 11883 44143 11889
rect 44085 11880 44097 11883
rect 43395 11852 44097 11880
rect 43395 11849 43407 11852
rect 43349 11843 43407 11849
rect 44085 11849 44097 11852
rect 44131 11880 44143 11883
rect 44450 11880 44456 11892
rect 44131 11852 44456 11880
rect 44131 11849 44143 11852
rect 44085 11843 44143 11849
rect 44450 11840 44456 11852
rect 44508 11840 44514 11892
rect 46750 11840 46756 11892
rect 46808 11840 46814 11892
rect 47581 11883 47639 11889
rect 47581 11849 47593 11883
rect 47627 11880 47639 11883
rect 48314 11880 48320 11892
rect 47627 11852 48320 11880
rect 47627 11849 47639 11852
rect 47581 11843 47639 11849
rect 48314 11840 48320 11852
rect 48372 11840 48378 11892
rect 49050 11840 49056 11892
rect 49108 11840 49114 11892
rect 55125 11883 55183 11889
rect 55125 11849 55137 11883
rect 55171 11880 55183 11883
rect 55306 11880 55312 11892
rect 55171 11852 55312 11880
rect 55171 11849 55183 11852
rect 55125 11843 55183 11849
rect 55306 11840 55312 11852
rect 55364 11840 55370 11892
rect 56226 11880 56232 11892
rect 55416 11852 56232 11880
rect 23658 11812 23664 11824
rect 7340 11784 9076 11812
rect 7340 11772 7346 11784
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3068 11716 3525 11744
rect 2225 11707 2283 11713
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 4706 11744 4712 11756
rect 3513 11707 3571 11713
rect 4356 11716 4712 11744
rect 4356 11676 4384 11716
rect 4706 11704 4712 11716
rect 4764 11744 4770 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4764 11716 4997 11744
rect 4764 11704 4770 11716
rect 4985 11713 4997 11716
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 7466 11704 7472 11756
rect 7524 11753 7530 11756
rect 7524 11707 7536 11753
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 7791 11716 8064 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 7524 11704 7530 11707
rect 8036 11688 8064 11716
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 3160 11648 4384 11676
rect 3160 11620 3188 11648
rect 4798 11636 4804 11688
rect 4856 11636 4862 11688
rect 5074 11636 5080 11688
rect 5132 11636 5138 11688
rect 7926 11636 7932 11688
rect 7984 11636 7990 11688
rect 8018 11636 8024 11688
rect 8076 11636 8082 11688
rect 3142 11568 3148 11620
rect 3200 11568 3206 11620
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 5092 11608 5120 11636
rect 4120 11580 5120 11608
rect 8680 11608 8708 11704
rect 9048 11685 9076 11784
rect 9140 11784 23664 11812
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9140 11608 9168 11784
rect 23658 11772 23664 11784
rect 23716 11772 23722 11824
rect 11330 11704 11336 11756
rect 11388 11704 11394 11756
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11773 11747 11831 11753
rect 11773 11744 11785 11747
rect 11664 11716 11785 11744
rect 11664 11704 11670 11716
rect 11773 11713 11785 11716
rect 11819 11713 11831 11747
rect 11773 11707 11831 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12342 11744 12348 11756
rect 12124 11716 12348 11744
rect 12124 11704 12130 11716
rect 12342 11704 12348 11716
rect 12400 11744 12406 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12400 11716 13093 11744
rect 12400 11704 12406 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10962 11676 10968 11688
rect 10376 11648 10968 11676
rect 10376 11636 10382 11648
rect 10962 11636 10968 11648
rect 11020 11676 11026 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11020 11648 11529 11676
rect 11020 11636 11026 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 13648 11676 13676 11707
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 13780 11716 15117 11744
rect 13780 11704 13786 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11744 15439 11747
rect 16298 11744 16304 11756
rect 15427 11716 16304 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 16356 11716 17632 11744
rect 16356 11704 16362 11716
rect 13648 11648 13952 11676
rect 11517 11639 11575 11645
rect 8680 11580 9168 11608
rect 10888 11580 11560 11608
rect 4120 11568 4126 11580
rect 10888 11552 10916 11580
rect 2869 11543 2927 11549
rect 2869 11509 2881 11543
rect 2915 11540 2927 11543
rect 3418 11540 3424 11552
rect 2915 11512 3424 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 3418 11500 3424 11512
rect 3476 11540 3482 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 3476 11512 4997 11540
rect 3476 11500 3482 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 5994 11540 6000 11552
rect 5399 11512 6000 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6365 11543 6423 11549
rect 6365 11509 6377 11543
rect 6411 11540 6423 11543
rect 6638 11540 6644 11552
rect 6411 11512 6644 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 8570 11500 8576 11552
rect 8628 11500 8634 11552
rect 10594 11500 10600 11552
rect 10652 11500 10658 11552
rect 10870 11500 10876 11552
rect 10928 11500 10934 11552
rect 10962 11500 10968 11552
rect 11020 11500 11026 11552
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 11112 11512 11161 11540
rect 11112 11500 11118 11512
rect 11149 11509 11161 11512
rect 11195 11509 11207 11543
rect 11532 11540 11560 11580
rect 13924 11552 13952 11648
rect 17494 11636 17500 11688
rect 17552 11636 17558 11688
rect 17604 11676 17632 11716
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18509 11747 18567 11753
rect 18509 11744 18521 11747
rect 18196 11716 18521 11744
rect 18196 11704 18202 11716
rect 18509 11713 18521 11716
rect 18555 11713 18567 11747
rect 19794 11744 19800 11756
rect 18509 11707 18567 11713
rect 18616 11716 19800 11744
rect 18616 11676 18644 11716
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19944 11716 20361 11744
rect 19944 11704 19950 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 17604 11648 18644 11676
rect 19153 11679 19211 11685
rect 19153 11645 19165 11679
rect 19199 11676 19211 11679
rect 20070 11676 20076 11688
rect 19199 11648 20076 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 20162 11636 20168 11688
rect 20220 11676 20226 11688
rect 23768 11676 23796 11840
rect 24572 11815 24630 11821
rect 24572 11781 24584 11815
rect 24618 11812 24630 11815
rect 24964 11812 24992 11840
rect 24618 11784 24992 11812
rect 24618 11781 24630 11784
rect 24572 11775 24630 11781
rect 29638 11772 29644 11824
rect 29696 11812 29702 11824
rect 29825 11815 29883 11821
rect 29825 11812 29837 11815
rect 29696 11784 29837 11812
rect 29696 11772 29702 11784
rect 29825 11781 29837 11784
rect 29871 11781 29883 11815
rect 29825 11775 29883 11781
rect 31662 11772 31668 11824
rect 31720 11812 31726 11824
rect 35434 11812 35440 11824
rect 31720 11784 35440 11812
rect 31720 11772 31726 11784
rect 35434 11772 35440 11784
rect 35492 11772 35498 11824
rect 54012 11815 54070 11821
rect 54012 11781 54024 11815
rect 54058 11812 54070 11815
rect 54110 11812 54116 11824
rect 54058 11784 54116 11812
rect 54058 11781 54070 11784
rect 54012 11775 54070 11781
rect 54110 11772 54116 11784
rect 54168 11772 54174 11824
rect 24320 11716 25452 11744
rect 24320 11685 24348 11716
rect 20220 11648 23796 11676
rect 24305 11679 24363 11685
rect 20220 11636 20226 11648
rect 24305 11645 24317 11679
rect 24351 11645 24363 11679
rect 24305 11639 24363 11645
rect 25424 11620 25452 11716
rect 29178 11704 29184 11756
rect 29236 11704 29242 11756
rect 35066 11704 35072 11756
rect 35124 11704 35130 11756
rect 38102 11704 38108 11756
rect 38160 11704 38166 11756
rect 46934 11704 46940 11756
rect 46992 11704 46998 11756
rect 48705 11747 48763 11753
rect 48705 11713 48717 11747
rect 48751 11744 48763 11747
rect 48866 11744 48872 11756
rect 48751 11716 48872 11744
rect 48751 11713 48763 11716
rect 48705 11707 48763 11713
rect 48866 11704 48872 11716
rect 48924 11704 48930 11756
rect 48961 11747 49019 11753
rect 48961 11713 48973 11747
rect 49007 11744 49019 11747
rect 49970 11744 49976 11756
rect 49007 11716 49976 11744
rect 49007 11713 49019 11716
rect 48961 11707 49019 11713
rect 49970 11704 49976 11716
rect 50028 11704 50034 11756
rect 50430 11704 50436 11756
rect 50488 11704 50494 11756
rect 51166 11704 51172 11756
rect 51224 11704 51230 11756
rect 55416 11744 55444 11852
rect 56226 11840 56232 11852
rect 56284 11840 56290 11892
rect 57054 11840 57060 11892
rect 57112 11880 57118 11892
rect 57112 11852 57284 11880
rect 57112 11840 57118 11852
rect 53760 11716 55444 11744
rect 53760 11688 53788 11716
rect 56134 11704 56140 11756
rect 56192 11753 56198 11756
rect 57256 11753 57284 11852
rect 56192 11747 56241 11753
rect 56192 11713 56195 11747
rect 56229 11713 56241 11747
rect 56192 11707 56241 11713
rect 57241 11747 57299 11753
rect 57241 11713 57253 11747
rect 57287 11713 57299 11747
rect 57241 11707 57299 11713
rect 56192 11704 56198 11707
rect 58526 11704 58532 11756
rect 58584 11704 58590 11756
rect 26510 11636 26516 11688
rect 26568 11676 26574 11688
rect 28445 11679 28503 11685
rect 28445 11676 28457 11679
rect 26568 11648 28457 11676
rect 26568 11636 26574 11648
rect 28445 11645 28457 11648
rect 28491 11676 28503 11679
rect 28718 11676 28724 11688
rect 28491 11648 28724 11676
rect 28491 11645 28503 11648
rect 28445 11639 28503 11645
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 30098 11636 30104 11688
rect 30156 11676 30162 11688
rect 30193 11679 30251 11685
rect 30193 11676 30205 11679
rect 30156 11648 30205 11676
rect 30156 11636 30162 11648
rect 30193 11645 30205 11648
rect 30239 11645 30251 11679
rect 30193 11639 30251 11645
rect 31570 11636 31576 11688
rect 31628 11636 31634 11688
rect 33594 11636 33600 11688
rect 33652 11636 33658 11688
rect 33778 11636 33784 11688
rect 33836 11636 33842 11688
rect 34790 11636 34796 11688
rect 34848 11676 34854 11688
rect 36078 11676 36084 11688
rect 34848 11648 36084 11676
rect 34848 11636 34854 11648
rect 36078 11636 36084 11648
rect 36136 11636 36142 11688
rect 36170 11636 36176 11688
rect 36228 11636 36234 11688
rect 36354 11636 36360 11688
rect 36412 11636 36418 11688
rect 37826 11636 37832 11688
rect 37884 11636 37890 11688
rect 40862 11636 40868 11688
rect 40920 11636 40926 11688
rect 42978 11636 42984 11688
rect 43036 11636 43042 11688
rect 45462 11636 45468 11688
rect 45520 11636 45526 11688
rect 45646 11636 45652 11688
rect 45704 11636 45710 11688
rect 45922 11636 45928 11688
rect 45980 11636 45986 11688
rect 49602 11636 49608 11688
rect 49660 11636 49666 11688
rect 52454 11636 52460 11688
rect 52512 11636 52518 11688
rect 53282 11636 53288 11688
rect 53340 11636 53346 11688
rect 53742 11636 53748 11688
rect 53800 11636 53806 11688
rect 56045 11679 56103 11685
rect 56045 11676 56057 11679
rect 55600 11648 56057 11676
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 16850 11608 16856 11620
rect 14976 11580 16856 11608
rect 14976 11568 14982 11580
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 20438 11608 20444 11620
rect 16908 11580 20444 11608
rect 16908 11568 16914 11580
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 25406 11568 25412 11620
rect 25464 11608 25470 11620
rect 25464 11580 26004 11608
rect 25464 11568 25470 11580
rect 25976 11552 26004 11580
rect 32122 11568 32128 11620
rect 32180 11608 32186 11620
rect 32401 11611 32459 11617
rect 32401 11608 32413 11611
rect 32180 11580 32413 11608
rect 32180 11568 32186 11580
rect 32401 11577 32413 11580
rect 32447 11608 32459 11611
rect 32674 11608 32680 11620
rect 32447 11580 32680 11608
rect 32447 11577 32459 11580
rect 32401 11571 32459 11577
rect 32674 11568 32680 11580
rect 32732 11608 32738 11620
rect 32769 11611 32827 11617
rect 32769 11608 32781 11611
rect 32732 11580 32781 11608
rect 32732 11568 32738 11580
rect 32769 11577 32781 11580
rect 32815 11608 32827 11611
rect 34808 11608 34836 11636
rect 32815 11580 34836 11608
rect 32815 11577 32827 11580
rect 32769 11571 32827 11577
rect 36814 11568 36820 11620
rect 36872 11608 36878 11620
rect 37277 11611 37335 11617
rect 37277 11608 37289 11611
rect 36872 11580 37289 11608
rect 36872 11568 36878 11580
rect 37277 11577 37289 11580
rect 37323 11577 37335 11611
rect 45480 11608 45508 11636
rect 55600 11620 55628 11648
rect 56045 11645 56057 11648
rect 56091 11645 56103 11679
rect 56045 11639 56103 11645
rect 56321 11679 56379 11685
rect 56321 11645 56333 11679
rect 56367 11676 56379 11679
rect 56502 11676 56508 11688
rect 56367 11648 56508 11676
rect 56367 11645 56379 11648
rect 56321 11639 56379 11645
rect 56502 11636 56508 11648
rect 56560 11636 56566 11688
rect 57054 11636 57060 11688
rect 57112 11636 57118 11688
rect 47121 11611 47179 11617
rect 47121 11608 47133 11611
rect 45480 11580 47133 11608
rect 37277 11571 37335 11577
rect 47121 11577 47133 11580
rect 47167 11577 47179 11611
rect 47121 11571 47179 11577
rect 55582 11568 55588 11620
rect 55640 11568 55646 11620
rect 56594 11568 56600 11620
rect 56652 11608 56658 11620
rect 56870 11608 56876 11620
rect 56652 11580 56876 11608
rect 56652 11568 56658 11580
rect 56870 11568 56876 11580
rect 56928 11568 56934 11620
rect 11698 11540 11704 11552
rect 11532 11512 11704 11540
rect 11149 11503 11207 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13814 11540 13820 11552
rect 12943 11512 13820 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 13906 11500 13912 11552
rect 13964 11500 13970 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 14366 11540 14372 11552
rect 14139 11512 14372 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14608 11512 14657 11540
rect 14608 11500 14614 11512
rect 14645 11509 14657 11512
rect 14691 11540 14703 11543
rect 14734 11540 14740 11552
rect 14691 11512 14740 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 18322 11540 18328 11552
rect 18279 11512 18328 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 19576 11512 20545 11540
rect 19576 11500 19582 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 24486 11540 24492 11552
rect 21324 11512 24492 11540
rect 21324 11500 21330 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 25685 11543 25743 11549
rect 25685 11540 25697 11543
rect 25556 11512 25697 11540
rect 25556 11500 25562 11512
rect 25685 11509 25697 11512
rect 25731 11509 25743 11543
rect 25685 11503 25743 11509
rect 25958 11500 25964 11552
rect 26016 11500 26022 11552
rect 27706 11500 27712 11552
rect 27764 11540 27770 11552
rect 28077 11543 28135 11549
rect 28077 11540 28089 11543
rect 27764 11512 28089 11540
rect 27764 11500 27770 11512
rect 28077 11509 28089 11512
rect 28123 11509 28135 11543
rect 28077 11503 28135 11509
rect 28997 11543 29055 11549
rect 28997 11509 29009 11543
rect 29043 11540 29055 11543
rect 29086 11540 29092 11552
rect 29043 11512 29092 11540
rect 29043 11509 29055 11512
rect 28997 11503 29055 11509
rect 29086 11500 29092 11512
rect 29144 11540 29150 11552
rect 30558 11540 30564 11552
rect 29144 11512 30564 11540
rect 29144 11500 29150 11512
rect 30558 11500 30564 11512
rect 30616 11500 30622 11552
rect 30834 11500 30840 11552
rect 30892 11500 30898 11552
rect 31018 11500 31024 11552
rect 31076 11500 31082 11552
rect 33042 11500 33048 11552
rect 33100 11500 33106 11552
rect 34422 11500 34428 11552
rect 34480 11500 34486 11552
rect 35618 11500 35624 11552
rect 35676 11500 35682 11552
rect 36630 11500 36636 11552
rect 36688 11540 36694 11552
rect 37001 11543 37059 11549
rect 37001 11540 37013 11543
rect 36688 11512 37013 11540
rect 36688 11500 36694 11512
rect 37001 11509 37013 11512
rect 37047 11509 37059 11543
rect 37001 11503 37059 11509
rect 40034 11500 40040 11552
rect 40092 11540 40098 11552
rect 40313 11543 40371 11549
rect 40313 11540 40325 11543
rect 40092 11512 40325 11540
rect 40092 11500 40098 11512
rect 40313 11509 40325 11512
rect 40359 11509 40371 11543
rect 40313 11503 40371 11509
rect 42150 11500 42156 11552
rect 42208 11540 42214 11552
rect 42429 11543 42487 11549
rect 42429 11540 42441 11543
rect 42208 11512 42441 11540
rect 42208 11500 42214 11512
rect 42429 11509 42441 11512
rect 42475 11509 42487 11543
rect 42429 11503 42487 11509
rect 42794 11500 42800 11552
rect 42852 11540 42858 11552
rect 43714 11540 43720 11552
rect 42852 11512 43720 11540
rect 42852 11500 42858 11512
rect 43714 11500 43720 11512
rect 43772 11500 43778 11552
rect 45094 11500 45100 11552
rect 45152 11500 45158 11552
rect 45554 11500 45560 11552
rect 45612 11540 45618 11552
rect 46477 11543 46535 11549
rect 46477 11540 46489 11543
rect 45612 11512 46489 11540
rect 45612 11500 45618 11512
rect 46477 11509 46489 11512
rect 46523 11540 46535 11543
rect 47302 11540 47308 11552
rect 46523 11512 47308 11540
rect 46523 11509 46535 11512
rect 46477 11503 46535 11509
rect 47302 11500 47308 11512
rect 47360 11500 47366 11552
rect 48314 11500 48320 11552
rect 48372 11540 48378 11552
rect 49418 11540 49424 11552
rect 48372 11512 49424 11540
rect 48372 11500 48378 11512
rect 49418 11500 49424 11512
rect 49476 11540 49482 11552
rect 50249 11543 50307 11549
rect 50249 11540 50261 11543
rect 49476 11512 50261 11540
rect 49476 11500 49482 11512
rect 50249 11509 50261 11512
rect 50295 11509 50307 11543
rect 50249 11503 50307 11509
rect 50706 11500 50712 11552
rect 50764 11540 50770 11552
rect 50982 11540 50988 11552
rect 50764 11512 50988 11540
rect 50764 11500 50770 11512
rect 50982 11500 50988 11512
rect 51040 11500 51046 11552
rect 51902 11500 51908 11552
rect 51960 11500 51966 11552
rect 52730 11500 52736 11552
rect 52788 11500 52794 11552
rect 55401 11543 55459 11549
rect 55401 11509 55413 11543
rect 55447 11540 55459 11543
rect 56686 11540 56692 11552
rect 55447 11512 56692 11540
rect 55447 11509 55459 11512
rect 55401 11503 55459 11509
rect 56686 11500 56692 11512
rect 56744 11500 56750 11552
rect 57422 11500 57428 11552
rect 57480 11540 57486 11552
rect 58345 11543 58403 11549
rect 58345 11540 58357 11543
rect 57480 11512 58357 11540
rect 57480 11500 57486 11512
rect 58345 11509 58357 11512
rect 58391 11509 58403 11543
rect 58345 11503 58403 11509
rect 1104 11450 58880 11472
rect 1104 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 22616 11450
rect 22668 11398 22680 11450
rect 22732 11398 22744 11450
rect 22796 11398 22808 11450
rect 22860 11398 22872 11450
rect 22924 11398 37060 11450
rect 37112 11398 37124 11450
rect 37176 11398 37188 11450
rect 37240 11398 37252 11450
rect 37304 11398 37316 11450
rect 37368 11398 51504 11450
rect 51556 11398 51568 11450
rect 51620 11398 51632 11450
rect 51684 11398 51696 11450
rect 51748 11398 51760 11450
rect 51812 11398 58880 11450
rect 1104 11376 58880 11398
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4798 11336 4804 11348
rect 4387 11308 4804 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7984 11308 8033 11336
rect 7984 11296 7990 11308
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 8021 11299 8079 11305
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9950 11336 9956 11348
rect 8987 11308 9956 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10336 11308 11560 11336
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 2866 11268 2872 11280
rect 2363 11240 2872 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 7576 11268 7604 11296
rect 4488 11240 4660 11268
rect 4488 11228 4494 11240
rect 3068 11172 4292 11200
rect 2498 11092 2504 11144
rect 2556 11092 2562 11144
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 3068 11141 3096 11172
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3418 11132 3424 11144
rect 3283 11104 3424 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3786 11092 3792 11144
rect 3844 11141 3850 11144
rect 3844 11135 3867 11141
rect 3855 11101 3867 11135
rect 3844 11095 3867 11101
rect 3844 11092 3850 11095
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4062 11092 4068 11144
rect 4120 11092 4126 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4264 11132 4292 11172
rect 4264 11104 4384 11132
rect 4157 11095 4215 11101
rect 2685 11067 2743 11073
rect 2685 11033 2697 11067
rect 2731 11033 2743 11067
rect 3436 11064 3464 11092
rect 4172 11064 4200 11095
rect 3436 11036 4200 11064
rect 2685 11027 2743 11033
rect 2700 10996 2728 11027
rect 2866 10996 2872 11008
rect 2700 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10996 3479 10999
rect 3510 10996 3516 11008
rect 3467 10968 3516 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4246 10996 4252 11008
rect 3844 10968 4252 10996
rect 3844 10956 3850 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4356 10996 4384 11104
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4632 11141 4660 11240
rect 7300 11240 7604 11268
rect 7300 11209 7328 11240
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 7742 11200 7748 11212
rect 7515 11172 7748 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 7852 11172 8585 11200
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 6972 11104 7205 11132
rect 6972 11092 6978 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7852 11073 7880 11172
rect 8573 11169 8585 11172
rect 8619 11169 8631 11203
rect 10336 11200 10364 11308
rect 8573 11163 8631 11169
rect 10244 11172 10364 11200
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8938 11132 8944 11144
rect 8435 11104 8944 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 10244 11132 10272 11172
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 11532 11200 11560 11308
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11756 11308 12434 11336
rect 11756 11296 11762 11308
rect 12406 11268 12434 11308
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 13964 11308 17540 11336
rect 13964 11296 13970 11308
rect 13354 11268 13360 11280
rect 12406 11240 13360 11268
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 16206 11268 16212 11280
rect 15252 11240 16212 11268
rect 15252 11228 15258 11240
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 16850 11228 16856 11280
rect 16908 11228 16914 11280
rect 17405 11271 17463 11277
rect 17405 11237 17417 11271
rect 17451 11237 17463 11271
rect 17512 11268 17540 11308
rect 18414 11296 18420 11348
rect 18472 11296 18478 11348
rect 23474 11336 23480 11348
rect 18524 11308 23480 11336
rect 18524 11268 18552 11308
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 23658 11296 23664 11348
rect 23716 11296 23722 11348
rect 24486 11296 24492 11348
rect 24544 11336 24550 11348
rect 24857 11339 24915 11345
rect 24857 11336 24869 11339
rect 24544 11308 24869 11336
rect 24544 11296 24550 11308
rect 24857 11305 24869 11308
rect 24903 11305 24915 11339
rect 24857 11299 24915 11305
rect 26789 11339 26847 11345
rect 26789 11305 26801 11339
rect 26835 11336 26847 11339
rect 27522 11336 27528 11348
rect 26835 11308 27528 11336
rect 26835 11305 26847 11308
rect 26789 11299 26847 11305
rect 27522 11296 27528 11308
rect 27580 11296 27586 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 27632 11308 29929 11336
rect 17512 11240 18552 11268
rect 17405 11231 17463 11237
rect 10560 11172 11100 11200
rect 10560 11160 10566 11172
rect 8996 11104 10272 11132
rect 8996 11092 9002 11104
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 11072 11141 11100 11172
rect 11210 11172 11560 11200
rect 11609 11203 11667 11209
rect 11210 11141 11238 11172
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11698 11200 11704 11212
rect 11655 11172 11704 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12069 11203 12127 11209
rect 12069 11169 12081 11203
rect 12115 11200 12127 11203
rect 13538 11200 13544 11212
rect 12115 11172 13544 11200
rect 12115 11169 12127 11172
rect 12069 11163 12127 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16623 11172 16773 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 16761 11169 16773 11172
rect 16807 11200 16819 11203
rect 16868 11200 16896 11228
rect 16807 11172 16896 11200
rect 17420 11200 17448 11231
rect 21450 11228 21456 11280
rect 21508 11228 21514 11280
rect 22370 11268 22376 11280
rect 21560 11240 22376 11268
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 17420 11172 17509 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 17497 11169 17509 11172
rect 17543 11169 17555 11203
rect 21468 11200 21496 11228
rect 17497 11163 17555 11169
rect 19306 11172 21496 11200
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11195 11135 11253 11141
rect 11195 11101 11207 11135
rect 11241 11101 11253 11135
rect 11195 11095 11253 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 11940 11104 12265 11132
rect 11940 11092 11946 11104
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7340 11036 7849 11064
rect 7340 11024 7346 11036
rect 7837 11033 7849 11036
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 8481 11067 8539 11073
rect 8481 11033 8493 11067
rect 8527 11064 8539 11067
rect 9950 11064 9956 11076
rect 8527 11036 9956 11064
rect 8527 11033 8539 11036
rect 8481 11027 8539 11033
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10076 11067 10134 11073
rect 10076 11033 10088 11067
rect 10122 11064 10134 11067
rect 10226 11064 10232 11076
rect 10122 11036 10232 11064
rect 10122 11033 10134 11036
rect 10076 11027 10134 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 12360 11064 12388 11095
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 12584 11104 13185 11132
rect 12584 11092 12590 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 19306 11132 19334 11172
rect 15304 11104 19334 11132
rect 15304 11064 15332 11104
rect 20346 11092 20352 11144
rect 20404 11092 20410 11144
rect 20438 11092 20444 11144
rect 20496 11132 20502 11144
rect 20496 11104 20852 11132
rect 20496 11092 20502 11104
rect 12360 11036 15332 11064
rect 4433 10999 4491 11005
rect 4433 10996 4445 10999
rect 4356 10968 4445 10996
rect 4433 10965 4445 10968
rect 4479 10965 4491 10999
rect 4433 10959 4491 10965
rect 6822 10956 6828 11008
rect 6880 10956 6886 11008
rect 10962 10956 10968 11008
rect 11020 10996 11026 11008
rect 11238 10996 11244 11008
rect 11020 10968 11244 10996
rect 11020 10956 11026 10968
rect 11238 10956 11244 10968
rect 11296 10996 11302 11008
rect 12360 10996 12388 11036
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 17000 11036 17724 11064
rect 17000 11024 17006 11036
rect 17696 11008 17724 11036
rect 19794 11024 19800 11076
rect 19852 11024 19858 11076
rect 20824 11064 20852 11104
rect 21174 11092 21180 11144
rect 21232 11092 21238 11144
rect 21450 11092 21456 11144
rect 21508 11092 21514 11144
rect 21560 11064 21588 11240
rect 22370 11228 22376 11240
rect 22428 11228 22434 11280
rect 23290 11228 23296 11280
rect 23348 11268 23354 11280
rect 23676 11268 23704 11296
rect 27632 11268 27660 11308
rect 29917 11305 29929 11308
rect 29963 11305 29975 11339
rect 29917 11299 29975 11305
rect 23348 11240 23612 11268
rect 23676 11240 27660 11268
rect 28629 11271 28687 11277
rect 23348 11228 23354 11240
rect 23584 11209 23612 11240
rect 28629 11237 28641 11271
rect 28675 11237 28687 11271
rect 28629 11231 28687 11237
rect 23569 11203 23627 11209
rect 20456 11036 20760 11064
rect 20824 11036 21588 11064
rect 21928 11172 23520 11200
rect 11296 10968 12388 10996
rect 11296 10956 11302 10968
rect 14366 10956 14372 11008
rect 14424 10956 14430 11008
rect 14550 10956 14556 11008
rect 14608 10956 14614 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 17037 10999 17095 11005
rect 17037 10996 17049 10999
rect 15344 10968 17049 10996
rect 15344 10956 15350 10968
rect 17037 10965 17049 10968
rect 17083 10996 17095 10999
rect 17126 10996 17132 11008
rect 17083 10968 17132 10996
rect 17083 10965 17095 10968
rect 17037 10959 17095 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17678 10956 17684 11008
rect 17736 10956 17742 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 18012 10968 18153 10996
rect 18012 10956 18018 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 20456 10996 20484 11036
rect 19300 10968 20484 10996
rect 19300 10956 19306 10968
rect 20530 10956 20536 11008
rect 20588 10996 20594 11008
rect 20625 10999 20683 11005
rect 20625 10996 20637 10999
rect 20588 10968 20637 10996
rect 20588 10956 20594 10968
rect 20625 10965 20637 10968
rect 20671 10965 20683 10999
rect 20732 10996 20760 11036
rect 21542 10996 21548 11008
rect 20732 10968 21548 10996
rect 20625 10959 20683 10965
rect 21542 10956 21548 10968
rect 21600 10996 21606 11008
rect 21928 10996 21956 11172
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 23492 11132 23520 11172
rect 23569 11169 23581 11203
rect 23615 11169 23627 11203
rect 23569 11163 23627 11169
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11200 28595 11203
rect 28644 11200 28672 11231
rect 28718 11228 28724 11280
rect 28776 11228 28782 11280
rect 28902 11228 28908 11280
rect 28960 11268 28966 11280
rect 29932 11268 29960 11299
rect 30098 11296 30104 11348
rect 30156 11296 30162 11348
rect 37553 11339 37611 11345
rect 37553 11305 37565 11339
rect 37599 11336 37611 11339
rect 37826 11336 37832 11348
rect 37599 11308 37832 11336
rect 37599 11305 37611 11308
rect 37553 11299 37611 11305
rect 37826 11296 37832 11308
rect 37884 11296 37890 11348
rect 41233 11339 41291 11345
rect 41233 11305 41245 11339
rect 41279 11336 41291 11339
rect 42978 11336 42984 11348
rect 41279 11308 42984 11336
rect 41279 11305 41291 11308
rect 41233 11299 41291 11305
rect 42978 11296 42984 11308
rect 43036 11296 43042 11348
rect 44450 11296 44456 11348
rect 44508 11336 44514 11348
rect 44634 11336 44640 11348
rect 44508 11308 44640 11336
rect 44508 11296 44514 11308
rect 44634 11296 44640 11308
rect 44692 11296 44698 11348
rect 45189 11339 45247 11345
rect 45189 11305 45201 11339
rect 45235 11336 45247 11339
rect 45646 11336 45652 11348
rect 45235 11308 45652 11336
rect 45235 11305 45247 11308
rect 45189 11299 45247 11305
rect 45646 11296 45652 11308
rect 45704 11296 45710 11348
rect 46293 11339 46351 11345
rect 46293 11305 46305 11339
rect 46339 11336 46351 11339
rect 46474 11336 46480 11348
rect 46339 11308 46480 11336
rect 46339 11305 46351 11308
rect 46293 11299 46351 11305
rect 35253 11271 35311 11277
rect 28960 11240 29868 11268
rect 29932 11240 30135 11268
rect 28960 11228 28966 11240
rect 28583 11172 28672 11200
rect 28736 11200 28764 11228
rect 29181 11203 29239 11209
rect 29181 11200 29193 11203
rect 28736 11172 29193 11200
rect 28583 11169 28595 11172
rect 28537 11163 28595 11169
rect 29181 11169 29193 11172
rect 29227 11169 29239 11203
rect 29181 11163 29239 11169
rect 25685 11135 25743 11141
rect 25685 11132 25697 11135
rect 23492 11104 25697 11132
rect 25685 11101 25697 11104
rect 25731 11132 25743 11135
rect 26418 11132 26424 11144
rect 25731 11104 26424 11132
rect 25731 11101 25743 11104
rect 25685 11095 25743 11101
rect 26418 11092 26424 11104
rect 26476 11092 26482 11144
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 22741 11067 22799 11073
rect 22741 11033 22753 11067
rect 22787 11064 22799 11067
rect 23198 11064 23204 11076
rect 22787 11036 23204 11064
rect 22787 11033 22799 11036
rect 22741 11027 22799 11033
rect 23198 11024 23204 11036
rect 23256 11024 23262 11076
rect 26510 11064 26516 11076
rect 23860 11036 26516 11064
rect 21600 10968 21956 10996
rect 21600 10956 21606 10968
rect 22002 10956 22008 11008
rect 22060 10956 22066 11008
rect 22922 10956 22928 11008
rect 22980 10956 22986 11008
rect 23658 10956 23664 11008
rect 23716 10996 23722 11008
rect 23860 11005 23888 11036
rect 26510 11024 26516 11036
rect 26568 11024 26574 11076
rect 26694 11024 26700 11076
rect 26752 11024 26758 11076
rect 27890 11024 27896 11076
rect 27948 11024 27954 11076
rect 29089 11067 29147 11073
rect 29089 11033 29101 11067
rect 29135 11064 29147 11067
rect 29178 11064 29184 11076
rect 29135 11036 29184 11064
rect 29135 11033 29147 11036
rect 29089 11027 29147 11033
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 23845 10999 23903 11005
rect 23845 10996 23857 10999
rect 23716 10968 23857 10996
rect 23716 10956 23722 10968
rect 23845 10965 23857 10968
rect 23891 10965 23903 10999
rect 23845 10959 23903 10965
rect 27157 10999 27215 11005
rect 27157 10965 27169 10999
rect 27203 10996 27215 10999
rect 27246 10996 27252 11008
rect 27203 10968 27252 10996
rect 27203 10965 27215 10968
rect 27157 10959 27215 10965
rect 27246 10956 27252 10968
rect 27304 10956 27310 11008
rect 28994 10956 29000 11008
rect 29052 10956 29058 11008
rect 29840 10996 29868 11240
rect 30107 11132 30135 11240
rect 35253 11237 35265 11271
rect 35299 11268 35311 11271
rect 35526 11268 35532 11280
rect 35299 11240 35532 11268
rect 35299 11237 35311 11240
rect 35253 11231 35311 11237
rect 35526 11228 35532 11240
rect 35584 11228 35590 11280
rect 37461 11271 37519 11277
rect 37461 11237 37473 11271
rect 37507 11268 37519 11271
rect 37642 11268 37648 11280
rect 37507 11240 37648 11268
rect 37507 11237 37519 11240
rect 37461 11231 37519 11237
rect 37642 11228 37648 11240
rect 37700 11228 37706 11280
rect 43441 11271 43499 11277
rect 43441 11237 43453 11271
rect 43487 11268 43499 11271
rect 44174 11268 44180 11280
rect 43487 11240 44180 11268
rect 43487 11237 43499 11240
rect 43441 11231 43499 11237
rect 44174 11228 44180 11240
rect 44232 11228 44238 11280
rect 30742 11160 30748 11212
rect 30800 11160 30806 11212
rect 31662 11160 31668 11212
rect 31720 11160 31726 11212
rect 32398 11200 32404 11212
rect 31772 11172 32404 11200
rect 30929 11135 30987 11141
rect 30929 11132 30941 11135
rect 30107 11104 30941 11132
rect 30929 11101 30941 11104
rect 30975 11101 30987 11135
rect 30929 11095 30987 11101
rect 30466 11024 30472 11076
rect 30524 11024 30530 11076
rect 30561 11067 30619 11073
rect 30561 11033 30573 11067
rect 30607 11064 30619 11067
rect 31018 11064 31024 11076
rect 30607 11036 31024 11064
rect 30607 11033 30619 11036
rect 30561 11027 30619 11033
rect 31018 11024 31024 11036
rect 31076 11064 31082 11076
rect 31772 11064 31800 11172
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 33597 11203 33655 11209
rect 33597 11169 33609 11203
rect 33643 11200 33655 11203
rect 34790 11200 34796 11212
rect 33643 11172 34796 11200
rect 33643 11169 33655 11172
rect 33597 11163 33655 11169
rect 34790 11160 34796 11172
rect 34848 11160 34854 11212
rect 35434 11160 35440 11212
rect 35492 11200 35498 11212
rect 35805 11203 35863 11209
rect 35805 11200 35817 11203
rect 35492 11172 35817 11200
rect 35492 11160 35498 11172
rect 35805 11169 35817 11172
rect 35851 11169 35863 11203
rect 35805 11163 35863 11169
rect 37734 11160 37740 11212
rect 37792 11200 37798 11212
rect 38105 11203 38163 11209
rect 38105 11200 38117 11203
rect 37792 11172 38117 11200
rect 37792 11160 37798 11172
rect 38105 11169 38117 11172
rect 38151 11200 38163 11203
rect 38151 11172 39804 11200
rect 38151 11169 38163 11172
rect 38105 11163 38163 11169
rect 33781 11135 33839 11141
rect 33781 11132 33793 11135
rect 31076 11036 31800 11064
rect 32140 11104 33793 11132
rect 31076 11024 31082 11036
rect 32140 10996 32168 11104
rect 33781 11101 33793 11104
rect 33827 11132 33839 11135
rect 33827 11104 34468 11132
rect 33827 11101 33839 11104
rect 33781 11095 33839 11101
rect 33352 11067 33410 11073
rect 33352 11033 33364 11067
rect 33398 11064 33410 11067
rect 33502 11064 33508 11076
rect 33398 11036 33508 11064
rect 33398 11033 33410 11036
rect 33352 11027 33410 11033
rect 33502 11024 33508 11036
rect 33560 11024 33566 11076
rect 34054 11024 34060 11076
rect 34112 11064 34118 11076
rect 34330 11064 34336 11076
rect 34112 11036 34336 11064
rect 34112 11024 34118 11036
rect 34330 11024 34336 11036
rect 34388 11024 34394 11076
rect 34440 11064 34468 11104
rect 36078 11092 36084 11144
rect 36136 11132 36142 11144
rect 37550 11132 37556 11144
rect 36136 11104 37556 11132
rect 36136 11092 36142 11104
rect 37550 11092 37556 11104
rect 37608 11092 37614 11144
rect 39022 11092 39028 11144
rect 39080 11092 39086 11144
rect 39776 11132 39804 11172
rect 39850 11160 39856 11212
rect 39908 11160 39914 11212
rect 41598 11160 41604 11212
rect 41656 11200 41662 11212
rect 42058 11200 42064 11212
rect 41656 11172 42064 11200
rect 41656 11160 41662 11172
rect 42058 11160 42064 11172
rect 42116 11160 42122 11212
rect 45833 11203 45891 11209
rect 45833 11169 45845 11203
rect 45879 11200 45891 11203
rect 46308 11200 46336 11299
rect 46474 11296 46480 11308
rect 46532 11296 46538 11348
rect 48130 11336 48136 11348
rect 46768 11308 48136 11336
rect 45879 11172 46336 11200
rect 46768 11200 46796 11308
rect 48130 11296 48136 11308
rect 48188 11296 48194 11348
rect 48774 11296 48780 11348
rect 48832 11296 48838 11348
rect 48866 11296 48872 11348
rect 48924 11296 48930 11348
rect 49145 11339 49203 11345
rect 49145 11305 49157 11339
rect 49191 11336 49203 11339
rect 49602 11336 49608 11348
rect 49191 11308 49608 11336
rect 49191 11305 49203 11308
rect 49145 11299 49203 11305
rect 49602 11296 49608 11308
rect 49660 11296 49666 11348
rect 50522 11296 50528 11348
rect 50580 11336 50586 11348
rect 50709 11339 50767 11345
rect 50709 11336 50721 11339
rect 50580 11308 50721 11336
rect 50580 11296 50586 11308
rect 50709 11305 50721 11308
rect 50755 11305 50767 11339
rect 50709 11299 50767 11305
rect 52362 11296 52368 11348
rect 52420 11296 52426 11348
rect 52454 11296 52460 11348
rect 52512 11296 52518 11348
rect 53466 11296 53472 11348
rect 53524 11296 53530 11348
rect 47670 11228 47676 11280
rect 47728 11268 47734 11280
rect 48222 11268 48228 11280
rect 47728 11240 48228 11268
rect 47728 11228 47734 11240
rect 48222 11228 48228 11240
rect 48280 11228 48286 11280
rect 47123 11203 47181 11209
rect 47123 11200 47135 11203
rect 46768 11172 47135 11200
rect 45879 11169 45891 11172
rect 45833 11163 45891 11169
rect 47123 11169 47135 11172
rect 47169 11169 47181 11203
rect 47123 11163 47181 11169
rect 47762 11160 47768 11212
rect 47820 11200 47826 11212
rect 48317 11203 48375 11209
rect 48317 11200 48329 11203
rect 47820 11172 48329 11200
rect 47820 11160 47826 11172
rect 48317 11169 48329 11172
rect 48363 11169 48375 11203
rect 48317 11163 48375 11169
rect 48590 11160 48596 11212
rect 48648 11160 48654 11212
rect 39776 11104 40356 11132
rect 34885 11067 34943 11073
rect 34885 11064 34897 11067
rect 34440 11036 34897 11064
rect 34885 11033 34897 11036
rect 34931 11033 34943 11067
rect 34885 11027 34943 11033
rect 35621 11067 35679 11073
rect 35621 11033 35633 11067
rect 35667 11064 35679 11067
rect 35986 11064 35992 11076
rect 35667 11036 35992 11064
rect 35667 11033 35679 11036
rect 35621 11027 35679 11033
rect 35986 11024 35992 11036
rect 36044 11024 36050 11076
rect 36348 11067 36406 11073
rect 36348 11033 36360 11067
rect 36394 11064 36406 11067
rect 36814 11064 36820 11076
rect 36394 11036 36820 11064
rect 36394 11033 36406 11036
rect 36348 11027 36406 11033
rect 36814 11024 36820 11036
rect 36872 11024 36878 11076
rect 38378 11024 38384 11076
rect 38436 11024 38442 11076
rect 40120 11067 40178 11073
rect 40120 11033 40132 11067
rect 40166 11064 40178 11067
rect 40218 11064 40224 11076
rect 40166 11036 40224 11064
rect 40166 11033 40178 11036
rect 40120 11027 40178 11033
rect 40218 11024 40224 11036
rect 40276 11024 40282 11076
rect 40328 11064 40356 11104
rect 41322 11092 41328 11144
rect 41380 11092 41386 11144
rect 44082 11092 44088 11144
rect 44140 11092 44146 11144
rect 45554 11092 45560 11144
rect 45612 11092 45618 11144
rect 47277 11141 47283 11144
rect 47259 11135 47283 11141
rect 47259 11101 47271 11135
rect 47259 11095 47283 11101
rect 47277 11092 47283 11095
rect 47335 11092 47341 11144
rect 47394 11092 47400 11144
rect 47452 11092 47458 11144
rect 48792 11141 48820 11296
rect 48884 11268 48912 11296
rect 49237 11271 49295 11277
rect 49237 11268 49249 11271
rect 48884 11240 49249 11268
rect 49237 11237 49249 11240
rect 49283 11237 49295 11271
rect 49237 11231 49295 11237
rect 52914 11160 52920 11212
rect 52972 11160 52978 11212
rect 53101 11203 53159 11209
rect 53101 11169 53113 11203
rect 53147 11200 53159 11203
rect 53484 11200 53512 11296
rect 57609 11271 57667 11277
rect 57609 11237 57621 11271
rect 57655 11268 57667 11271
rect 58434 11268 58440 11280
rect 57655 11240 58440 11268
rect 57655 11237 57667 11240
rect 57609 11231 57667 11237
rect 58434 11228 58440 11240
rect 58492 11228 58498 11280
rect 53147 11172 53512 11200
rect 53147 11169 53159 11172
rect 53101 11163 53159 11169
rect 53742 11160 53748 11212
rect 53800 11160 53806 11212
rect 56226 11160 56232 11212
rect 56284 11160 56290 11212
rect 48133 11135 48191 11141
rect 48133 11101 48145 11135
rect 48179 11132 48191 11135
rect 48777 11135 48835 11141
rect 48777 11132 48789 11135
rect 48179 11104 48789 11132
rect 48179 11101 48191 11104
rect 48133 11095 48191 11101
rect 48777 11101 48789 11104
rect 48823 11101 48835 11135
rect 48777 11095 48835 11101
rect 49694 11092 49700 11144
rect 49752 11132 49758 11144
rect 49789 11135 49847 11141
rect 49789 11132 49801 11135
rect 49752 11104 49801 11132
rect 49752 11092 49758 11104
rect 49789 11101 49801 11104
rect 49835 11101 49847 11135
rect 49789 11095 49847 11101
rect 50985 11135 51043 11141
rect 50985 11101 50997 11135
rect 51031 11132 51043 11135
rect 53760 11132 53788 11160
rect 51031 11104 53788 11132
rect 51031 11101 51043 11104
rect 50985 11095 51043 11101
rect 41782 11064 41788 11076
rect 40328 11036 41788 11064
rect 41782 11024 41788 11036
rect 41840 11024 41846 11076
rect 42328 11067 42386 11073
rect 42328 11033 42340 11067
rect 42374 11064 42386 11067
rect 43898 11064 43904 11076
rect 42374 11036 43904 11064
rect 42374 11033 42386 11036
rect 42328 11027 42386 11033
rect 43898 11024 43904 11036
rect 43956 11024 43962 11076
rect 46474 11024 46480 11076
rect 46532 11024 46538 11076
rect 51184 11008 51212 11104
rect 55858 11092 55864 11144
rect 55916 11092 55922 11144
rect 57330 11092 57336 11144
rect 57388 11132 57394 11144
rect 58253 11135 58311 11141
rect 58253 11132 58265 11135
rect 57388 11104 58265 11132
rect 57388 11092 57394 11104
rect 58253 11101 58265 11104
rect 58299 11101 58311 11135
rect 58253 11095 58311 11101
rect 51252 11067 51310 11073
rect 51252 11033 51264 11067
rect 51298 11064 51310 11067
rect 51902 11064 51908 11076
rect 51298 11036 51908 11064
rect 51298 11033 51310 11036
rect 51252 11027 51310 11033
rect 51902 11024 51908 11036
rect 51960 11024 51966 11076
rect 54012 11067 54070 11073
rect 54012 11033 54024 11067
rect 54058 11064 54070 11067
rect 55309 11067 55367 11073
rect 55309 11064 55321 11067
rect 54058 11036 55321 11064
rect 54058 11033 54070 11036
rect 54012 11027 54070 11033
rect 55309 11033 55321 11036
rect 55355 11033 55367 11067
rect 55309 11027 55367 11033
rect 56496 11067 56554 11073
rect 56496 11033 56508 11067
rect 56542 11064 56554 11067
rect 57701 11067 57759 11073
rect 57701 11064 57713 11067
rect 56542 11036 57713 11064
rect 56542 11033 56554 11036
rect 56496 11027 56554 11033
rect 57701 11033 57713 11036
rect 57747 11033 57759 11067
rect 57701 11027 57759 11033
rect 29840 10968 32168 10996
rect 32214 10956 32220 11008
rect 32272 10956 32278 11008
rect 35713 10999 35771 11005
rect 35713 10965 35725 10999
rect 35759 10996 35771 10999
rect 35802 10996 35808 11008
rect 35759 10968 35808 10996
rect 35759 10965 35771 10968
rect 35713 10959 35771 10965
rect 35802 10956 35808 10968
rect 35860 10996 35866 11008
rect 37918 10996 37924 11008
rect 35860 10968 37924 10996
rect 35860 10956 35866 10968
rect 37918 10956 37924 10968
rect 37976 10956 37982 11008
rect 38010 10956 38016 11008
rect 38068 10956 38074 11008
rect 39298 10956 39304 11008
rect 39356 10956 39362 11008
rect 41966 10956 41972 11008
rect 42024 10956 42030 11008
rect 43530 10956 43536 11008
rect 43588 10956 43594 11008
rect 45646 10956 45652 11008
rect 45704 10956 45710 11008
rect 46566 10956 46572 11008
rect 46624 10996 46630 11008
rect 47118 10996 47124 11008
rect 46624 10968 47124 10996
rect 46624 10956 46630 10968
rect 47118 10956 47124 10968
rect 47176 10956 47182 11008
rect 48682 10956 48688 11008
rect 48740 10956 48746 11008
rect 51166 10956 51172 11008
rect 51224 10956 51230 11008
rect 52822 10956 52828 11008
rect 52880 10956 52886 11008
rect 55122 10956 55128 11008
rect 55180 10956 55186 11008
rect 1104 10906 59040 10928
rect 1104 10854 15394 10906
rect 15446 10854 15458 10906
rect 15510 10854 15522 10906
rect 15574 10854 15586 10906
rect 15638 10854 15650 10906
rect 15702 10854 29838 10906
rect 29890 10854 29902 10906
rect 29954 10854 29966 10906
rect 30018 10854 30030 10906
rect 30082 10854 30094 10906
rect 30146 10854 44282 10906
rect 44334 10854 44346 10906
rect 44398 10854 44410 10906
rect 44462 10854 44474 10906
rect 44526 10854 44538 10906
rect 44590 10854 58726 10906
rect 58778 10854 58790 10906
rect 58842 10854 58854 10906
rect 58906 10854 58918 10906
rect 58970 10854 58982 10906
rect 59034 10854 59040 10906
rect 1104 10832 59040 10854
rect 2774 10752 2780 10804
rect 2832 10752 2838 10804
rect 2866 10752 2872 10804
rect 2924 10752 2930 10804
rect 3881 10795 3939 10801
rect 3881 10761 3893 10795
rect 3927 10792 3939 10795
rect 3970 10792 3976 10804
rect 3927 10764 3976 10792
rect 3927 10761 3939 10764
rect 3881 10755 3939 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10761 4215 10795
rect 4157 10755 4215 10761
rect 2884 10724 2912 10752
rect 2884 10696 3740 10724
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 2823 10628 3065 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 3053 10625 3065 10628
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 2608 10588 2636 10619
rect 2608 10560 2774 10588
rect 2746 10452 2774 10560
rect 3068 10532 3096 10619
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3510 10656 3516 10668
rect 3384 10628 3516 10656
rect 3384 10616 3390 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3712 10665 3740 10696
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 4172 10724 4200 10755
rect 4246 10752 4252 10804
rect 4304 10752 4310 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7466 10792 7472 10804
rect 7423 10764 7472 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7742 10752 7748 10804
rect 7800 10752 7806 10804
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10594 10792 10600 10804
rect 10275 10764 10600 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 11020 10764 14473 10792
rect 11020 10752 11026 10764
rect 3844 10696 4200 10724
rect 8288 10727 8346 10733
rect 3844 10684 3850 10696
rect 8288 10693 8300 10727
rect 8334 10724 8346 10727
rect 8570 10724 8576 10736
rect 8334 10696 8576 10724
rect 8334 10693 8346 10696
rect 8288 10687 8346 10693
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 9968 10724 9996 10752
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 9968 10696 10333 10724
rect 10321 10693 10333 10696
rect 10367 10724 10379 10727
rect 11698 10724 11704 10736
rect 10367 10696 11704 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 11698 10684 11704 10696
rect 11756 10724 11762 10736
rect 13633 10727 13691 10733
rect 13633 10724 13645 10727
rect 11756 10696 13645 10724
rect 11756 10684 11762 10696
rect 13633 10693 13645 10696
rect 13679 10693 13691 10727
rect 13633 10687 13691 10693
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3743 10628 3985 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3200 10560 3433 10588
rect 3200 10548 3206 10560
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 3786 10588 3792 10600
rect 3651 10560 3792 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 3050 10480 3056 10532
rect 3108 10480 3114 10532
rect 3436 10520 3464 10551
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 4080 10520 4108 10619
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4212 10628 4353 10656
rect 4212 10616 4218 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 6822 10616 6828 10668
rect 6880 10616 6886 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 11330 10656 11336 10668
rect 10652 10628 11336 10656
rect 10652 10616 10658 10628
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 11784 10659 11842 10665
rect 11784 10625 11796 10659
rect 11830 10656 11842 10659
rect 12066 10656 12072 10668
rect 11830 10628 12072 10656
rect 11830 10625 11842 10628
rect 11784 10619 11842 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 8018 10548 8024 10600
rect 8076 10548 8082 10600
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9824 10560 10149 10588
rect 9824 10548 9830 10560
rect 10137 10557 10149 10560
rect 10183 10588 10195 10591
rect 10962 10588 10968 10600
rect 10183 10560 10968 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11422 10588 11428 10600
rect 11204 10560 11428 10588
rect 11204 10548 11210 10560
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 13725 10591 13783 10597
rect 13725 10588 13737 10591
rect 11517 10551 11575 10557
rect 12544 10560 13737 10588
rect 3436 10492 4108 10520
rect 9858 10480 9864 10532
rect 9916 10520 9922 10532
rect 10318 10520 10324 10532
rect 9916 10492 10324 10520
rect 9916 10480 9922 10492
rect 10318 10480 10324 10492
rect 10376 10520 10382 10532
rect 11532 10520 11560 10551
rect 10376 10492 11560 10520
rect 10376 10480 10382 10492
rect 10980 10464 11008 10492
rect 12544 10464 12572 10560
rect 13725 10557 13737 10560
rect 13771 10557 13783 10591
rect 14292 10588 14320 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 15194 10792 15200 10804
rect 14691 10764 15200 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 17494 10792 17500 10804
rect 16715 10764 17500 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 19518 10752 19524 10804
rect 19576 10752 19582 10804
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 20346 10792 20352 10804
rect 19935 10764 20352 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 21450 10752 21456 10804
rect 21508 10792 21514 10804
rect 21637 10795 21695 10801
rect 21637 10792 21649 10795
rect 21508 10764 21649 10792
rect 21508 10752 21514 10764
rect 21637 10761 21649 10764
rect 21683 10761 21695 10795
rect 21637 10755 21695 10761
rect 26329 10795 26387 10801
rect 26329 10761 26341 10795
rect 26375 10792 26387 10795
rect 27982 10792 27988 10804
rect 26375 10764 27988 10792
rect 26375 10761 26387 10764
rect 26329 10755 26387 10761
rect 27982 10752 27988 10764
rect 28040 10752 28046 10804
rect 30392 10764 32168 10792
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 14424 10696 15761 10724
rect 14424 10684 14430 10696
rect 15749 10693 15761 10696
rect 15795 10724 15807 10727
rect 27614 10724 27620 10736
rect 15795 10696 18092 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 15010 10616 15016 10668
rect 15068 10616 15074 10668
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 16485 10659 16543 10665
rect 16485 10656 16497 10659
rect 15151 10628 16497 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 16485 10625 16497 10628
rect 16531 10656 16543 10659
rect 16758 10656 16764 10668
rect 16531 10628 16764 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17793 10659 17851 10665
rect 17793 10625 17805 10659
rect 17839 10656 17851 10659
rect 17954 10656 17960 10668
rect 17839 10628 17960 10656
rect 17839 10625 17851 10628
rect 17793 10619 17851 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18064 10665 18092 10696
rect 20272 10696 21496 10724
rect 20272 10668 20300 10696
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 20254 10616 20260 10668
rect 20312 10616 20318 10668
rect 20530 10665 20536 10668
rect 20524 10656 20536 10665
rect 20491 10628 20536 10656
rect 20524 10619 20536 10628
rect 20530 10616 20536 10619
rect 20588 10616 20594 10668
rect 21468 10600 21496 10696
rect 22112 10696 23796 10724
rect 22112 10665 22140 10696
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22364 10659 22422 10665
rect 22364 10625 22376 10659
rect 22410 10656 22422 10659
rect 22922 10656 22928 10668
rect 22410 10628 22928 10656
rect 22410 10625 22422 10628
rect 22364 10619 22422 10625
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14292 10560 15209 10588
rect 13725 10551 13783 10557
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 15746 10548 15752 10600
rect 15804 10548 15810 10600
rect 15838 10548 15844 10600
rect 15896 10548 15902 10600
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19024 10560 19257 10588
rect 19024 10548 19030 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 15764 10520 15792 10548
rect 16574 10520 16580 10532
rect 15764 10492 16580 10520
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 18984 10520 19012 10548
rect 18064 10492 19012 10520
rect 3234 10452 3240 10464
rect 2746 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 4062 10452 4068 10464
rect 3292 10424 4068 10452
rect 3292 10412 3298 10424
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 6454 10412 6460 10464
rect 6512 10452 6518 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6512 10424 6561 10452
rect 6512 10412 6518 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 10686 10412 10692 10464
rect 10744 10412 10750 10464
rect 10962 10412 10968 10464
rect 11020 10412 11026 10464
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 12526 10452 12532 10464
rect 11379 10424 12532 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 13170 10412 13176 10464
rect 13228 10412 13234 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 18064 10452 18092 10492
rect 14792 10424 18092 10452
rect 14792 10412 14798 10424
rect 18138 10412 18144 10464
rect 18196 10412 18202 10464
rect 19260 10452 19288 10551
rect 19426 10548 19432 10600
rect 19484 10548 19490 10600
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 22112 10588 22140 10619
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 23768 10600 23796 10696
rect 27172 10696 27620 10724
rect 24210 10616 24216 10668
rect 24268 10616 24274 10668
rect 26237 10659 26295 10665
rect 26237 10625 26249 10659
rect 26283 10656 26295 10659
rect 26326 10656 26332 10668
rect 26283 10628 26332 10656
rect 26283 10625 26295 10628
rect 26237 10619 26295 10625
rect 26326 10616 26332 10628
rect 26384 10616 26390 10668
rect 21508 10560 22140 10588
rect 21508 10548 21514 10560
rect 23750 10548 23756 10600
rect 23808 10548 23814 10600
rect 25777 10591 25835 10597
rect 25777 10557 25789 10591
rect 25823 10588 25835 10591
rect 25823 10560 25912 10588
rect 25823 10557 25835 10560
rect 25777 10551 25835 10557
rect 25884 10529 25912 10560
rect 26418 10548 26424 10600
rect 26476 10548 26482 10600
rect 27172 10597 27200 10696
rect 27614 10684 27620 10696
rect 27672 10684 27678 10736
rect 29730 10684 29736 10736
rect 29788 10724 29794 10736
rect 30392 10733 30420 10764
rect 30377 10727 30435 10733
rect 30377 10724 30389 10727
rect 29788 10696 30389 10724
rect 29788 10684 29794 10696
rect 30377 10693 30389 10696
rect 30423 10693 30435 10727
rect 30377 10687 30435 10693
rect 30742 10684 30748 10736
rect 30800 10684 30806 10736
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 27413 10659 27471 10665
rect 27413 10656 27425 10659
rect 27304 10628 27425 10656
rect 27304 10616 27310 10628
rect 27413 10625 27425 10628
rect 27459 10625 27471 10659
rect 27413 10619 27471 10625
rect 27706 10616 27712 10668
rect 27764 10656 27770 10668
rect 28629 10659 28687 10665
rect 28629 10656 28641 10659
rect 27764 10628 28641 10656
rect 27764 10616 27770 10628
rect 28629 10625 28641 10628
rect 28675 10625 28687 10659
rect 28629 10619 28687 10625
rect 27157 10591 27215 10597
rect 27157 10557 27169 10591
rect 27203 10557 27215 10591
rect 30760 10588 30788 10684
rect 32140 10668 32168 10764
rect 33594 10752 33600 10804
rect 33652 10752 33658 10804
rect 34057 10795 34115 10801
rect 34057 10761 34069 10795
rect 34103 10792 34115 10795
rect 34422 10792 34428 10804
rect 34103 10764 34428 10792
rect 34103 10761 34115 10764
rect 34057 10755 34115 10761
rect 34422 10752 34428 10764
rect 34480 10752 34486 10804
rect 35066 10752 35072 10804
rect 35124 10792 35130 10804
rect 35710 10792 35716 10804
rect 35124 10764 35716 10792
rect 35124 10752 35130 10764
rect 35710 10752 35716 10764
rect 35768 10752 35774 10804
rect 35894 10752 35900 10804
rect 35952 10752 35958 10804
rect 36170 10752 36176 10804
rect 36228 10752 36234 10804
rect 36630 10752 36636 10804
rect 36688 10752 36694 10804
rect 39209 10795 39267 10801
rect 39209 10761 39221 10795
rect 39255 10792 39267 10795
rect 39298 10792 39304 10804
rect 39255 10764 39304 10792
rect 39255 10761 39267 10764
rect 39209 10755 39267 10761
rect 39298 10752 39304 10764
rect 39356 10752 39362 10804
rect 40773 10795 40831 10801
rect 40773 10761 40785 10795
rect 40819 10761 40831 10795
rect 40773 10755 40831 10761
rect 32392 10727 32450 10733
rect 32392 10693 32404 10727
rect 32438 10724 32450 10727
rect 33042 10724 33048 10736
rect 32438 10696 33048 10724
rect 32438 10693 32450 10696
rect 32392 10687 32450 10693
rect 33042 10684 33048 10696
rect 33100 10684 33106 10736
rect 34968 10727 35026 10733
rect 34968 10693 34980 10727
rect 35014 10724 35026 10727
rect 35618 10724 35624 10736
rect 35014 10696 35624 10724
rect 35014 10693 35026 10696
rect 34968 10687 35026 10693
rect 35618 10684 35624 10696
rect 35676 10684 35682 10736
rect 35912 10724 35940 10752
rect 36541 10727 36599 10733
rect 36541 10724 36553 10727
rect 35912 10696 36553 10724
rect 36541 10693 36553 10696
rect 36587 10693 36599 10727
rect 37550 10724 37556 10736
rect 36541 10687 36599 10693
rect 37548 10684 37556 10724
rect 37608 10724 37614 10736
rect 39316 10724 39344 10752
rect 37608 10696 39344 10724
rect 37608 10684 37614 10696
rect 30926 10616 30932 10668
rect 30984 10616 30990 10668
rect 32122 10616 32128 10668
rect 32180 10616 32186 10668
rect 33962 10616 33968 10668
rect 34020 10616 34026 10668
rect 34701 10659 34759 10665
rect 34701 10625 34713 10659
rect 34747 10656 34759 10659
rect 34790 10656 34796 10668
rect 34747 10628 34796 10656
rect 34747 10625 34759 10628
rect 34701 10619 34759 10625
rect 34790 10616 34796 10628
rect 34848 10616 34854 10668
rect 31297 10591 31355 10597
rect 31297 10588 31309 10591
rect 30760 10560 31309 10588
rect 27157 10551 27215 10557
rect 31297 10557 31309 10560
rect 31343 10557 31355 10591
rect 31297 10551 31355 10557
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 23032 10492 24041 10520
rect 21266 10452 21272 10464
rect 19260 10424 21272 10452
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 23032 10452 23060 10492
rect 24029 10489 24041 10492
rect 24075 10489 24087 10523
rect 24029 10483 24087 10489
rect 25869 10523 25927 10529
rect 25869 10489 25881 10523
rect 25915 10489 25927 10523
rect 25869 10483 25927 10489
rect 27172 10464 27200 10551
rect 33778 10548 33784 10600
rect 33836 10548 33842 10600
rect 34149 10591 34207 10597
rect 34149 10557 34161 10591
rect 34195 10557 34207 10591
rect 34149 10551 34207 10557
rect 33505 10523 33563 10529
rect 33505 10489 33517 10523
rect 33551 10520 33563 10523
rect 33796 10520 33824 10548
rect 33551 10492 33824 10520
rect 33551 10489 33563 10492
rect 33505 10483 33563 10489
rect 34164 10464 34192 10551
rect 36354 10548 36360 10600
rect 36412 10548 36418 10600
rect 36538 10548 36544 10600
rect 36596 10588 36602 10600
rect 36725 10591 36783 10597
rect 36725 10588 36737 10591
rect 36596 10560 36737 10588
rect 36596 10548 36602 10560
rect 36725 10557 36737 10560
rect 36771 10557 36783 10591
rect 36725 10551 36783 10557
rect 37461 10591 37519 10597
rect 37461 10557 37473 10591
rect 37507 10588 37519 10591
rect 37548 10588 37576 10684
rect 37728 10659 37786 10665
rect 37728 10625 37740 10659
rect 37774 10656 37786 10659
rect 38562 10656 38568 10668
rect 37774 10628 38568 10656
rect 37774 10625 37786 10628
rect 37728 10619 37786 10625
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 39316 10656 39344 10696
rect 39660 10727 39718 10733
rect 39660 10693 39672 10727
rect 39706 10724 39718 10727
rect 40034 10724 40040 10736
rect 39706 10696 40040 10724
rect 39706 10693 39718 10696
rect 39660 10687 39718 10693
rect 40034 10684 40040 10696
rect 40092 10684 40098 10736
rect 40788 10724 40816 10755
rect 40862 10752 40868 10804
rect 40920 10752 40926 10804
rect 41322 10752 41328 10804
rect 41380 10752 41386 10804
rect 41969 10795 42027 10801
rect 41969 10761 41981 10795
rect 42015 10792 42027 10795
rect 42610 10792 42616 10804
rect 42015 10764 42616 10792
rect 42015 10761 42027 10764
rect 41969 10755 42027 10761
rect 41340 10724 41368 10752
rect 40788 10696 41368 10724
rect 39393 10659 39451 10665
rect 39393 10656 39405 10659
rect 39316 10628 39405 10656
rect 39393 10625 39405 10628
rect 39439 10625 39451 10659
rect 39393 10619 39451 10625
rect 41233 10659 41291 10665
rect 41233 10625 41245 10659
rect 41279 10625 41291 10659
rect 41233 10619 41291 10625
rect 37507 10560 37576 10588
rect 37507 10557 37519 10560
rect 37461 10551 37519 10557
rect 36081 10523 36139 10529
rect 36081 10489 36093 10523
rect 36127 10520 36139 10523
rect 36372 10520 36400 10548
rect 36127 10492 36400 10520
rect 41248 10520 41276 10619
rect 41322 10548 41328 10600
rect 41380 10548 41386 10600
rect 41509 10591 41567 10597
rect 41509 10557 41521 10591
rect 41555 10588 41567 10591
rect 41984 10588 42012 10755
rect 42610 10752 42616 10764
rect 42668 10752 42674 10804
rect 43898 10752 43904 10804
rect 43956 10752 43962 10804
rect 45922 10752 45928 10804
rect 45980 10792 45986 10804
rect 46017 10795 46075 10801
rect 46017 10792 46029 10795
rect 45980 10764 46029 10792
rect 45980 10752 45986 10764
rect 46017 10761 46029 10764
rect 46063 10761 46075 10795
rect 46017 10755 46075 10761
rect 47762 10752 47768 10804
rect 47820 10792 47826 10804
rect 47857 10795 47915 10801
rect 47857 10792 47869 10795
rect 47820 10764 47869 10792
rect 47820 10752 47826 10764
rect 47857 10761 47869 10764
rect 47903 10761 47915 10795
rect 47857 10755 47915 10761
rect 47949 10795 48007 10801
rect 47949 10761 47961 10795
rect 47995 10792 48007 10795
rect 48682 10792 48688 10804
rect 47995 10764 48688 10792
rect 47995 10761 48007 10764
rect 47949 10755 48007 10761
rect 42696 10727 42754 10733
rect 42696 10693 42708 10727
rect 42742 10724 42754 10727
rect 43530 10724 43536 10736
rect 42742 10696 43536 10724
rect 42742 10693 42754 10696
rect 42696 10687 42754 10693
rect 43530 10684 43536 10696
rect 43588 10684 43594 10736
rect 44904 10727 44962 10733
rect 44904 10693 44916 10727
rect 44950 10724 44962 10727
rect 45094 10724 45100 10736
rect 44950 10696 45100 10724
rect 44950 10693 44962 10696
rect 44904 10687 44962 10693
rect 45094 10684 45100 10696
rect 45152 10684 45158 10736
rect 46569 10727 46627 10733
rect 46569 10693 46581 10727
rect 46615 10724 46627 10727
rect 47394 10724 47400 10736
rect 46615 10696 47400 10724
rect 46615 10693 46627 10696
rect 46569 10687 46627 10693
rect 47394 10684 47400 10696
rect 47452 10684 47458 10736
rect 42058 10616 42064 10668
rect 42116 10656 42122 10668
rect 42429 10659 42487 10665
rect 42429 10656 42441 10659
rect 42116 10628 42441 10656
rect 42116 10616 42122 10628
rect 42429 10625 42441 10628
rect 42475 10625 42487 10659
rect 42429 10619 42487 10625
rect 44634 10616 44640 10668
rect 44692 10616 44698 10668
rect 45646 10616 45652 10668
rect 45704 10656 45710 10668
rect 46477 10659 46535 10665
rect 46477 10656 46489 10659
rect 45704 10628 46489 10656
rect 45704 10616 45710 10628
rect 46477 10625 46489 10628
rect 46523 10656 46535 10659
rect 47964 10656 47992 10755
rect 48682 10752 48688 10764
rect 48740 10752 48746 10804
rect 49697 10795 49755 10801
rect 49697 10761 49709 10795
rect 49743 10792 49755 10795
rect 49786 10792 49792 10804
rect 49743 10764 49792 10792
rect 49743 10761 49755 10764
rect 49697 10755 49755 10761
rect 49786 10752 49792 10764
rect 49844 10752 49850 10804
rect 51994 10792 52000 10804
rect 51046 10764 52000 10792
rect 48130 10684 48136 10736
rect 48188 10684 48194 10736
rect 48590 10684 48596 10736
rect 48648 10724 48654 10736
rect 51046 10724 51074 10764
rect 51994 10752 52000 10764
rect 52052 10792 52058 10804
rect 53374 10792 53380 10804
rect 52052 10764 53380 10792
rect 52052 10752 52058 10764
rect 53374 10752 53380 10764
rect 53432 10752 53438 10804
rect 55033 10795 55091 10801
rect 55033 10761 55045 10795
rect 55079 10792 55091 10795
rect 55858 10792 55864 10804
rect 55079 10764 55864 10792
rect 55079 10761 55091 10764
rect 55033 10755 55091 10761
rect 55858 10752 55864 10764
rect 55916 10752 55922 10804
rect 56502 10752 56508 10804
rect 56560 10752 56566 10804
rect 56965 10795 57023 10801
rect 56965 10761 56977 10795
rect 57011 10792 57023 10795
rect 57054 10792 57060 10804
rect 57011 10764 57060 10792
rect 57011 10761 57023 10764
rect 56965 10755 57023 10761
rect 57054 10752 57060 10764
rect 57112 10752 57118 10804
rect 57330 10752 57336 10804
rect 57388 10752 57394 10804
rect 48648 10696 51074 10724
rect 51436 10727 51494 10733
rect 48648 10684 48654 10696
rect 51436 10693 51448 10727
rect 51482 10724 51494 10727
rect 52730 10724 52736 10736
rect 51482 10696 52736 10724
rect 51482 10693 51494 10696
rect 51436 10687 51494 10693
rect 52730 10684 52736 10696
rect 52788 10684 52794 10736
rect 54573 10727 54631 10733
rect 54573 10693 54585 10727
rect 54619 10724 54631 10727
rect 55769 10727 55827 10733
rect 55769 10724 55781 10727
rect 54619 10696 55781 10724
rect 54619 10693 54631 10696
rect 54573 10687 54631 10693
rect 55769 10693 55781 10696
rect 55815 10724 55827 10727
rect 56520 10724 56548 10752
rect 55815 10696 56548 10724
rect 57072 10724 57100 10752
rect 57885 10727 57943 10733
rect 57885 10724 57897 10727
rect 57072 10696 57897 10724
rect 55815 10693 55827 10696
rect 55769 10687 55827 10693
rect 57885 10693 57897 10696
rect 57931 10693 57943 10727
rect 57885 10687 57943 10693
rect 46523 10628 47992 10656
rect 46523 10625 46535 10628
rect 46477 10619 46535 10625
rect 41555 10560 42012 10588
rect 41555 10557 41567 10560
rect 41509 10551 41567 10557
rect 44450 10548 44456 10600
rect 44508 10548 44514 10600
rect 46661 10591 46719 10597
rect 46661 10588 46673 10591
rect 46032 10560 46673 10588
rect 41966 10520 41972 10532
rect 41248 10492 41972 10520
rect 36127 10489 36139 10492
rect 36081 10483 36139 10489
rect 41966 10480 41972 10492
rect 42024 10480 42030 10532
rect 43732 10492 44680 10520
rect 22152 10424 23060 10452
rect 23477 10455 23535 10461
rect 22152 10412 22158 10424
rect 23477 10421 23489 10455
rect 23523 10452 23535 10455
rect 23842 10452 23848 10464
rect 23523 10424 23848 10452
rect 23523 10421 23535 10424
rect 23477 10415 23535 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 25130 10412 25136 10464
rect 25188 10412 25194 10464
rect 27154 10412 27160 10464
rect 27212 10412 27218 10464
rect 28534 10412 28540 10464
rect 28592 10412 28598 10464
rect 29546 10412 29552 10464
rect 29604 10452 29610 10464
rect 34146 10452 34152 10464
rect 29604 10424 34152 10452
rect 29604 10412 29610 10424
rect 34146 10412 34152 10424
rect 34204 10412 34210 10464
rect 38838 10412 38844 10464
rect 38896 10412 38902 10464
rect 40770 10412 40776 10464
rect 40828 10452 40834 10464
rect 42702 10452 42708 10464
rect 40828 10424 42708 10452
rect 40828 10412 40834 10424
rect 42702 10412 42708 10424
rect 42760 10452 42766 10464
rect 43732 10452 43760 10492
rect 42760 10424 43760 10452
rect 42760 10412 42766 10424
rect 43806 10412 43812 10464
rect 43864 10412 43870 10464
rect 44652 10452 44680 10492
rect 46032 10452 46060 10560
rect 46661 10557 46673 10560
rect 46707 10588 46719 10591
rect 47121 10591 47179 10597
rect 47121 10588 47133 10591
rect 46707 10560 47133 10588
rect 46707 10557 46719 10560
rect 46661 10551 46719 10557
rect 47121 10557 47133 10560
rect 47167 10557 47179 10591
rect 47121 10551 47179 10557
rect 47765 10591 47823 10597
rect 47765 10557 47777 10591
rect 47811 10588 47823 10591
rect 47946 10588 47952 10600
rect 47811 10560 47952 10588
rect 47811 10557 47823 10560
rect 47765 10551 47823 10557
rect 44652 10424 46060 10452
rect 46106 10412 46112 10464
rect 46164 10412 46170 10464
rect 47136 10452 47164 10551
rect 47946 10548 47952 10560
rect 48004 10548 48010 10600
rect 48148 10588 48176 10684
rect 48222 10616 48228 10668
rect 48280 10656 48286 10668
rect 49421 10659 49479 10665
rect 49421 10656 49433 10659
rect 48280 10628 49433 10656
rect 48280 10616 48286 10628
rect 49421 10625 49433 10628
rect 49467 10656 49479 10659
rect 49467 10628 49832 10656
rect 49467 10625 49479 10628
rect 49421 10619 49479 10625
rect 48961 10591 49019 10597
rect 48961 10588 48973 10591
rect 48148 10560 48973 10588
rect 48961 10557 48973 10560
rect 49007 10557 49019 10591
rect 48961 10551 49019 10557
rect 49694 10548 49700 10600
rect 49752 10548 49758 10600
rect 49804 10588 49832 10628
rect 49878 10616 49884 10668
rect 49936 10616 49942 10668
rect 50522 10656 50528 10668
rect 49988 10628 50528 10656
rect 49988 10588 50016 10628
rect 50522 10616 50528 10628
rect 50580 10616 50586 10668
rect 51166 10616 51172 10668
rect 51224 10616 51230 10668
rect 53098 10616 53104 10668
rect 53156 10656 53162 10668
rect 53561 10659 53619 10665
rect 53561 10656 53573 10659
rect 53156 10628 53573 10656
rect 53156 10616 53162 10628
rect 53561 10625 53573 10628
rect 53607 10625 53619 10659
rect 53561 10619 53619 10625
rect 54036 10628 54248 10656
rect 49804 10560 50016 10588
rect 50246 10548 50252 10600
rect 50304 10548 50310 10600
rect 52730 10548 52736 10600
rect 52788 10588 52794 10600
rect 53193 10591 53251 10597
rect 53193 10588 53205 10591
rect 52788 10560 53205 10588
rect 52788 10548 52794 10560
rect 53193 10557 53205 10560
rect 53239 10557 53251 10591
rect 53193 10551 53251 10557
rect 53374 10548 53380 10600
rect 53432 10588 53438 10600
rect 54036 10588 54064 10628
rect 53432 10560 54064 10588
rect 54113 10591 54171 10597
rect 53432 10548 53438 10560
rect 54113 10557 54125 10591
rect 54159 10557 54171 10591
rect 54113 10551 54171 10557
rect 48317 10523 48375 10529
rect 48317 10489 48329 10523
rect 48363 10520 48375 10523
rect 49712 10520 49740 10548
rect 48363 10492 49740 10520
rect 52549 10523 52607 10529
rect 48363 10489 48375 10492
rect 48317 10483 48375 10489
rect 52549 10489 52561 10523
rect 52595 10520 52607 10523
rect 54128 10520 54156 10551
rect 52595 10492 54156 10520
rect 54220 10520 54248 10628
rect 54662 10616 54668 10668
rect 54720 10656 54726 10668
rect 56873 10659 56931 10665
rect 56873 10656 56885 10659
rect 54720 10628 56885 10656
rect 54720 10616 54726 10628
rect 56873 10625 56885 10628
rect 56919 10656 56931 10659
rect 56962 10656 56968 10668
rect 56919 10628 56968 10656
rect 56919 10625 56931 10628
rect 56873 10619 56931 10625
rect 56962 10616 56968 10628
rect 57020 10616 57026 10668
rect 58434 10616 58440 10668
rect 58492 10616 58498 10668
rect 54294 10548 54300 10600
rect 54352 10588 54358 10600
rect 54481 10591 54539 10597
rect 54481 10588 54493 10591
rect 54352 10560 54493 10588
rect 54352 10548 54358 10560
rect 54481 10557 54493 10560
rect 54527 10588 54539 10591
rect 55030 10588 55036 10600
rect 54527 10560 55036 10588
rect 54527 10557 54539 10560
rect 54481 10551 54539 10557
rect 55030 10548 55036 10560
rect 55088 10548 55094 10600
rect 55122 10548 55128 10600
rect 55180 10588 55186 10600
rect 55217 10591 55275 10597
rect 55217 10588 55229 10591
rect 55180 10560 55229 10588
rect 55180 10548 55186 10560
rect 55217 10557 55229 10560
rect 55263 10557 55275 10591
rect 55217 10551 55275 10557
rect 56505 10591 56563 10597
rect 56505 10557 56517 10591
rect 56551 10588 56563 10591
rect 56778 10588 56784 10600
rect 56551 10560 56784 10588
rect 56551 10557 56563 10560
rect 56505 10551 56563 10557
rect 56520 10520 56548 10551
rect 56778 10548 56784 10560
rect 56836 10548 56842 10600
rect 54220 10492 56548 10520
rect 52595 10489 52607 10492
rect 52549 10483 52607 10489
rect 48038 10452 48044 10464
rect 47136 10424 48044 10452
rect 48038 10412 48044 10424
rect 48096 10412 48102 10464
rect 50798 10412 50804 10464
rect 50856 10412 50862 10464
rect 52733 10455 52791 10461
rect 52733 10421 52745 10455
rect 52779 10452 52791 10455
rect 53282 10452 53288 10464
rect 52779 10424 53288 10452
rect 52779 10421 52791 10424
rect 52733 10415 52791 10421
rect 53282 10412 53288 10424
rect 53340 10412 53346 10464
rect 1104 10362 58880 10384
rect 1104 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 22616 10362
rect 22668 10310 22680 10362
rect 22732 10310 22744 10362
rect 22796 10310 22808 10362
rect 22860 10310 22872 10362
rect 22924 10310 37060 10362
rect 37112 10310 37124 10362
rect 37176 10310 37188 10362
rect 37240 10310 37252 10362
rect 37304 10310 37316 10362
rect 37368 10310 51504 10362
rect 51556 10310 51568 10362
rect 51620 10310 51632 10362
rect 51684 10310 51696 10362
rect 51748 10310 51760 10362
rect 51812 10310 58880 10362
rect 1104 10288 58880 10310
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3326 10248 3332 10260
rect 3191 10220 3332 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3418 10208 3424 10260
rect 3476 10208 3482 10260
rect 4522 10208 4528 10260
rect 4580 10208 4586 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8076 10220 8769 10248
rect 8076 10208 8082 10220
rect 8757 10217 8769 10220
rect 8803 10248 8815 10251
rect 9858 10248 9864 10260
rect 8803 10220 9864 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 10100 10220 10149 10248
rect 10100 10208 10106 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 10284 10220 10425 10248
rect 10284 10208 10290 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 10686 10208 10692 10260
rect 10744 10208 10750 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 12124 10220 12541 10248
rect 12124 10208 12130 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 12529 10211 12587 10217
rect 13170 10208 13176 10260
rect 13228 10208 13234 10260
rect 15473 10251 15531 10257
rect 15473 10217 15485 10251
rect 15519 10248 15531 10251
rect 15838 10248 15844 10260
rect 15519 10220 15844 10248
rect 15519 10217 15531 10220
rect 15473 10211 15531 10217
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 17862 10248 17868 10260
rect 16132 10220 17868 10248
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 5353 10183 5411 10189
rect 5353 10180 5365 10183
rect 3108 10152 3464 10180
rect 3108 10140 3114 10152
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3436 10112 3464 10152
rect 4080 10152 5365 10180
rect 4080 10112 4108 10152
rect 5353 10149 5365 10152
rect 5399 10149 5411 10183
rect 6362 10180 6368 10192
rect 5353 10143 5411 10149
rect 5828 10152 6368 10180
rect 3283 10084 3372 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3050 9936 3056 9988
rect 3108 9936 3114 9988
rect 3344 9920 3372 10084
rect 3436 10084 4108 10112
rect 3436 10053 3464 10084
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3786 10004 3792 10056
rect 3844 10004 3850 10056
rect 3988 10053 4016 10084
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4264 10044 4292 10072
rect 5828 10053 5856 10152
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 7006 10140 7012 10192
rect 7064 10140 7070 10192
rect 8938 10140 8944 10192
rect 8996 10140 9002 10192
rect 9398 10140 9404 10192
rect 9456 10140 9462 10192
rect 6730 10112 6736 10124
rect 5920 10084 6736 10112
rect 5920 10053 5948 10084
rect 6288 10053 6316 10084
rect 6730 10072 6736 10084
rect 6788 10112 6794 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6788 10084 7113 10112
rect 6788 10072 6794 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 9416 10112 9444 10140
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9416 10084 9505 10112
rect 7101 10075 7159 10081
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10704 10112 10732 10208
rect 10965 10115 11023 10121
rect 10965 10112 10977 10115
rect 10008 10084 10456 10112
rect 10704 10084 10977 10112
rect 10008 10072 10014 10084
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 4264 10016 4353 10044
rect 4341 10013 4353 10016
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5491 10016 5549 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5812 10047 5870 10053
rect 5812 10013 5824 10047
rect 5858 10013 5870 10047
rect 5812 10007 5870 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 6272 10047 6330 10053
rect 6272 10044 6284 10047
rect 6251 10016 6284 10044
rect 5905 10007 5963 10013
rect 6272 10013 6284 10016
rect 6318 10013 6330 10047
rect 6272 10007 6330 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 3804 9976 3832 10004
rect 5276 9976 5304 10007
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 3804 9948 6009 9976
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6380 9920 6408 10007
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6880 10047 6938 10053
rect 6880 10044 6892 10047
rect 6512 10016 6892 10044
rect 6512 10004 6518 10016
rect 6880 10013 6892 10016
rect 6926 10013 6938 10047
rect 6880 10007 6938 10013
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 10428 10044 10456 10084
rect 10965 10081 10977 10084
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11882 10072 11888 10124
rect 11940 10072 11946 10124
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 13188 10121 13216 10208
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 16022 10180 16028 10192
rect 15344 10152 16028 10180
rect 15344 10140 15350 10152
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13814 10072 13820 10124
rect 13872 10072 13878 10124
rect 16132 10112 16160 10220
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18509 10251 18567 10257
rect 18509 10217 18521 10251
rect 18555 10248 18567 10251
rect 18690 10248 18696 10260
rect 18555 10220 18696 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 21450 10208 21456 10260
rect 21508 10208 21514 10260
rect 22462 10248 22468 10260
rect 21836 10220 22468 10248
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16132 10084 16497 10112
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 16758 10072 16764 10124
rect 16816 10072 16822 10124
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 17000 10084 17049 10112
rect 17000 10072 17006 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 17184 10084 17632 10112
rect 17184 10072 17190 10084
rect 10870 10044 10876 10056
rect 10428 10016 10876 10044
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11756 10016 11805 10044
rect 11756 10004 11762 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11900 10044 11928 10072
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 11900 10016 13277 10044
rect 11793 10007 11851 10013
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 6546 9936 6552 9988
rect 6604 9976 6610 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6604 9948 6745 9976
rect 6604 9936 6610 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 7469 9979 7527 9985
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 12250 9976 12256 9988
rect 7515 9948 12256 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 14108 9976 14136 10007
rect 16574 10004 16580 10056
rect 16632 10053 16638 10056
rect 16632 10047 16681 10053
rect 16632 10013 16635 10047
rect 16669 10013 16681 10047
rect 16632 10007 16681 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10013 17555 10047
rect 17604 10044 17632 10084
rect 17678 10072 17684 10124
rect 17736 10072 17742 10124
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10112 18015 10115
rect 18414 10112 18420 10124
rect 18003 10084 18420 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 21836 10112 21864 10220
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 29825 10251 29883 10257
rect 29825 10248 29837 10251
rect 26476 10220 29837 10248
rect 26476 10208 26482 10220
rect 29825 10217 29837 10220
rect 29871 10248 29883 10251
rect 30926 10248 30932 10260
rect 29871 10220 30932 10248
rect 29871 10217 29883 10220
rect 29825 10211 29883 10217
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 31389 10251 31447 10257
rect 31389 10217 31401 10251
rect 31435 10248 31447 10251
rect 31570 10248 31576 10260
rect 31435 10220 31576 10248
rect 31435 10217 31447 10220
rect 31389 10211 31447 10217
rect 31570 10208 31576 10220
rect 31628 10208 31634 10260
rect 34146 10208 34152 10260
rect 34204 10248 34210 10260
rect 34425 10251 34483 10257
rect 34425 10248 34437 10251
rect 34204 10220 34437 10248
rect 34204 10208 34210 10220
rect 34425 10217 34437 10220
rect 34471 10217 34483 10251
rect 34425 10211 34483 10217
rect 36538 10208 36544 10260
rect 36596 10248 36602 10260
rect 36596 10220 38608 10248
rect 36596 10208 36602 10220
rect 23566 10180 23572 10192
rect 23124 10152 23572 10180
rect 23124 10124 23152 10152
rect 23566 10140 23572 10152
rect 23624 10140 23630 10192
rect 24213 10183 24271 10189
rect 24213 10149 24225 10183
rect 24259 10180 24271 10183
rect 24259 10152 24992 10180
rect 24259 10149 24271 10152
rect 24213 10143 24271 10149
rect 22465 10115 22523 10121
rect 21836 10084 22232 10112
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 17604 10016 18061 10044
rect 17497 10007 17555 10013
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 20254 10044 20260 10056
rect 19475 10016 20260 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 16632 10004 16638 10007
rect 13832 9948 14136 9976
rect 14360 9979 14418 9985
rect 13832 9920 13860 9948
rect 14360 9945 14372 9979
rect 14406 9976 14418 9979
rect 14550 9976 14556 9988
rect 14406 9948 14556 9976
rect 14406 9945 14418 9948
rect 14360 9939 14418 9945
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 17512 9976 17540 10007
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 22204 10053 22232 10084
rect 22465 10081 22477 10115
rect 22511 10112 22523 10115
rect 22646 10112 22652 10124
rect 22511 10084 22652 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 23106 10112 23112 10124
rect 22787 10084 23112 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23256 10084 23520 10112
rect 23256 10072 23262 10084
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22278 10004 22284 10056
rect 22336 10053 22342 10056
rect 22336 10047 22385 10053
rect 22336 10013 22339 10047
rect 22373 10013 22385 10047
rect 22336 10007 22385 10013
rect 22336 10004 22342 10007
rect 23382 10004 23388 10056
rect 23440 10004 23446 10056
rect 23492 10044 23520 10084
rect 23658 10072 23664 10124
rect 23716 10072 23722 10124
rect 24964 10121 24992 10152
rect 32674 10140 32680 10192
rect 32732 10140 32738 10192
rect 33612 10152 34376 10180
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10081 25007 10115
rect 27154 10112 27160 10124
rect 24949 10075 25007 10081
rect 26252 10084 27160 10112
rect 23845 10047 23903 10053
rect 23845 10044 23857 10047
rect 23492 10016 23857 10044
rect 23845 10013 23857 10016
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 25096 10016 25237 10044
rect 25096 10004 25102 10016
rect 25225 10013 25237 10016
rect 25271 10044 25283 10047
rect 25958 10044 25964 10056
rect 25271 10016 25964 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 25958 10004 25964 10016
rect 26016 10044 26022 10056
rect 26252 10044 26280 10084
rect 27154 10072 27160 10084
rect 27212 10072 27218 10124
rect 27801 10115 27859 10121
rect 27801 10081 27813 10115
rect 27847 10112 27859 10115
rect 27982 10112 27988 10124
rect 27847 10084 27988 10112
rect 27847 10081 27859 10084
rect 27801 10075 27859 10081
rect 27982 10072 27988 10084
rect 28040 10072 28046 10124
rect 28077 10115 28135 10121
rect 28077 10081 28089 10115
rect 28123 10112 28135 10115
rect 28166 10112 28172 10124
rect 28123 10084 28172 10112
rect 28123 10081 28135 10084
rect 28077 10075 28135 10081
rect 28166 10072 28172 10084
rect 28224 10072 28230 10124
rect 28537 10115 28595 10121
rect 28537 10081 28549 10115
rect 28583 10112 28595 10115
rect 28994 10112 29000 10124
rect 28583 10084 29000 10112
rect 28583 10081 28595 10084
rect 28537 10075 28595 10081
rect 28994 10072 29000 10084
rect 29052 10072 29058 10124
rect 29365 10115 29423 10121
rect 29365 10081 29377 10115
rect 29411 10112 29423 10115
rect 29730 10112 29736 10124
rect 29411 10084 29736 10112
rect 29411 10081 29423 10084
rect 29365 10075 29423 10081
rect 29730 10072 29736 10084
rect 29788 10112 29794 10124
rect 30009 10115 30067 10121
rect 30009 10112 30021 10115
rect 29788 10084 30021 10112
rect 29788 10072 29794 10084
rect 30009 10081 30021 10084
rect 30055 10081 30067 10115
rect 30009 10075 30067 10081
rect 31938 10072 31944 10124
rect 31996 10112 32002 10124
rect 32263 10115 32321 10121
rect 32263 10112 32275 10115
rect 31996 10084 32275 10112
rect 31996 10072 32002 10084
rect 32263 10081 32275 10084
rect 32309 10081 32321 10115
rect 32263 10075 32321 10081
rect 32398 10072 32404 10124
rect 32456 10072 32462 10124
rect 33612 10121 33640 10152
rect 34348 10124 34376 10152
rect 37918 10140 37924 10192
rect 37976 10180 37982 10192
rect 37976 10152 38516 10180
rect 37976 10140 37982 10152
rect 33597 10115 33655 10121
rect 33597 10081 33609 10115
rect 33643 10081 33655 10115
rect 33597 10075 33655 10081
rect 33689 10115 33747 10121
rect 33689 10081 33701 10115
rect 33735 10112 33747 10115
rect 33962 10112 33968 10124
rect 33735 10084 33968 10112
rect 33735 10081 33747 10084
rect 33689 10075 33747 10081
rect 33962 10072 33968 10084
rect 34020 10072 34026 10124
rect 34330 10072 34336 10124
rect 34388 10072 34394 10124
rect 34422 10072 34428 10124
rect 34480 10072 34486 10124
rect 35986 10072 35992 10124
rect 36044 10112 36050 10124
rect 37047 10115 37105 10121
rect 37047 10112 37059 10115
rect 36044 10084 37059 10112
rect 36044 10072 36050 10084
rect 37047 10081 37059 10084
rect 37093 10081 37105 10115
rect 37047 10075 37105 10081
rect 37366 10072 37372 10124
rect 37424 10112 37430 10124
rect 37461 10115 37519 10121
rect 37461 10112 37473 10115
rect 37424 10084 37473 10112
rect 37424 10072 37430 10084
rect 37461 10081 37473 10084
rect 37507 10112 37519 10115
rect 37826 10112 37832 10124
rect 37507 10084 37832 10112
rect 37507 10081 37519 10084
rect 37461 10075 37519 10081
rect 37826 10072 37832 10084
rect 37884 10072 37890 10124
rect 38010 10072 38016 10124
rect 38068 10112 38074 10124
rect 38105 10115 38163 10121
rect 38105 10112 38117 10115
rect 38068 10084 38117 10112
rect 38068 10072 38074 10084
rect 38105 10081 38117 10084
rect 38151 10081 38163 10115
rect 38105 10075 38163 10081
rect 38286 10072 38292 10124
rect 38344 10072 38350 10124
rect 38488 10121 38516 10152
rect 38473 10115 38531 10121
rect 38473 10081 38485 10115
rect 38519 10081 38531 10115
rect 38473 10075 38531 10081
rect 26016 10016 26280 10044
rect 26016 10004 26022 10016
rect 27522 10004 27528 10056
rect 27580 10004 27586 10056
rect 27706 10053 27712 10056
rect 27684 10047 27712 10053
rect 27684 10013 27696 10047
rect 27684 10007 27712 10013
rect 27706 10004 27712 10007
rect 27764 10004 27770 10056
rect 28718 10004 28724 10056
rect 28776 10004 28782 10056
rect 30276 10047 30334 10053
rect 30276 10013 30288 10047
rect 30322 10044 30334 10047
rect 30834 10044 30840 10056
rect 30322 10016 30840 10044
rect 30322 10013 30334 10016
rect 30276 10007 30334 10013
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 32122 10004 32128 10056
rect 32180 10004 32186 10056
rect 33137 10047 33195 10053
rect 33137 10013 33149 10047
rect 33183 10013 33195 10047
rect 33137 10007 33195 10013
rect 33321 10047 33379 10053
rect 33321 10013 33333 10047
rect 33367 10044 33379 10047
rect 34440 10044 34468 10072
rect 33367 10016 34468 10044
rect 34701 10047 34759 10053
rect 33367 10013 33379 10016
rect 33321 10007 33379 10013
rect 34701 10013 34713 10047
rect 34747 10044 34759 10047
rect 34790 10044 34796 10056
rect 34747 10016 34796 10044
rect 34747 10013 34759 10016
rect 34701 10007 34759 10013
rect 19696 9979 19754 9985
rect 17512 9948 18184 9976
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 4154 9908 4160 9920
rect 3384 9880 4160 9908
rect 3384 9868 3390 9880
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 7834 9908 7840 9920
rect 6420 9880 7840 9908
rect 6420 9868 6426 9880
rect 7834 9868 7840 9880
rect 7892 9908 7898 9920
rect 8754 9908 8760 9920
rect 7892 9880 8760 9908
rect 7892 9868 7898 9880
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 11422 9868 11428 9920
rect 11480 9868 11486 9920
rect 13814 9868 13820 9920
rect 13872 9868 13878 9920
rect 15841 9911 15899 9917
rect 15841 9877 15853 9911
rect 15887 9908 15899 9911
rect 17954 9908 17960 9920
rect 15887 9880 17960 9908
rect 15887 9877 15899 9880
rect 15841 9871 15899 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 18156 9917 18184 9948
rect 19696 9945 19708 9979
rect 19742 9976 19754 9979
rect 19886 9976 19892 9988
rect 19742 9948 19892 9976
rect 19742 9945 19754 9948
rect 19696 9939 19754 9945
rect 19886 9936 19892 9948
rect 19944 9936 19950 9988
rect 23198 9936 23204 9988
rect 23256 9976 23262 9988
rect 23753 9979 23811 9985
rect 23753 9976 23765 9979
rect 23256 9948 23765 9976
rect 23256 9936 23262 9948
rect 23753 9945 23765 9948
rect 23799 9945 23811 9979
rect 23753 9939 23811 9945
rect 25130 9936 25136 9988
rect 25188 9976 25194 9988
rect 25470 9979 25528 9985
rect 25470 9976 25482 9979
rect 25188 9948 25482 9976
rect 25188 9936 25194 9948
rect 25470 9945 25482 9948
rect 25516 9945 25528 9979
rect 33152 9976 33180 10007
rect 34790 10004 34796 10016
rect 34848 10004 34854 10056
rect 36906 10004 36912 10056
rect 36964 10004 36970 10056
rect 37182 10004 37188 10056
rect 37240 10004 37246 10056
rect 37921 10047 37979 10053
rect 37921 10013 37933 10047
rect 37967 10013 37979 10047
rect 38580 10044 38608 10220
rect 38838 10208 38844 10260
rect 38896 10208 38902 10260
rect 42150 10248 42156 10260
rect 40696 10220 42156 10248
rect 38856 10112 38884 10208
rect 40696 10121 40724 10220
rect 42150 10208 42156 10220
rect 42208 10208 42214 10260
rect 43901 10251 43959 10257
rect 43901 10217 43913 10251
rect 43947 10248 43959 10251
rect 44450 10248 44456 10260
rect 43947 10220 44456 10248
rect 43947 10217 43959 10220
rect 43901 10211 43959 10217
rect 44450 10208 44456 10220
rect 44508 10208 44514 10260
rect 47394 10208 47400 10260
rect 47452 10248 47458 10260
rect 47673 10251 47731 10257
rect 47673 10248 47685 10251
rect 47452 10220 47685 10248
rect 47452 10208 47458 10220
rect 47673 10217 47685 10220
rect 47719 10217 47731 10251
rect 47673 10211 47731 10217
rect 47946 10208 47952 10260
rect 48004 10208 48010 10260
rect 48038 10208 48044 10260
rect 48096 10248 48102 10260
rect 49145 10251 49203 10257
rect 49145 10248 49157 10251
rect 48096 10220 49157 10248
rect 48096 10208 48102 10220
rect 49145 10217 49157 10220
rect 49191 10217 49203 10251
rect 49145 10211 49203 10217
rect 46661 10183 46719 10189
rect 46661 10149 46673 10183
rect 46707 10149 46719 10183
rect 46661 10143 46719 10149
rect 39577 10115 39635 10121
rect 39577 10112 39589 10115
rect 38856 10084 39589 10112
rect 39577 10081 39589 10084
rect 39623 10081 39635 10115
rect 39577 10075 39635 10081
rect 40681 10115 40739 10121
rect 40681 10081 40693 10115
rect 40727 10081 40739 10115
rect 40681 10075 40739 10081
rect 40770 10072 40776 10124
rect 40828 10072 40834 10124
rect 41966 10072 41972 10124
rect 42024 10121 42030 10124
rect 42024 10115 42073 10121
rect 42024 10081 42027 10115
rect 42061 10081 42073 10115
rect 42024 10075 42073 10081
rect 42024 10072 42030 10075
rect 42150 10072 42156 10124
rect 42208 10072 42214 10124
rect 42426 10072 42432 10124
rect 42484 10072 42490 10124
rect 43254 10072 43260 10124
rect 43312 10072 43318 10124
rect 44174 10072 44180 10124
rect 44232 10112 44238 10124
rect 44545 10115 44603 10121
rect 44545 10112 44557 10115
rect 44232 10084 44557 10112
rect 44232 10072 44238 10084
rect 44545 10081 44557 10084
rect 44591 10081 44603 10115
rect 44545 10075 44603 10081
rect 44634 10072 44640 10124
rect 44692 10112 44698 10124
rect 45094 10112 45100 10124
rect 44692 10084 45100 10112
rect 44692 10072 44698 10084
rect 45094 10072 45100 10084
rect 45152 10112 45158 10124
rect 45281 10115 45339 10121
rect 45281 10112 45293 10115
rect 45152 10084 45293 10112
rect 45152 10072 45158 10084
rect 45281 10081 45293 10084
rect 45327 10081 45339 10115
rect 46676 10112 46704 10143
rect 47029 10115 47087 10121
rect 47029 10112 47041 10115
rect 46676 10084 47041 10112
rect 45281 10075 45339 10081
rect 47029 10081 47041 10084
rect 47075 10081 47087 10115
rect 49160 10112 49188 10211
rect 50246 10208 50252 10260
rect 50304 10208 50310 10260
rect 54205 10251 54263 10257
rect 54205 10248 54217 10251
rect 50816 10220 54217 10248
rect 50816 10121 50844 10220
rect 54205 10217 54217 10220
rect 54251 10248 54263 10251
rect 54294 10248 54300 10260
rect 54251 10220 54300 10248
rect 54251 10217 54263 10220
rect 54205 10211 54263 10217
rect 54294 10208 54300 10220
rect 54352 10208 54358 10260
rect 55398 10208 55404 10260
rect 55456 10248 55462 10260
rect 56318 10248 56324 10260
rect 55456 10220 56324 10248
rect 55456 10208 55462 10220
rect 56318 10208 56324 10220
rect 56376 10208 56382 10260
rect 53098 10140 53104 10192
rect 53156 10140 53162 10192
rect 53285 10183 53343 10189
rect 53285 10149 53297 10183
rect 53331 10180 53343 10183
rect 53374 10180 53380 10192
rect 53331 10152 53380 10180
rect 53331 10149 53343 10152
rect 53285 10143 53343 10149
rect 53374 10140 53380 10152
rect 53432 10140 53438 10192
rect 50801 10115 50859 10121
rect 50801 10112 50813 10115
rect 49160 10084 50813 10112
rect 47029 10075 47087 10081
rect 50801 10081 50813 10084
rect 50847 10081 50859 10115
rect 51997 10115 52055 10121
rect 51997 10112 52009 10115
rect 50801 10075 50859 10081
rect 51046 10084 52009 10112
rect 40037 10047 40095 10053
rect 40037 10044 40049 10047
rect 38580 10016 40049 10044
rect 37921 10007 37979 10013
rect 40037 10013 40049 10016
rect 40083 10044 40095 10047
rect 40788 10044 40816 10072
rect 40083 10016 40816 10044
rect 40083 10013 40095 10016
rect 40037 10007 40095 10013
rect 33594 9976 33600 9988
rect 33152 9948 33600 9976
rect 25470 9939 25528 9945
rect 33594 9936 33600 9948
rect 33652 9976 33658 9988
rect 33781 9979 33839 9985
rect 33781 9976 33793 9979
rect 33652 9948 33793 9976
rect 33652 9936 33658 9948
rect 33781 9945 33793 9948
rect 33827 9945 33839 9979
rect 33781 9939 33839 9945
rect 34968 9979 35026 9985
rect 34968 9945 34980 9979
rect 35014 9976 35026 9979
rect 35250 9976 35256 9988
rect 35014 9948 35256 9976
rect 35014 9945 35026 9948
rect 34968 9939 35026 9945
rect 35250 9936 35256 9948
rect 35308 9936 35314 9988
rect 37936 9976 37964 10007
rect 41874 10004 41880 10056
rect 41932 10004 41938 10056
rect 42889 10047 42947 10053
rect 42889 10013 42901 10047
rect 42935 10013 42947 10047
rect 42889 10007 42947 10013
rect 43073 10047 43131 10053
rect 43073 10013 43085 10047
rect 43119 10044 43131 10047
rect 43346 10044 43352 10056
rect 43119 10016 43352 10044
rect 43119 10013 43131 10016
rect 43073 10007 43131 10013
rect 38565 9979 38623 9985
rect 38565 9976 38577 9979
rect 35360 9948 36400 9976
rect 37936 9948 38577 9976
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18230 9908 18236 9920
rect 18187 9880 18236 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18966 9868 18972 9920
rect 19024 9868 19030 9920
rect 20806 9868 20812 9920
rect 20864 9868 20870 9920
rect 21545 9911 21603 9917
rect 21545 9877 21557 9911
rect 21591 9908 21603 9911
rect 23658 9908 23664 9920
rect 21591 9880 23664 9908
rect 21591 9877 21603 9880
rect 21545 9871 21603 9877
rect 23658 9868 23664 9880
rect 23716 9868 23722 9920
rect 24394 9868 24400 9920
rect 24452 9868 24458 9920
rect 26602 9868 26608 9920
rect 26660 9868 26666 9920
rect 26881 9911 26939 9917
rect 26881 9877 26893 9911
rect 26927 9908 26939 9911
rect 28074 9908 28080 9920
rect 26927 9880 28080 9908
rect 26927 9877 26939 9880
rect 26881 9871 26939 9877
rect 28074 9868 28080 9880
rect 28132 9868 28138 9920
rect 31481 9911 31539 9917
rect 31481 9877 31493 9911
rect 31527 9908 31539 9911
rect 32950 9908 32956 9920
rect 31527 9880 32956 9908
rect 31527 9877 31539 9880
rect 31481 9871 31539 9877
rect 32950 9868 32956 9880
rect 33008 9868 33014 9920
rect 34146 9868 34152 9920
rect 34204 9868 34210 9920
rect 34422 9868 34428 9920
rect 34480 9908 34486 9920
rect 35360 9908 35388 9948
rect 34480 9880 35388 9908
rect 34480 9868 34486 9880
rect 36078 9868 36084 9920
rect 36136 9868 36142 9920
rect 36262 9868 36268 9920
rect 36320 9868 36326 9920
rect 36372 9908 36400 9948
rect 38565 9945 38577 9948
rect 38611 9976 38623 9979
rect 39025 9979 39083 9985
rect 39025 9976 39037 9979
rect 38611 9948 39037 9976
rect 38611 9945 38623 9948
rect 38565 9939 38623 9945
rect 39025 9945 39037 9948
rect 39071 9945 39083 9979
rect 39025 9939 39083 9945
rect 40589 9979 40647 9985
rect 40589 9945 40601 9979
rect 40635 9976 40647 9979
rect 41322 9976 41328 9988
rect 40635 9948 41328 9976
rect 40635 9945 40647 9948
rect 40589 9939 40647 9945
rect 41322 9936 41328 9948
rect 41380 9936 41386 9988
rect 42904 9976 42932 10007
rect 43346 10004 43352 10016
rect 43404 10004 43410 10056
rect 49421 10047 49479 10053
rect 49421 10013 49433 10047
rect 49467 10044 49479 10047
rect 49694 10044 49700 10056
rect 49467 10016 49700 10044
rect 49467 10013 49479 10016
rect 49421 10007 49479 10013
rect 49694 10004 49700 10016
rect 49752 10004 49758 10056
rect 50614 10004 50620 10056
rect 50672 10004 50678 10056
rect 51046 10044 51074 10084
rect 51997 10081 52009 10084
rect 52043 10081 52055 10115
rect 51997 10075 52055 10081
rect 52273 10115 52331 10121
rect 52273 10081 52285 10115
rect 52319 10112 52331 10115
rect 52733 10115 52791 10121
rect 52319 10084 52684 10112
rect 52319 10081 52331 10084
rect 52273 10075 52331 10081
rect 50724 10016 51074 10044
rect 43533 9979 43591 9985
rect 43533 9976 43545 9979
rect 42904 9948 43545 9976
rect 43533 9945 43545 9948
rect 43579 9976 43591 9979
rect 43993 9979 44051 9985
rect 43993 9976 44005 9979
rect 43579 9948 44005 9976
rect 43579 9945 43591 9948
rect 43533 9939 43591 9945
rect 43993 9945 44005 9948
rect 44039 9945 44051 9979
rect 43993 9939 44051 9945
rect 45548 9979 45606 9985
rect 45548 9945 45560 9979
rect 45594 9976 45606 9979
rect 45830 9976 45836 9988
rect 45594 9948 45836 9976
rect 45594 9945 45606 9948
rect 45548 9939 45606 9945
rect 45830 9936 45836 9948
rect 45888 9936 45894 9988
rect 48130 9936 48136 9988
rect 48188 9936 48194 9988
rect 50724 9985 50752 10016
rect 51718 10004 51724 10056
rect 51776 10004 51782 10056
rect 51902 10053 51908 10056
rect 51880 10047 51908 10053
rect 51880 10013 51892 10047
rect 51880 10007 51908 10013
rect 51902 10004 51908 10007
rect 51960 10004 51966 10056
rect 52656 10044 52684 10084
rect 52733 10081 52745 10115
rect 52779 10112 52791 10115
rect 53116 10112 53144 10140
rect 52779 10084 53144 10112
rect 52779 10081 52791 10084
rect 52733 10075 52791 10081
rect 57238 10072 57244 10124
rect 57296 10112 57302 10124
rect 57517 10115 57575 10121
rect 57517 10112 57529 10115
rect 57296 10084 57529 10112
rect 57296 10072 57302 10084
rect 57517 10081 57529 10084
rect 57563 10081 57575 10115
rect 57517 10075 57575 10081
rect 52656 10016 52776 10044
rect 49973 9979 50031 9985
rect 49973 9945 49985 9979
rect 50019 9976 50031 9979
rect 50709 9979 50767 9985
rect 50709 9976 50721 9979
rect 50019 9948 50721 9976
rect 50019 9945 50031 9948
rect 49973 9939 50031 9945
rect 50709 9945 50721 9948
rect 50755 9945 50767 9979
rect 51166 9976 51172 9988
rect 50709 9939 50767 9945
rect 50816 9948 51172 9976
rect 38286 9908 38292 9920
rect 36372 9880 38292 9908
rect 38286 9868 38292 9880
rect 38344 9868 38350 9920
rect 38930 9868 38936 9920
rect 38988 9868 38994 9920
rect 40221 9911 40279 9917
rect 40221 9877 40233 9911
rect 40267 9908 40279 9911
rect 40494 9908 40500 9920
rect 40267 9880 40500 9908
rect 40267 9877 40279 9880
rect 40221 9871 40279 9877
rect 40494 9868 40500 9880
rect 40552 9868 40558 9920
rect 41233 9911 41291 9917
rect 41233 9877 41245 9911
rect 41279 9908 41291 9911
rect 42886 9908 42892 9920
rect 41279 9880 42892 9908
rect 41279 9877 41291 9880
rect 41233 9871 41291 9877
rect 42886 9868 42892 9880
rect 42944 9868 42950 9920
rect 43438 9868 43444 9920
rect 43496 9868 43502 9920
rect 47854 9868 47860 9920
rect 47912 9908 47918 9920
rect 48148 9908 48176 9936
rect 50816 9908 50844 9948
rect 51166 9936 51172 9948
rect 51224 9936 51230 9988
rect 52748 9976 52776 10016
rect 52914 10004 52920 10056
rect 52972 10004 52978 10056
rect 55306 9976 55312 9988
rect 52748 9948 55312 9976
rect 55306 9936 55312 9948
rect 55364 9936 55370 9988
rect 47912 9880 50844 9908
rect 51077 9911 51135 9917
rect 47912 9868 47918 9880
rect 51077 9877 51089 9911
rect 51123 9908 51135 9911
rect 51994 9908 52000 9920
rect 51123 9880 52000 9908
rect 51123 9877 51135 9880
rect 51077 9871 51135 9877
rect 51994 9868 52000 9880
rect 52052 9868 52058 9920
rect 56962 9868 56968 9920
rect 57020 9868 57026 9920
rect 1104 9818 59040 9840
rect 1104 9766 15394 9818
rect 15446 9766 15458 9818
rect 15510 9766 15522 9818
rect 15574 9766 15586 9818
rect 15638 9766 15650 9818
rect 15702 9766 29838 9818
rect 29890 9766 29902 9818
rect 29954 9766 29966 9818
rect 30018 9766 30030 9818
rect 30082 9766 30094 9818
rect 30146 9766 44282 9818
rect 44334 9766 44346 9818
rect 44398 9766 44410 9818
rect 44462 9766 44474 9818
rect 44526 9766 44538 9818
rect 44590 9766 58726 9818
rect 58778 9766 58790 9818
rect 58842 9766 58854 9818
rect 58906 9766 58918 9818
rect 58970 9766 58982 9818
rect 59034 9766 59040 9818
rect 1104 9744 59040 9766
rect 3326 9664 3332 9716
rect 3384 9664 3390 9716
rect 6089 9707 6147 9713
rect 6089 9673 6101 9707
rect 6135 9704 6147 9707
rect 6362 9704 6368 9716
rect 6135 9676 6368 9704
rect 6135 9673 6147 9676
rect 6089 9667 6147 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 11698 9704 11704 9716
rect 10928 9676 11704 9704
rect 10928 9664 10934 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11793 9707 11851 9713
rect 11793 9673 11805 9707
rect 11839 9704 11851 9707
rect 11974 9704 11980 9716
rect 11839 9676 11980 9704
rect 11839 9673 11851 9676
rect 11793 9667 11851 9673
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 13265 9707 13323 9713
rect 13265 9673 13277 9707
rect 13311 9704 13323 9707
rect 13538 9704 13544 9716
rect 13311 9676 13544 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15252 9676 15761 9704
rect 15252 9664 15258 9676
rect 15749 9673 15761 9676
rect 15795 9704 15807 9707
rect 16022 9704 16028 9716
rect 15795 9676 16028 9704
rect 15795 9673 15807 9676
rect 15749 9667 15807 9673
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 16574 9664 16580 9716
rect 16632 9664 16638 9716
rect 22278 9704 22284 9716
rect 22066 9676 22284 9704
rect 7006 9636 7012 9648
rect 6196 9608 7012 9636
rect 6196 9580 6224 9608
rect 7006 9596 7012 9608
rect 7064 9636 7070 9648
rect 7745 9639 7803 9645
rect 7064 9608 7144 9636
rect 7064 9596 7070 9608
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3252 9376 3280 9531
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 6420 9540 6469 9568
rect 6420 9528 6426 9540
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7116 9577 7144 9608
rect 7745 9605 7757 9639
rect 7791 9636 7803 9639
rect 11238 9636 11244 9648
rect 7791 9608 11244 9636
rect 7791 9605 7803 9608
rect 7745 9599 7803 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 11333 9639 11391 9645
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 11606 9636 11612 9648
rect 11379 9608 11612 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 11606 9596 11612 9608
rect 11664 9596 11670 9648
rect 12529 9639 12587 9645
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 13722 9636 13728 9648
rect 12575 9608 13728 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 15657 9639 15715 9645
rect 14016 9608 15608 9636
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7834 9528 7840 9580
rect 7892 9528 7898 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10134 9568 10140 9580
rect 9907 9540 10140 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 11422 9568 11428 9580
rect 10827 9540 11428 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 12713 9571 12771 9577
rect 11808 9540 12434 9568
rect 8018 9460 8024 9512
rect 8076 9460 8082 9512
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 11808 9500 11836 9540
rect 9953 9463 10011 9469
rect 10152 9472 11836 9500
rect 11885 9503 11943 9509
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 9968 9432 9996 9463
rect 10042 9432 10048 9444
rect 7156 9404 9904 9432
rect 9968 9404 10048 9432
rect 7156 9392 7162 9404
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 8754 9324 8760 9376
rect 8812 9324 8818 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 8938 9364 8944 9376
rect 8895 9336 8944 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 9876 9364 9904 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10152 9364 10180 9472
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 12406 9500 12434 9540
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 12894 9568 12900 9580
rect 12759 9540 12900 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 14016 9568 14044 9608
rect 13740 9540 14044 9568
rect 14084 9571 14142 9577
rect 13740 9500 13768 9540
rect 14084 9537 14096 9571
rect 14130 9568 14142 9571
rect 14366 9568 14372 9580
rect 14130 9540 14372 9568
rect 14130 9537 14142 9540
rect 14084 9531 14142 9537
rect 14366 9528 14372 9540
rect 14424 9528 14430 9580
rect 15580 9568 15608 9608
rect 15657 9605 15669 9639
rect 15703 9636 15715 9639
rect 16592 9636 16620 9664
rect 15703 9608 16620 9636
rect 17804 9639 17862 9645
rect 15703 9605 15715 9608
rect 15657 9599 15715 9605
rect 17804 9605 17816 9639
rect 17850 9636 17862 9639
rect 18138 9636 18144 9648
rect 17850 9608 18144 9636
rect 17850 9605 17862 9608
rect 17804 9599 17862 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 19644 9639 19702 9645
rect 19644 9605 19656 9639
rect 19690 9636 19702 9639
rect 19794 9636 19800 9648
rect 19690 9608 19800 9636
rect 19690 9605 19702 9608
rect 19644 9599 19702 9605
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 20441 9639 20499 9645
rect 20441 9605 20453 9639
rect 20487 9636 20499 9639
rect 22066 9636 22094 9676
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 22373 9707 22431 9713
rect 22373 9673 22385 9707
rect 22419 9673 22431 9707
rect 22373 9667 22431 9673
rect 20487 9608 22094 9636
rect 20487 9605 20499 9608
rect 20441 9599 20499 9605
rect 22186 9596 22192 9648
rect 22244 9636 22250 9648
rect 22388 9636 22416 9667
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 24762 9704 24768 9716
rect 22520 9676 24768 9704
rect 22520 9664 22526 9676
rect 22244 9608 22416 9636
rect 22244 9596 22250 9608
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 15580 9540 16313 9568
rect 16301 9537 16313 9540
rect 16347 9568 16359 9571
rect 16942 9568 16948 9580
rect 16347 9540 16948 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 20548 9540 21281 9568
rect 20548 9512 20576 9540
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9568 21419 9571
rect 22002 9568 22008 9580
rect 21407 9540 22008 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 12406 9472 13768 9500
rect 13817 9503 13875 9509
rect 11885 9463 11943 9469
rect 13817 9469 13829 9503
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 10226 9392 10232 9444
rect 10284 9432 10290 9444
rect 11900 9432 11928 9463
rect 10284 9404 11928 9432
rect 10284 9392 10290 9404
rect 13832 9376 13860 9463
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15896 9472 15945 9500
rect 15896 9460 15902 9472
rect 15933 9469 15945 9472
rect 15979 9500 15991 9503
rect 16482 9500 16488 9512
rect 15979 9472 16488 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 19889 9503 19947 9509
rect 18095 9472 18460 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 15197 9435 15255 9441
rect 15197 9401 15209 9435
rect 15243 9432 15255 9435
rect 15470 9432 15476 9444
rect 15243 9404 15476 9432
rect 15243 9401 15255 9404
rect 15197 9395 15255 9401
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 18432 9376 18460 9472
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 19904 9432 19932 9463
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 21284 9500 21312 9531
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9568 22155 9571
rect 22480 9568 22508 9664
rect 23508 9639 23566 9645
rect 23508 9605 23520 9639
rect 23554 9636 23566 9639
rect 24394 9636 24400 9648
rect 23554 9608 24400 9636
rect 23554 9605 23566 9608
rect 23508 9599 23566 9605
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 24504 9636 24532 9676
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 31938 9664 31944 9716
rect 31996 9664 32002 9716
rect 32122 9664 32128 9716
rect 32180 9704 32186 9716
rect 32180 9676 33456 9704
rect 32180 9664 32186 9676
rect 24504 9608 26556 9636
rect 22143 9540 22508 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 21284 9472 21404 9500
rect 21266 9432 21272 9444
rect 19904 9404 21272 9432
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 21376 9432 21404 9472
rect 21542 9460 21548 9512
rect 21600 9460 21606 9512
rect 22186 9432 22192 9444
rect 21376 9404 22192 9432
rect 22186 9392 22192 9404
rect 22244 9392 22250 9444
rect 9876 9336 10180 9364
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 11054 9364 11060 9376
rect 10643 9336 11060 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 13725 9367 13783 9373
rect 13725 9333 13737 9367
rect 13771 9364 13783 9367
rect 13814 9364 13820 9376
rect 13771 9336 13820 9364
rect 13771 9333 13783 9336
rect 13725 9327 13783 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 15286 9324 15292 9376
rect 15344 9324 15350 9376
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15746 9364 15752 9376
rect 15620 9336 15752 9364
rect 15620 9324 15626 9336
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16666 9324 16672 9376
rect 16724 9324 16730 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 18046 9364 18052 9376
rect 17736 9336 18052 9364
rect 17736 9324 17742 9336
rect 18046 9324 18052 9336
rect 18104 9364 18110 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18104 9336 18337 9364
rect 18104 9324 18110 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 18414 9324 18420 9376
rect 18472 9324 18478 9376
rect 18506 9324 18512 9376
rect 18564 9324 18570 9376
rect 20073 9367 20131 9373
rect 20073 9333 20085 9367
rect 20119 9364 20131 9367
rect 20438 9364 20444 9376
rect 20119 9336 20444 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 20901 9367 20959 9373
rect 20901 9333 20913 9367
rect 20947 9364 20959 9367
rect 21174 9364 21180 9376
rect 20947 9336 21180 9364
rect 20947 9333 20959 9336
rect 20901 9327 20959 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21634 9324 21640 9376
rect 21692 9364 21698 9376
rect 22296 9364 22324 9540
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 23900 9540 24501 9568
rect 23900 9528 23906 9540
rect 24489 9537 24501 9540
rect 24535 9537 24547 9571
rect 24489 9531 24547 9537
rect 25038 9528 25044 9580
rect 25096 9528 25102 9580
rect 25308 9571 25366 9577
rect 25308 9537 25320 9571
rect 25354 9568 25366 9571
rect 25590 9568 25596 9580
rect 25354 9540 25596 9568
rect 25354 9537 25366 9540
rect 25308 9531 25366 9537
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 23750 9460 23756 9512
rect 23808 9500 23814 9512
rect 25056 9500 25084 9528
rect 23808 9472 25084 9500
rect 23808 9460 23814 9472
rect 26528 9376 26556 9608
rect 27154 9596 27160 9648
rect 27212 9636 27218 9648
rect 27249 9639 27307 9645
rect 27249 9636 27261 9639
rect 27212 9608 27261 9636
rect 27212 9596 27218 9608
rect 27249 9605 27261 9608
rect 27295 9636 27307 9639
rect 27295 9608 29868 9636
rect 27295 9605 27307 9608
rect 27249 9599 27307 9605
rect 27632 9577 27660 9608
rect 27890 9577 27896 9580
rect 27617 9571 27675 9577
rect 27617 9537 27629 9571
rect 27663 9537 27675 9571
rect 27884 9568 27896 9577
rect 27851 9540 27896 9568
rect 27617 9531 27675 9537
rect 27884 9531 27896 9540
rect 27890 9528 27896 9531
rect 27948 9528 27954 9580
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29840 9577 29868 9608
rect 33428 9580 33456 9676
rect 33594 9664 33600 9716
rect 33652 9704 33658 9716
rect 33689 9707 33747 9713
rect 33689 9704 33701 9707
rect 33652 9676 33701 9704
rect 33652 9664 33658 9676
rect 33689 9673 33701 9676
rect 33735 9673 33747 9707
rect 33689 9667 33747 9673
rect 35250 9664 35256 9716
rect 35308 9664 35314 9716
rect 35986 9664 35992 9716
rect 36044 9704 36050 9716
rect 36633 9707 36691 9713
rect 36633 9704 36645 9707
rect 36044 9676 36645 9704
rect 36044 9664 36050 9676
rect 36633 9673 36645 9676
rect 36679 9673 36691 9707
rect 36633 9667 36691 9673
rect 38010 9664 38016 9716
rect 38068 9704 38074 9716
rect 38473 9707 38531 9713
rect 38473 9704 38485 9707
rect 38068 9676 38485 9704
rect 38068 9664 38074 9676
rect 38473 9673 38485 9676
rect 38519 9673 38531 9707
rect 38473 9667 38531 9673
rect 38562 9664 38568 9716
rect 38620 9664 38626 9716
rect 40954 9704 40960 9716
rect 38672 9676 40960 9704
rect 33502 9596 33508 9648
rect 33560 9636 33566 9648
rect 33781 9639 33839 9645
rect 33781 9636 33793 9639
rect 33560 9608 33793 9636
rect 33560 9596 33566 9608
rect 33781 9605 33793 9608
rect 33827 9605 33839 9639
rect 33781 9599 33839 9605
rect 38286 9596 38292 9648
rect 38344 9636 38350 9648
rect 38672 9636 38700 9676
rect 40954 9664 40960 9676
rect 41012 9704 41018 9716
rect 41012 9676 41276 9704
rect 41012 9664 41018 9676
rect 38344 9608 38700 9636
rect 38344 9596 38350 9608
rect 40218 9596 40224 9648
rect 40276 9596 40282 9648
rect 29089 9571 29147 9577
rect 29089 9568 29101 9571
rect 29052 9540 29101 9568
rect 29052 9528 29058 9540
rect 29089 9537 29101 9540
rect 29135 9537 29147 9571
rect 29089 9531 29147 9537
rect 29825 9571 29883 9577
rect 29825 9537 29837 9571
rect 29871 9537 29883 9571
rect 29825 9531 29883 9537
rect 30092 9571 30150 9577
rect 30092 9537 30104 9571
rect 30138 9568 30150 9571
rect 32125 9571 32183 9577
rect 32125 9568 32137 9571
rect 30138 9540 32137 9568
rect 30138 9537 30150 9540
rect 30092 9531 30150 9537
rect 32125 9537 32137 9540
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 32214 9528 32220 9580
rect 32272 9568 32278 9580
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32272 9540 33057 9568
rect 32272 9528 32278 9540
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 33410 9528 33416 9580
rect 33468 9528 33474 9580
rect 34146 9528 34152 9580
rect 34204 9568 34210 9580
rect 34333 9571 34391 9577
rect 34333 9568 34345 9571
rect 34204 9540 34345 9568
rect 34204 9528 34210 9540
rect 34333 9537 34345 9540
rect 34379 9537 34391 9571
rect 34333 9531 34391 9537
rect 34517 9571 34575 9577
rect 34517 9537 34529 9571
rect 34563 9568 34575 9571
rect 34698 9568 34704 9580
rect 34563 9540 34704 9568
rect 34563 9537 34575 9540
rect 34517 9531 34575 9537
rect 34698 9528 34704 9540
rect 34756 9528 34762 9580
rect 34974 9528 34980 9580
rect 35032 9568 35038 9580
rect 35161 9571 35219 9577
rect 35161 9568 35173 9571
rect 35032 9540 35173 9568
rect 35032 9528 35038 9540
rect 35161 9537 35173 9540
rect 35207 9537 35219 9571
rect 35161 9531 35219 9537
rect 35526 9528 35532 9580
rect 35584 9568 35590 9580
rect 35897 9571 35955 9577
rect 35897 9568 35909 9571
rect 35584 9540 35909 9568
rect 35584 9528 35590 9540
rect 35897 9537 35909 9540
rect 35943 9537 35955 9571
rect 35897 9531 35955 9537
rect 36078 9528 36084 9580
rect 36136 9528 36142 9580
rect 37642 9528 37648 9580
rect 37700 9568 37706 9580
rect 37829 9571 37887 9577
rect 37829 9568 37841 9571
rect 37700 9540 37841 9568
rect 37700 9528 37706 9540
rect 37829 9537 37841 9540
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 38930 9528 38936 9580
rect 38988 9568 38994 9580
rect 39117 9571 39175 9577
rect 39117 9568 39129 9571
rect 38988 9540 39129 9568
rect 38988 9528 38994 9540
rect 39117 9537 39129 9540
rect 39163 9537 39175 9571
rect 39117 9531 39175 9537
rect 40494 9528 40500 9580
rect 40552 9568 40558 9580
rect 40773 9571 40831 9577
rect 40773 9568 40785 9571
rect 40552 9540 40785 9568
rect 40552 9528 40558 9540
rect 40773 9537 40785 9540
rect 40819 9537 40831 9571
rect 41248 9568 41276 9676
rect 41322 9664 41328 9716
rect 41380 9704 41386 9716
rect 42797 9707 42855 9713
rect 42797 9704 42809 9707
rect 41380 9676 42809 9704
rect 41380 9664 41386 9676
rect 42797 9673 42809 9676
rect 42843 9704 42855 9707
rect 43438 9704 43444 9716
rect 42843 9676 43444 9704
rect 42843 9673 42855 9676
rect 42797 9667 42855 9673
rect 43438 9664 43444 9676
rect 43496 9664 43502 9716
rect 45094 9664 45100 9716
rect 45152 9664 45158 9716
rect 45830 9664 45836 9716
rect 45888 9664 45894 9716
rect 49694 9664 49700 9716
rect 49752 9664 49758 9716
rect 50614 9664 50620 9716
rect 50672 9704 50678 9716
rect 54205 9707 54263 9713
rect 50672 9676 51304 9704
rect 50672 9664 50678 9676
rect 41782 9596 41788 9648
rect 41840 9636 41846 9648
rect 42245 9639 42303 9645
rect 42245 9636 42257 9639
rect 41840 9608 42257 9636
rect 41840 9596 41846 9608
rect 42245 9605 42257 9608
rect 42291 9636 42303 9639
rect 42705 9639 42763 9645
rect 42291 9608 42656 9636
rect 42291 9605 42303 9608
rect 42245 9599 42303 9605
rect 41248 9540 42564 9568
rect 40773 9531 40831 9537
rect 29641 9503 29699 9509
rect 29641 9469 29653 9503
rect 29687 9469 29699 9503
rect 31297 9503 31355 9509
rect 31297 9500 31309 9503
rect 29641 9463 29699 9469
rect 31220 9472 31309 9500
rect 28997 9435 29055 9441
rect 28997 9401 29009 9435
rect 29043 9432 29055 9435
rect 29656 9432 29684 9463
rect 31220 9441 31248 9472
rect 31297 9469 31309 9472
rect 31343 9469 31355 9503
rect 31297 9463 31355 9469
rect 32674 9460 32680 9512
rect 32732 9460 32738 9512
rect 42426 9500 42432 9512
rect 41386 9472 42432 9500
rect 29043 9404 29684 9432
rect 31205 9435 31263 9441
rect 29043 9401 29055 9404
rect 28997 9395 29055 9401
rect 31205 9401 31217 9435
rect 31251 9401 31263 9435
rect 31205 9395 31263 9401
rect 37274 9392 37280 9444
rect 37332 9432 37338 9444
rect 37332 9404 37596 9432
rect 37332 9392 37338 9404
rect 21692 9336 22324 9364
rect 21692 9324 21698 9336
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23440 9336 23857 9364
rect 23440 9324 23446 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 26418 9324 26424 9376
rect 26476 9324 26482 9376
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 26697 9367 26755 9373
rect 26697 9364 26709 9367
rect 26568 9336 26709 9364
rect 26568 9324 26574 9336
rect 26697 9333 26709 9336
rect 26743 9364 26755 9367
rect 27522 9364 27528 9376
rect 26743 9336 27528 9364
rect 26743 9333 26755 9336
rect 26697 9327 26755 9333
rect 27522 9324 27528 9336
rect 27580 9324 27586 9376
rect 36722 9324 36728 9376
rect 36780 9364 36786 9376
rect 36909 9367 36967 9373
rect 36909 9364 36921 9367
rect 36780 9336 36921 9364
rect 36780 9324 36786 9336
rect 36909 9333 36921 9336
rect 36955 9364 36967 9367
rect 37366 9364 37372 9376
rect 36955 9336 37372 9364
rect 36955 9333 36967 9336
rect 36909 9327 36967 9333
rect 37366 9324 37372 9336
rect 37424 9324 37430 9376
rect 37568 9373 37596 9404
rect 37553 9367 37611 9373
rect 37553 9333 37565 9367
rect 37599 9364 37611 9367
rect 37642 9364 37648 9376
rect 37599 9336 37648 9364
rect 37599 9333 37611 9336
rect 37553 9327 37611 9333
rect 37642 9324 37648 9336
rect 37700 9324 37706 9376
rect 40126 9324 40132 9376
rect 40184 9364 40190 9376
rect 41141 9367 41199 9373
rect 41141 9364 41153 9367
rect 40184 9336 41153 9364
rect 40184 9324 40190 9336
rect 41141 9333 41153 9336
rect 41187 9364 41199 9367
rect 41386 9364 41414 9472
rect 42426 9460 42432 9472
rect 42484 9460 42490 9512
rect 42536 9432 42564 9540
rect 42628 9509 42656 9608
rect 42705 9605 42717 9639
rect 42751 9636 42763 9639
rect 43346 9636 43352 9648
rect 42751 9608 43352 9636
rect 42751 9605 42763 9608
rect 42705 9599 42763 9605
rect 43346 9596 43352 9608
rect 43404 9596 43410 9648
rect 45112 9636 45140 9664
rect 46753 9639 46811 9645
rect 46753 9636 46765 9639
rect 45112 9608 46765 9636
rect 46753 9605 46765 9608
rect 46799 9605 46811 9639
rect 46753 9599 46811 9605
rect 50798 9596 50804 9648
rect 50856 9645 50862 9648
rect 50856 9636 50868 9645
rect 50856 9608 50901 9636
rect 50856 9599 50868 9608
rect 50856 9596 50862 9599
rect 43806 9528 43812 9580
rect 43864 9568 43870 9580
rect 43901 9571 43959 9577
rect 43901 9568 43913 9571
rect 43864 9540 43913 9568
rect 43864 9528 43870 9540
rect 43901 9537 43913 9540
rect 43947 9537 43959 9571
rect 43901 9531 43959 9537
rect 46106 9528 46112 9580
rect 46164 9568 46170 9580
rect 46385 9571 46443 9577
rect 46385 9568 46397 9571
rect 46164 9540 46397 9568
rect 46164 9528 46170 9540
rect 46385 9537 46397 9540
rect 46431 9537 46443 9571
rect 51276 9568 51304 9676
rect 54205 9673 54217 9707
rect 54251 9704 54263 9707
rect 54662 9704 54668 9716
rect 54251 9676 54668 9704
rect 54251 9673 54263 9676
rect 54205 9667 54263 9673
rect 54662 9664 54668 9676
rect 54720 9664 54726 9716
rect 56873 9707 56931 9713
rect 56873 9673 56885 9707
rect 56919 9704 56931 9707
rect 57054 9704 57060 9716
rect 56919 9676 57060 9704
rect 56919 9673 56931 9676
rect 56873 9667 56931 9673
rect 57054 9664 57060 9676
rect 57112 9664 57118 9716
rect 51537 9639 51595 9645
rect 51537 9605 51549 9639
rect 51583 9636 51595 9639
rect 51902 9636 51908 9648
rect 51583 9608 51908 9636
rect 51583 9605 51595 9608
rect 51537 9599 51595 9605
rect 51902 9596 51908 9608
rect 51960 9636 51966 9648
rect 52733 9639 52791 9645
rect 52733 9636 52745 9639
rect 51960 9608 52745 9636
rect 51960 9596 51966 9608
rect 52733 9605 52745 9608
rect 52779 9605 52791 9639
rect 55582 9636 55588 9648
rect 52733 9599 52791 9605
rect 54036 9608 55588 9636
rect 51276 9540 51396 9568
rect 46385 9531 46443 9537
rect 42613 9503 42671 9509
rect 42613 9469 42625 9503
rect 42659 9500 42671 9503
rect 47946 9500 47952 9512
rect 42659 9472 47952 9500
rect 42659 9469 42671 9472
rect 42613 9463 42671 9469
rect 47946 9460 47952 9472
rect 48004 9460 48010 9512
rect 48130 9460 48136 9512
rect 48188 9460 48194 9512
rect 51074 9460 51080 9512
rect 51132 9460 51138 9512
rect 51258 9460 51264 9512
rect 51316 9460 51322 9512
rect 51368 9500 51396 9540
rect 51718 9528 51724 9580
rect 51776 9568 51782 9580
rect 52273 9571 52331 9577
rect 52273 9568 52285 9571
rect 51776 9540 52285 9568
rect 51776 9528 51782 9540
rect 52273 9537 52285 9540
rect 52319 9568 52331 9571
rect 54036 9568 54064 9608
rect 55582 9596 55588 9608
rect 55640 9596 55646 9648
rect 52319 9540 54064 9568
rect 54297 9571 54355 9577
rect 52319 9537 52331 9540
rect 52273 9531 52331 9537
rect 54297 9537 54309 9571
rect 54343 9568 54355 9571
rect 56134 9568 56140 9580
rect 54343 9540 56140 9568
rect 54343 9537 54355 9540
rect 54297 9531 54355 9537
rect 56134 9528 56140 9540
rect 56192 9528 56198 9580
rect 56336 9540 57100 9568
rect 56336 9512 56364 9540
rect 51445 9503 51503 9509
rect 51445 9500 51457 9503
rect 51368 9472 51457 9500
rect 51445 9469 51457 9472
rect 51491 9500 51503 9503
rect 52730 9500 52736 9512
rect 51491 9472 52736 9500
rect 51491 9469 51503 9472
rect 51445 9463 51503 9469
rect 52730 9460 52736 9472
rect 52788 9460 52794 9512
rect 53282 9460 53288 9512
rect 53340 9460 53346 9512
rect 54021 9503 54079 9509
rect 54021 9500 54033 9503
rect 53852 9472 54033 9500
rect 43165 9435 43223 9441
rect 42536 9404 42840 9432
rect 41187 9336 41414 9364
rect 41187 9333 41199 9336
rect 41141 9327 41199 9333
rect 41598 9324 41604 9376
rect 41656 9324 41662 9376
rect 42812 9364 42840 9404
rect 43165 9401 43177 9435
rect 43211 9432 43223 9435
rect 44082 9432 44088 9444
rect 43211 9404 44088 9432
rect 43211 9401 43223 9404
rect 43165 9395 43223 9401
rect 44082 9392 44088 9404
rect 44140 9392 44146 9444
rect 43254 9364 43260 9376
rect 42812 9336 43260 9364
rect 43254 9324 43260 9336
rect 43312 9324 43318 9376
rect 47210 9324 47216 9376
rect 47268 9324 47274 9376
rect 48038 9324 48044 9376
rect 48096 9324 48102 9376
rect 48222 9324 48228 9376
rect 48280 9364 48286 9376
rect 48777 9367 48835 9373
rect 48777 9364 48789 9367
rect 48280 9336 48789 9364
rect 48280 9324 48286 9336
rect 48777 9333 48789 9336
rect 48823 9333 48835 9367
rect 48777 9327 48835 9333
rect 50154 9324 50160 9376
rect 50212 9364 50218 9376
rect 51092 9364 51120 9460
rect 51166 9392 51172 9444
rect 51224 9432 51230 9444
rect 51718 9432 51724 9444
rect 51224 9404 51724 9432
rect 51224 9392 51230 9404
rect 51718 9392 51724 9404
rect 51776 9392 51782 9444
rect 53852 9376 53880 9472
rect 54021 9469 54033 9472
rect 54067 9469 54079 9503
rect 55309 9503 55367 9509
rect 55309 9500 55321 9503
rect 54021 9463 54079 9469
rect 54680 9472 55321 9500
rect 54680 9441 54708 9472
rect 55309 9469 55321 9472
rect 55355 9469 55367 9503
rect 55309 9463 55367 9469
rect 55490 9460 55496 9512
rect 55548 9460 55554 9512
rect 56318 9460 56324 9512
rect 56376 9460 56382 9512
rect 57072 9509 57100 9540
rect 56965 9503 57023 9509
rect 56965 9469 56977 9503
rect 57011 9469 57023 9503
rect 56965 9463 57023 9469
rect 57057 9503 57115 9509
rect 57057 9469 57069 9503
rect 57103 9469 57115 9503
rect 57057 9463 57115 9469
rect 54665 9435 54723 9441
rect 54665 9401 54677 9435
rect 54711 9401 54723 9435
rect 56980 9432 57008 9463
rect 57146 9432 57152 9444
rect 56980 9404 57152 9432
rect 54665 9395 54723 9401
rect 57146 9392 57152 9404
rect 57204 9392 57210 9444
rect 50212 9336 51120 9364
rect 50212 9324 50218 9336
rect 51902 9324 51908 9376
rect 51960 9324 51966 9376
rect 53834 9324 53840 9376
rect 53892 9324 53898 9376
rect 54754 9324 54760 9376
rect 54812 9324 54818 9376
rect 56226 9324 56232 9376
rect 56284 9364 56290 9376
rect 56505 9367 56563 9373
rect 56505 9364 56517 9367
rect 56284 9336 56517 9364
rect 56284 9324 56290 9336
rect 56505 9333 56517 9336
rect 56551 9333 56563 9367
rect 56505 9327 56563 9333
rect 1104 9274 58880 9296
rect 1104 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 22616 9274
rect 22668 9222 22680 9274
rect 22732 9222 22744 9274
rect 22796 9222 22808 9274
rect 22860 9222 22872 9274
rect 22924 9222 37060 9274
rect 37112 9222 37124 9274
rect 37176 9222 37188 9274
rect 37240 9222 37252 9274
rect 37304 9222 37316 9274
rect 37368 9222 51504 9274
rect 51556 9222 51568 9274
rect 51620 9222 51632 9274
rect 51684 9222 51696 9274
rect 51748 9222 51760 9274
rect 51812 9222 58880 9274
rect 1104 9200 58880 9222
rect 3142 9120 3148 9172
rect 3200 9120 3206 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 4062 9160 4068 9172
rect 3559 9132 4068 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3160 9064 3893 9092
rect 3160 9036 3188 9064
rect 3881 9061 3893 9064
rect 3927 9092 3939 9095
rect 5828 9092 5856 9123
rect 6546 9120 6552 9172
rect 6604 9120 6610 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7374 9160 7380 9172
rect 7055 9132 7380 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7708 9132 7849 9160
rect 7708 9120 7714 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10100 9132 10701 9160
rect 10100 9120 10106 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 10796 9132 12434 9160
rect 6178 9092 6184 9104
rect 3927 9064 6184 9092
rect 3927 9061 3939 9064
rect 3881 9055 3939 9061
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 6641 9095 6699 9101
rect 6641 9061 6653 9095
rect 6687 9092 6699 9095
rect 6687 9064 6960 9092
rect 6687 9061 6699 9064
rect 6641 9055 6699 9061
rect 6932 9036 6960 9064
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 7248 9064 7481 9092
rect 7248 9052 7254 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 8570 9092 8576 9104
rect 7469 9055 7527 9061
rect 7576 9064 8576 9092
rect 2685 9027 2743 9033
rect 2685 9024 2697 9027
rect 2332 8996 2697 9024
rect 2332 8832 2360 8996
rect 2685 8993 2697 8996
rect 2731 9024 2743 9027
rect 2731 8996 3096 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 3068 8956 3096 8996
rect 3142 8984 3148 9036
rect 3200 8984 3206 9036
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4304 8996 4629 9024
rect 4304 8984 4310 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 4663 8996 6224 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 3234 8956 3240 8968
rect 3068 8928 3240 8956
rect 2777 8919 2835 8925
rect 2792 8888 2820 8919
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8956 3387 8959
rect 3786 8956 3792 8968
rect 3375 8928 3792 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3344 8888 3372 8919
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8925 6147 8959
rect 6196 8956 6224 8996
rect 6730 8984 6736 9036
rect 6788 8984 6794 9036
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 7208 8956 7236 9052
rect 6196 8928 7236 8956
rect 6089 8919 6147 8925
rect 2792 8860 3372 8888
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 2314 8780 2320 8832
rect 2372 8780 2378 8832
rect 3528 8820 3556 8851
rect 5258 8848 5264 8900
rect 5316 8888 5322 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 5316 8860 5457 8888
rect 5316 8848 5322 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 6104 8888 6132 8919
rect 7576 8888 7604 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 8665 9095 8723 9101
rect 8665 9061 8677 9095
rect 8711 9092 8723 9095
rect 9214 9092 9220 9104
rect 8711 9064 9220 9092
rect 8711 9061 8723 9064
rect 8665 9055 8723 9061
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 10796 9024 10824 9132
rect 12406 9092 12434 9132
rect 14366 9120 14372 9172
rect 14424 9160 14430 9172
rect 14737 9163 14795 9169
rect 14737 9160 14749 9163
rect 14424 9132 14749 9160
rect 14424 9120 14430 9132
rect 14737 9129 14749 9132
rect 14783 9129 14795 9163
rect 14737 9123 14795 9129
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15344 9132 15424 9160
rect 15344 9120 15350 9132
rect 12406 9064 15240 9092
rect 8343 8996 10824 9024
rect 12069 9027 12127 9033
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 9048 8965 9076 8996
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12342 9024 12348 9036
rect 12115 8996 12348 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12342 8984 12348 8996
rect 12400 9024 12406 9036
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 12400 8996 13737 9024
rect 12400 8984 12406 8996
rect 13725 8993 13737 8996
rect 13771 9024 13783 9027
rect 13814 9024 13820 9036
rect 13771 8996 13820 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 13814 8984 13820 8996
rect 13872 9024 13878 9036
rect 14274 9024 14280 9036
rect 13872 8996 14280 9024
rect 13872 8984 13878 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 6104 8860 7604 8888
rect 7668 8928 8401 8956
rect 5445 8851 5503 8857
rect 7668 8832 7696 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11900 8928 12633 8956
rect 7742 8848 7748 8900
rect 7800 8848 7806 8900
rect 8220 8860 8616 8888
rect 8220 8832 8248 8860
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3528 8792 3801 8820
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 5822 8823 5880 8829
rect 5822 8789 5834 8823
rect 5868 8820 5880 8823
rect 6362 8820 6368 8832
rect 5868 8792 6368 8820
rect 5868 8789 5880 8792
rect 5822 8783 5880 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 7650 8780 7656 8832
rect 7708 8780 7714 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 8588 8820 8616 8860
rect 8662 8848 8668 8900
rect 8720 8848 8726 8900
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 8812 8860 9597 8888
rect 8812 8848 8818 8860
rect 9585 8857 9597 8860
rect 9631 8888 9643 8891
rect 10502 8888 10508 8900
rect 9631 8860 10508 8888
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 10597 8891 10655 8897
rect 10597 8857 10609 8891
rect 10643 8888 10655 8891
rect 11802 8891 11860 8897
rect 11802 8888 11814 8891
rect 10643 8860 11814 8888
rect 10643 8857 10655 8860
rect 10597 8851 10655 8857
rect 11802 8857 11814 8860
rect 11848 8857 11860 8891
rect 11802 8851 11860 8857
rect 11238 8820 11244 8832
rect 8588 8792 11244 8820
rect 11238 8780 11244 8792
rect 11296 8820 11302 8832
rect 11900 8820 11928 8928
rect 12621 8925 12633 8928
rect 12667 8956 12679 8959
rect 12667 8928 15148 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 12492 8860 13277 8888
rect 12492 8848 12498 8860
rect 13265 8857 13277 8860
rect 13311 8888 13323 8891
rect 14458 8888 14464 8900
rect 13311 8860 14464 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 11296 8792 11928 8820
rect 15120 8820 15148 8928
rect 15212 8888 15240 9064
rect 15396 9033 15424 9132
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 16117 9163 16175 9169
rect 15528 9132 15608 9160
rect 15528 9120 15534 9132
rect 15580 9033 15608 9132
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16574 9160 16580 9172
rect 16163 9132 16580 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9160 18199 9163
rect 18230 9160 18236 9172
rect 18187 9132 18236 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 18472 9132 18521 9160
rect 18472 9120 18478 9132
rect 18509 9129 18521 9132
rect 18555 9160 18567 9163
rect 20254 9160 20260 9172
rect 18555 9132 20260 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20438 9120 20444 9172
rect 20496 9120 20502 9172
rect 21361 9163 21419 9169
rect 21361 9129 21373 9163
rect 21407 9160 21419 9163
rect 22278 9160 22284 9172
rect 21407 9132 22284 9160
rect 21407 9129 21419 9132
rect 21361 9123 21419 9129
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 22370 9120 22376 9172
rect 22428 9120 22434 9172
rect 23290 9120 23296 9172
rect 23348 9120 23354 9172
rect 23750 9120 23756 9172
rect 23808 9160 23814 9172
rect 23845 9163 23903 9169
rect 23845 9160 23857 9163
rect 23808 9132 23857 9160
rect 23808 9120 23814 9132
rect 23845 9129 23857 9132
rect 23891 9129 23903 9163
rect 23845 9123 23903 9129
rect 27709 9163 27767 9169
rect 27709 9129 27721 9163
rect 27755 9160 27767 9163
rect 27798 9160 27804 9172
rect 27755 9132 27804 9160
rect 27755 9129 27767 9132
rect 27709 9123 27767 9129
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 29730 9120 29736 9172
rect 29788 9160 29794 9172
rect 30101 9163 30159 9169
rect 30101 9160 30113 9163
rect 29788 9132 30113 9160
rect 29788 9120 29794 9132
rect 30101 9129 30113 9132
rect 30147 9129 30159 9163
rect 30101 9123 30159 9129
rect 31297 9163 31355 9169
rect 31297 9129 31309 9163
rect 31343 9160 31355 9163
rect 32674 9160 32680 9172
rect 31343 9132 32680 9160
rect 31343 9129 31355 9132
rect 31297 9123 31355 9129
rect 32674 9120 32680 9132
rect 32732 9120 32738 9172
rect 34422 9120 34428 9172
rect 34480 9120 34486 9172
rect 34790 9120 34796 9172
rect 34848 9160 34854 9172
rect 34885 9163 34943 9169
rect 34885 9160 34897 9163
rect 34848 9132 34897 9160
rect 34848 9120 34854 9132
rect 34885 9129 34897 9132
rect 34931 9129 34943 9163
rect 34885 9123 34943 9129
rect 36265 9163 36323 9169
rect 36265 9129 36277 9163
rect 36311 9160 36323 9163
rect 36538 9160 36544 9172
rect 36311 9132 36544 9160
rect 36311 9129 36323 9132
rect 36265 9123 36323 9129
rect 36538 9120 36544 9132
rect 36596 9120 36602 9172
rect 38197 9163 38255 9169
rect 38197 9129 38209 9163
rect 38243 9160 38255 9163
rect 38286 9160 38292 9172
rect 38243 9132 38292 9160
rect 38243 9129 38255 9132
rect 38197 9123 38255 9129
rect 38286 9120 38292 9132
rect 38344 9120 38350 9172
rect 38470 9120 38476 9172
rect 38528 9120 38534 9172
rect 38580 9132 51488 9160
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 8993 15623 9027
rect 16684 9024 16712 9120
rect 19886 9052 19892 9104
rect 19944 9052 19950 9104
rect 20456 9033 20484 9120
rect 38580 9092 38608 9132
rect 20548 9064 38608 9092
rect 43073 9095 43131 9101
rect 17497 9027 17555 9033
rect 17497 9024 17509 9027
rect 16684 8996 17509 9024
rect 15565 8987 15623 8993
rect 17497 8993 17509 8996
rect 17543 8993 17555 9027
rect 17497 8987 17555 8993
rect 20441 9027 20499 9033
rect 20441 8993 20453 9027
rect 20487 8993 20499 9027
rect 20441 8987 20499 8993
rect 20548 8956 20576 9064
rect 43073 9061 43085 9095
rect 43119 9092 43131 9095
rect 43254 9092 43260 9104
rect 43119 9064 43260 9092
rect 43119 9061 43131 9064
rect 43073 9055 43131 9061
rect 43254 9052 43260 9064
rect 43312 9052 43318 9104
rect 48038 9092 48044 9104
rect 46952 9064 48044 9092
rect 20806 8984 20812 9036
rect 20864 8984 20870 9036
rect 21729 9027 21787 9033
rect 21729 8993 21741 9027
rect 21775 9024 21787 9027
rect 21775 8996 22094 9024
rect 21775 8993 21787 8996
rect 21729 8987 21787 8993
rect 16408 8928 20576 8956
rect 22066 8956 22094 8996
rect 22370 8984 22376 9036
rect 22428 9024 22434 9036
rect 22649 9027 22707 9033
rect 22649 9024 22661 9027
rect 22428 8996 22661 9024
rect 22428 8984 22434 8996
rect 22649 8993 22661 8996
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 23382 9024 23388 9036
rect 22879 8996 23388 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 26329 9027 26387 9033
rect 26329 9024 26341 9027
rect 24872 8996 26341 9024
rect 23106 8956 23112 8968
rect 22066 8928 23112 8956
rect 16298 8888 16304 8900
rect 15212 8860 16304 8888
rect 16298 8848 16304 8860
rect 16356 8848 16362 8900
rect 16408 8820 16436 8928
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 19705 8891 19763 8897
rect 19705 8888 19717 8891
rect 16540 8860 19717 8888
rect 16540 8848 16546 8860
rect 19705 8857 19717 8860
rect 19751 8888 19763 8891
rect 20622 8888 20628 8900
rect 19751 8860 20628 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 20622 8848 20628 8860
rect 20680 8888 20686 8900
rect 24872 8897 24900 8996
rect 26329 8993 26341 8996
rect 26375 8993 26387 9027
rect 26329 8987 26387 8993
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 26973 9027 27031 9033
rect 26973 9024 26985 9027
rect 26660 8996 26985 9024
rect 26660 8984 26666 8996
rect 26973 8993 26985 8996
rect 27019 8993 27031 9027
rect 26973 8987 27031 8993
rect 27617 9027 27675 9033
rect 27617 8993 27629 9027
rect 27663 9024 27675 9027
rect 27982 9024 27988 9036
rect 27663 8996 27988 9024
rect 27663 8993 27675 8996
rect 27617 8987 27675 8993
rect 27982 8984 27988 8996
rect 28040 8984 28046 9036
rect 28258 9024 28264 9036
rect 28092 8996 28264 9024
rect 25130 8916 25136 8968
rect 25188 8916 25194 8968
rect 26145 8959 26203 8965
rect 26145 8925 26157 8959
rect 26191 8956 26203 8959
rect 27706 8956 27712 8968
rect 26191 8928 27712 8956
rect 26191 8925 26203 8928
rect 26145 8919 26203 8925
rect 27706 8916 27712 8928
rect 27764 8916 27770 8968
rect 27890 8916 27896 8968
rect 27948 8956 27954 8968
rect 28092 8956 28120 8996
rect 28258 8984 28264 8996
rect 28316 8984 28322 9036
rect 28534 8984 28540 9036
rect 28592 8984 28598 9036
rect 30466 8984 30472 9036
rect 30524 8984 30530 9036
rect 30745 9027 30803 9033
rect 30745 8993 30757 9027
rect 30791 9024 30803 9027
rect 31662 9024 31668 9036
rect 30791 8996 31668 9024
rect 30791 8993 30803 8996
rect 30745 8987 30803 8993
rect 31662 8984 31668 8996
rect 31720 8984 31726 9036
rect 32769 9027 32827 9033
rect 32769 8993 32781 9027
rect 32815 9024 32827 9027
rect 33226 9024 33232 9036
rect 32815 8996 33232 9024
rect 32815 8993 32827 8996
rect 32769 8987 32827 8993
rect 33226 8984 33232 8996
rect 33284 8984 33290 9036
rect 34882 8984 34888 9036
rect 34940 9024 34946 9036
rect 35897 9027 35955 9033
rect 35897 9024 35909 9027
rect 34940 8996 35909 9024
rect 34940 8984 34946 8996
rect 35897 8993 35909 8996
rect 35943 8993 35955 9027
rect 35897 8987 35955 8993
rect 35986 8984 35992 9036
rect 36044 9024 36050 9036
rect 36906 9024 36912 9036
rect 36044 8996 36912 9024
rect 36044 8984 36050 8996
rect 36906 8984 36912 8996
rect 36964 8984 36970 9036
rect 42242 9024 42248 9036
rect 41386 8996 42248 9024
rect 27948 8928 28120 8956
rect 28169 8959 28227 8965
rect 27948 8916 27954 8928
rect 28169 8925 28181 8959
rect 28215 8956 28227 8959
rect 28718 8956 28724 8968
rect 28215 8928 28724 8956
rect 28215 8925 28227 8928
rect 28169 8919 28227 8925
rect 28718 8916 28724 8928
rect 28776 8956 28782 8968
rect 29181 8959 29239 8965
rect 29181 8956 29193 8959
rect 28776 8928 29193 8956
rect 28776 8916 28782 8928
rect 29181 8925 29193 8928
rect 29227 8925 29239 8959
rect 30484 8956 30512 8984
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 30484 8928 30849 8956
rect 29181 8919 29239 8925
rect 30837 8925 30849 8928
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 32950 8916 32956 8968
rect 33008 8916 33014 8968
rect 33318 8916 33324 8968
rect 33376 8956 33382 8968
rect 34330 8956 34336 8968
rect 33376 8928 34336 8956
rect 33376 8916 33382 8928
rect 34330 8916 34336 8928
rect 34388 8956 34394 8968
rect 34388 8928 35756 8956
rect 34388 8916 34394 8928
rect 24857 8891 24915 8897
rect 24857 8888 24869 8891
rect 20680 8860 24869 8888
rect 20680 8848 20686 8860
rect 24857 8857 24869 8860
rect 24903 8857 24915 8891
rect 24857 8851 24915 8857
rect 26881 8891 26939 8897
rect 26881 8857 26893 8891
rect 26927 8888 26939 8891
rect 27062 8888 27068 8900
rect 26927 8860 27068 8888
rect 26927 8857 26939 8860
rect 26881 8851 26939 8857
rect 27062 8848 27068 8860
rect 27120 8888 27126 8900
rect 28258 8888 28264 8900
rect 27120 8860 28264 8888
rect 27120 8848 27126 8860
rect 28258 8848 28264 8860
rect 28316 8848 28322 8900
rect 30929 8891 30987 8897
rect 30929 8857 30941 8891
rect 30975 8888 30987 8891
rect 31938 8888 31944 8900
rect 30975 8860 31944 8888
rect 30975 8857 30987 8860
rect 30929 8851 30987 8857
rect 31938 8848 31944 8860
rect 31996 8848 32002 8900
rect 34606 8888 34612 8900
rect 33336 8860 34612 8888
rect 15120 8792 16436 8820
rect 11296 8780 11302 8792
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 22925 8823 22983 8829
rect 22925 8820 22937 8823
rect 22336 8792 22937 8820
rect 22336 8780 22342 8792
rect 22925 8789 22937 8792
rect 22971 8820 22983 8823
rect 23198 8820 23204 8832
rect 22971 8792 23204 8820
rect 22971 8789 22983 8792
rect 22925 8783 22983 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 26237 8823 26295 8829
rect 26237 8789 26249 8823
rect 26283 8820 26295 8823
rect 26326 8820 26332 8832
rect 26283 8792 26332 8820
rect 26283 8789 26295 8792
rect 26237 8783 26295 8789
rect 26326 8780 26332 8792
rect 26384 8820 26390 8832
rect 28077 8823 28135 8829
rect 28077 8820 28089 8823
rect 26384 8792 28089 8820
rect 26384 8780 26390 8792
rect 28077 8789 28089 8792
rect 28123 8820 28135 8823
rect 28626 8820 28632 8832
rect 28123 8792 28632 8820
rect 28123 8789 28135 8792
rect 28077 8783 28135 8789
rect 28626 8780 28632 8792
rect 28684 8820 28690 8832
rect 29178 8820 29184 8832
rect 28684 8792 29184 8820
rect 28684 8780 28690 8792
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 31662 8780 31668 8832
rect 31720 8820 31726 8832
rect 33336 8829 33364 8860
rect 34606 8848 34612 8860
rect 34664 8848 34670 8900
rect 35728 8888 35756 8928
rect 36354 8916 36360 8968
rect 36412 8916 36418 8968
rect 36814 8916 36820 8968
rect 36872 8956 36878 8968
rect 37185 8959 37243 8965
rect 37185 8956 37197 8959
rect 36872 8928 37197 8956
rect 36872 8916 36878 8928
rect 37185 8925 37197 8928
rect 37231 8925 37243 8959
rect 38933 8959 38991 8965
rect 38933 8956 38945 8959
rect 37185 8919 37243 8925
rect 37568 8928 38945 8956
rect 37568 8900 37596 8928
rect 38933 8925 38945 8928
rect 38979 8956 38991 8959
rect 39666 8956 39672 8968
rect 38979 8928 39672 8956
rect 38979 8925 38991 8928
rect 38933 8919 38991 8925
rect 39666 8916 39672 8928
rect 39724 8956 39730 8968
rect 41386 8956 41414 8996
rect 42242 8984 42248 8996
rect 42300 9024 42306 9036
rect 46952 9024 46980 9064
rect 48038 9052 48044 9064
rect 48096 9092 48102 9104
rect 50062 9092 50068 9104
rect 48096 9064 50068 9092
rect 48096 9052 48102 9064
rect 42300 8996 46980 9024
rect 42300 8984 42306 8996
rect 47026 8984 47032 9036
rect 47084 8984 47090 9036
rect 47854 8984 47860 9036
rect 47912 9024 47918 9036
rect 48516 9033 48544 9064
rect 50062 9052 50068 9064
rect 50120 9052 50126 9104
rect 48133 9027 48191 9033
rect 48133 9024 48145 9027
rect 47912 8996 48145 9024
rect 47912 8984 47918 8996
rect 48133 8993 48145 8996
rect 48179 8993 48191 9027
rect 48133 8987 48191 8993
rect 48501 9027 48559 9033
rect 48501 8993 48513 9027
rect 48547 9024 48559 9027
rect 48547 8996 48581 9024
rect 48547 8993 48559 8996
rect 48501 8987 48559 8993
rect 48682 8984 48688 9036
rect 48740 8984 48746 9036
rect 50154 8984 50160 9036
rect 50212 8984 50218 9036
rect 39724 8928 41414 8956
rect 39724 8916 39730 8928
rect 45646 8916 45652 8968
rect 45704 8956 45710 8968
rect 45925 8959 45983 8965
rect 45925 8956 45937 8959
rect 45704 8928 45937 8956
rect 45704 8916 45710 8928
rect 45925 8925 45937 8928
rect 45971 8925 45983 8959
rect 45925 8919 45983 8925
rect 46290 8916 46296 8968
rect 46348 8956 46354 8968
rect 46658 8956 46664 8968
rect 46348 8928 46664 8956
rect 46348 8916 46354 8928
rect 46658 8916 46664 8928
rect 46716 8916 46722 8968
rect 48593 8959 48651 8965
rect 48593 8925 48605 8959
rect 48639 8956 48651 8959
rect 48700 8956 48728 8984
rect 48639 8928 48728 8956
rect 49697 8959 49755 8965
rect 48639 8925 48651 8928
rect 48593 8919 48651 8925
rect 49697 8925 49709 8959
rect 49743 8925 49755 8959
rect 51460 8956 51488 9132
rect 53282 9120 53288 9172
rect 53340 9120 53346 9172
rect 55582 9120 55588 9172
rect 55640 9120 55646 9172
rect 56226 9120 56232 9172
rect 56284 9120 56290 9172
rect 56321 9163 56379 9169
rect 56321 9129 56333 9163
rect 56367 9160 56379 9163
rect 56594 9160 56600 9172
rect 56367 9132 56600 9160
rect 56367 9129 56379 9132
rect 56321 9123 56379 9129
rect 56594 9120 56600 9132
rect 56652 9120 56658 9172
rect 51537 9095 51595 9101
rect 51537 9061 51549 9095
rect 51583 9092 51595 9095
rect 53300 9092 53328 9120
rect 51583 9064 53328 9092
rect 51583 9061 51595 9064
rect 51537 9055 51595 9061
rect 51902 8984 51908 9036
rect 51960 9024 51966 9036
rect 52181 9027 52239 9033
rect 52181 9024 52193 9027
rect 51960 8996 52193 9024
rect 51960 8984 51966 8996
rect 52181 8993 52193 8996
rect 52227 8993 52239 9027
rect 52181 8987 52239 8993
rect 55769 9027 55827 9033
rect 55769 8993 55781 9027
rect 55815 9024 55827 9027
rect 56244 9024 56272 9120
rect 55815 8996 56272 9024
rect 55815 8993 55827 8996
rect 55769 8987 55827 8993
rect 55950 8956 55956 8968
rect 51460 8928 55956 8956
rect 49697 8919 49755 8925
rect 37550 8888 37556 8900
rect 35728 8860 37556 8888
rect 37550 8848 37556 8860
rect 37608 8848 37614 8900
rect 38565 8891 38623 8897
rect 38565 8857 38577 8891
rect 38611 8888 38623 8891
rect 39482 8888 39488 8900
rect 38611 8860 39488 8888
rect 38611 8857 38623 8860
rect 38565 8851 38623 8857
rect 39482 8848 39488 8860
rect 39540 8848 39546 8900
rect 47210 8888 47216 8900
rect 44928 8860 47216 8888
rect 44928 8832 44956 8860
rect 47210 8848 47216 8860
rect 47268 8888 47274 8900
rect 47305 8891 47363 8897
rect 47305 8888 47317 8891
rect 47268 8860 47317 8888
rect 47268 8848 47274 8860
rect 47305 8857 47317 8860
rect 47351 8857 47363 8891
rect 48685 8891 48743 8897
rect 48685 8888 48697 8891
rect 47305 8851 47363 8857
rect 48424 8860 48697 8888
rect 32861 8823 32919 8829
rect 32861 8820 32873 8823
rect 31720 8792 32873 8820
rect 31720 8780 31726 8792
rect 32861 8789 32873 8792
rect 32907 8789 32919 8823
rect 32861 8783 32919 8789
rect 33321 8823 33379 8829
rect 33321 8789 33333 8823
rect 33367 8789 33379 8823
rect 33321 8783 33379 8789
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 33597 8823 33655 8829
rect 33597 8820 33609 8823
rect 33468 8792 33609 8820
rect 33468 8780 33474 8792
rect 33597 8789 33609 8792
rect 33643 8789 33655 8823
rect 33597 8783 33655 8789
rect 34057 8823 34115 8829
rect 34057 8789 34069 8823
rect 34103 8820 34115 8823
rect 34146 8820 34152 8832
rect 34103 8792 34152 8820
rect 34103 8789 34115 8792
rect 34057 8783 34115 8789
rect 34146 8780 34152 8792
rect 34204 8780 34210 8832
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 36538 8780 36544 8832
rect 36596 8820 36602 8832
rect 37001 8823 37059 8829
rect 37001 8820 37013 8823
rect 36596 8792 37013 8820
rect 36596 8780 36602 8792
rect 37001 8789 37013 8792
rect 37047 8789 37059 8823
rect 37001 8783 37059 8789
rect 37826 8780 37832 8832
rect 37884 8780 37890 8832
rect 44910 8780 44916 8832
rect 44968 8780 44974 8832
rect 45370 8780 45376 8832
rect 45428 8780 45434 8832
rect 46290 8780 46296 8832
rect 46348 8780 46354 8832
rect 46477 8823 46535 8829
rect 46477 8789 46489 8823
rect 46523 8820 46535 8823
rect 46658 8820 46664 8832
rect 46523 8792 46664 8820
rect 46523 8789 46535 8792
rect 46477 8783 46535 8789
rect 46658 8780 46664 8792
rect 46716 8780 46722 8832
rect 47762 8780 47768 8832
rect 47820 8820 47826 8832
rect 48222 8820 48228 8832
rect 47820 8792 48228 8820
rect 47820 8780 47826 8792
rect 48222 8780 48228 8792
rect 48280 8820 48286 8832
rect 48424 8820 48452 8860
rect 48685 8857 48697 8860
rect 48731 8857 48743 8891
rect 49712 8888 49740 8919
rect 55950 8916 55956 8928
rect 56008 8916 56014 8968
rect 56226 8916 56232 8968
rect 56284 8956 56290 8968
rect 56413 8959 56471 8965
rect 56413 8956 56425 8959
rect 56284 8928 56425 8956
rect 56284 8916 56290 8928
rect 56413 8925 56425 8928
rect 56459 8925 56471 8959
rect 56413 8919 56471 8925
rect 57146 8916 57152 8968
rect 57204 8956 57210 8968
rect 57885 8959 57943 8965
rect 57885 8956 57897 8959
rect 57204 8928 57897 8956
rect 57204 8916 57210 8928
rect 57885 8925 57897 8928
rect 57931 8925 57943 8959
rect 57885 8919 57943 8925
rect 58434 8916 58440 8968
rect 58492 8916 58498 8968
rect 48685 8851 48743 8857
rect 49068 8860 49740 8888
rect 50424 8891 50482 8897
rect 49068 8829 49096 8860
rect 50424 8857 50436 8891
rect 50470 8888 50482 8891
rect 51629 8891 51687 8897
rect 51629 8888 51641 8891
rect 50470 8860 51641 8888
rect 50470 8857 50482 8860
rect 50424 8851 50482 8857
rect 51629 8857 51641 8860
rect 51675 8857 51687 8891
rect 51629 8851 51687 8857
rect 53377 8891 53435 8897
rect 53377 8857 53389 8891
rect 53423 8857 53435 8891
rect 53377 8851 53435 8857
rect 48280 8792 48452 8820
rect 49053 8823 49111 8829
rect 48280 8780 48286 8792
rect 49053 8789 49065 8823
rect 49099 8789 49111 8823
rect 49053 8783 49111 8789
rect 49142 8780 49148 8832
rect 49200 8780 49206 8832
rect 53190 8780 53196 8832
rect 53248 8820 53254 8832
rect 53392 8820 53420 8851
rect 54294 8848 54300 8900
rect 54352 8888 54358 8900
rect 55125 8891 55183 8897
rect 55125 8888 55137 8891
rect 54352 8860 55137 8888
rect 54352 8848 54358 8860
rect 55125 8857 55137 8860
rect 55171 8888 55183 8891
rect 56244 8888 56272 8916
rect 55171 8860 56272 8888
rect 56680 8891 56738 8897
rect 55171 8857 55183 8860
rect 55125 8851 55183 8857
rect 56680 8857 56692 8891
rect 56726 8888 56738 8891
rect 57238 8888 57244 8900
rect 56726 8860 57244 8888
rect 56726 8857 56738 8860
rect 56680 8851 56738 8857
rect 57238 8848 57244 8860
rect 57296 8848 57302 8900
rect 53248 8792 53420 8820
rect 53248 8780 53254 8792
rect 57790 8780 57796 8832
rect 57848 8780 57854 8832
rect 1104 8730 59040 8752
rect 1104 8678 15394 8730
rect 15446 8678 15458 8730
rect 15510 8678 15522 8730
rect 15574 8678 15586 8730
rect 15638 8678 15650 8730
rect 15702 8678 29838 8730
rect 29890 8678 29902 8730
rect 29954 8678 29966 8730
rect 30018 8678 30030 8730
rect 30082 8678 30094 8730
rect 30146 8678 44282 8730
rect 44334 8678 44346 8730
rect 44398 8678 44410 8730
rect 44462 8678 44474 8730
rect 44526 8678 44538 8730
rect 44590 8678 58726 8730
rect 58778 8678 58790 8730
rect 58842 8678 58854 8730
rect 58906 8678 58918 8730
rect 58970 8678 58982 8730
rect 59034 8678 59040 8730
rect 1104 8656 59040 8678
rect 2314 8576 2320 8628
rect 2372 8576 2378 8628
rect 4246 8616 4252 8628
rect 3436 8588 4252 8616
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3436 8480 3464 8588
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 7653 8619 7711 8625
rect 7653 8585 7665 8619
rect 7699 8616 7711 8619
rect 7834 8616 7840 8628
rect 7699 8588 7840 8616
rect 7699 8585 7711 8588
rect 7653 8579 7711 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9490 8616 9496 8628
rect 8536 8588 9496 8616
rect 8536 8576 8542 8588
rect 9490 8576 9496 8588
rect 9548 8616 9554 8628
rect 9548 8588 9996 8616
rect 9548 8576 9554 8588
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 6730 8548 6736 8560
rect 5276 8520 6736 8548
rect 5276 8492 5304 8520
rect 3099 8452 3464 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 5258 8440 5264 8492
rect 5316 8440 5322 8492
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6656 8489 6684 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 7009 8551 7067 8557
rect 7009 8517 7021 8551
rect 7055 8548 7067 8551
rect 8202 8548 8208 8560
rect 7055 8520 8208 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 9858 8548 9864 8560
rect 8404 8520 9864 8548
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6420 8452 6561 8480
rect 6420 8440 6426 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 8404 8489 8432 8520
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 9968 8548 9996 8588
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10100 8588 10609 8616
rect 10100 8576 10106 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 12342 8616 12348 8628
rect 11020 8588 12348 8616
rect 11020 8576 11026 8588
rect 10229 8551 10287 8557
rect 10229 8548 10241 8551
rect 9968 8520 10241 8548
rect 10229 8517 10241 8520
rect 10275 8517 10287 8551
rect 10229 8511 10287 8517
rect 11054 8508 11060 8560
rect 11112 8508 11118 8560
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8656 8483 8714 8489
rect 8656 8449 8668 8483
rect 8702 8480 8714 8483
rect 8938 8480 8944 8492
rect 8702 8452 8944 8480
rect 8702 8449 8714 8452
rect 8656 8443 8714 8449
rect 3142 8372 3148 8424
rect 3200 8372 3206 8424
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6236 8384 7113 8412
rect 6236 8372 6242 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7208 8412 7236 8440
rect 7576 8412 7604 8443
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11072 8480 11100 8508
rect 11624 8489 11652 8588
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 14332 8588 14381 8616
rect 14332 8576 14338 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15838 8616 15844 8628
rect 15243 8588 15844 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 16264 8588 17325 8616
rect 16264 8576 16270 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17770 8616 17776 8628
rect 17727 8588 17776 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17770 8576 17776 8588
rect 17828 8616 17834 8628
rect 18046 8616 18052 8628
rect 17828 8588 18052 8616
rect 17828 8576 17834 8588
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20312 8588 20913 8616
rect 20312 8576 20318 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21542 8616 21548 8628
rect 21407 8588 21548 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 24857 8619 24915 8625
rect 24857 8585 24869 8619
rect 24903 8616 24915 8619
rect 25222 8616 25228 8628
rect 24903 8588 25228 8616
rect 24903 8585 24915 8588
rect 24857 8579 24915 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 25590 8576 25596 8628
rect 25648 8576 25654 8628
rect 26605 8619 26663 8625
rect 26605 8585 26617 8619
rect 26651 8616 26663 8619
rect 27154 8616 27160 8628
rect 26651 8588 27160 8616
rect 26651 8585 26663 8588
rect 26605 8579 26663 8585
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 27617 8619 27675 8625
rect 27617 8585 27629 8619
rect 27663 8616 27675 8619
rect 27706 8616 27712 8628
rect 27663 8588 27712 8616
rect 27663 8585 27675 8588
rect 27617 8579 27675 8585
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 27890 8576 27896 8628
rect 27948 8576 27954 8628
rect 31726 8588 45048 8616
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 11716 8520 13921 8548
rect 11011 8452 11100 8480
rect 11609 8483 11667 8489
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 7834 8412 7840 8424
rect 7208 8384 7840 8412
rect 7101 8375 7159 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 7469 8279 7527 8285
rect 7469 8245 7481 8279
rect 7515 8276 7527 8279
rect 7650 8276 7656 8288
rect 7515 8248 7656 8276
rect 7515 8245 7527 8248
rect 7469 8239 7527 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 8312 8276 8340 8375
rect 10226 8372 10232 8424
rect 10284 8372 10290 8424
rect 10336 8412 10364 8443
rect 10502 8412 10508 8424
rect 10336 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10928 8384 11069 8412
rect 10928 8372 10934 8384
rect 11057 8381 11069 8384
rect 11103 8381 11115 8415
rect 11057 8375 11115 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11716 8412 11744 8520
rect 13909 8517 13921 8520
rect 13955 8548 13967 8551
rect 14182 8548 14188 8560
rect 13955 8520 14188 8548
rect 13955 8517 13967 8520
rect 13909 8511 13967 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 14829 8551 14887 8557
rect 14829 8517 14841 8551
rect 14875 8548 14887 8551
rect 31726 8548 31754 8588
rect 14875 8520 31754 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 11876 8483 11934 8489
rect 11876 8449 11888 8483
rect 11922 8480 11934 8483
rect 12802 8480 12808 8492
rect 11922 8452 12808 8480
rect 11922 8449 11934 8452
rect 11876 8443 11934 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 14844 8480 14872 8511
rect 33042 8508 33048 8560
rect 33100 8548 33106 8560
rect 34149 8551 34207 8557
rect 34149 8548 34161 8551
rect 33100 8520 34161 8548
rect 33100 8508 33106 8520
rect 34149 8517 34161 8520
rect 34195 8517 34207 8551
rect 34149 8511 34207 8517
rect 34882 8508 34888 8560
rect 34940 8508 34946 8560
rect 35802 8508 35808 8560
rect 35860 8508 35866 8560
rect 35986 8508 35992 8560
rect 36044 8508 36050 8560
rect 36170 8508 36176 8560
rect 36228 8548 36234 8560
rect 38105 8551 38163 8557
rect 38105 8548 38117 8551
rect 36228 8520 36308 8548
rect 36228 8508 36234 8520
rect 13320 8452 14872 8480
rect 15488 8452 16068 8480
rect 13320 8440 13326 8452
rect 15488 8424 15516 8452
rect 11195 8384 11744 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8344 9827 8347
rect 10244 8344 10272 8372
rect 11164 8344 11192 8375
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 15470 8412 15476 8424
rect 14240 8384 15476 8412
rect 14240 8372 14246 8384
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15746 8372 15752 8424
rect 15804 8372 15810 8424
rect 16040 8412 16068 8452
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16172 8452 16681 8480
rect 16172 8440 16178 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 25498 8440 25504 8492
rect 25556 8440 25562 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 26145 8483 26203 8489
rect 26145 8480 26157 8483
rect 25832 8452 26157 8480
rect 25832 8440 25838 8452
rect 26145 8449 26157 8452
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 26418 8440 26424 8492
rect 26476 8480 26482 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26476 8452 26985 8480
rect 26476 8440 26482 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 28350 8440 28356 8492
rect 28408 8440 28414 8492
rect 32769 8483 32827 8489
rect 32769 8449 32781 8483
rect 32815 8449 32827 8483
rect 32769 8443 32827 8449
rect 18322 8412 18328 8424
rect 16040 8384 18328 8412
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 21174 8412 21180 8424
rect 19306 8384 21180 8412
rect 9815 8316 10272 8344
rect 10980 8316 11192 8344
rect 12989 8347 13047 8353
rect 9815 8313 9827 8316
rect 9769 8307 9827 8313
rect 8570 8276 8576 8288
rect 8312 8248 8576 8276
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 10980 8276 11008 8316
rect 12989 8313 13001 8347
rect 13035 8344 13047 8347
rect 13814 8344 13820 8356
rect 13035 8316 13820 8344
rect 13035 8313 13047 8316
rect 12989 8307 13047 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 18340 8344 18368 8372
rect 19306 8344 19334 8384
rect 21174 8372 21180 8384
rect 21232 8412 21238 8424
rect 21232 8384 22223 8412
rect 21232 8372 21238 8384
rect 14516 8316 17632 8344
rect 18340 8316 19334 8344
rect 14516 8304 14522 8316
rect 17604 8288 17632 8316
rect 22094 8304 22100 8356
rect 22152 8304 22158 8356
rect 22195 8344 22223 8384
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22649 8415 22707 8421
rect 22649 8412 22661 8415
rect 22520 8384 22661 8412
rect 22520 8372 22526 8384
rect 22649 8381 22661 8384
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 23382 8372 23388 8424
rect 23440 8372 23446 8424
rect 28902 8372 28908 8424
rect 28960 8412 28966 8424
rect 29365 8415 29423 8421
rect 29365 8412 29377 8415
rect 28960 8384 29377 8412
rect 28960 8372 28966 8384
rect 29365 8381 29377 8384
rect 29411 8381 29423 8415
rect 29365 8375 29423 8381
rect 30098 8372 30104 8424
rect 30156 8412 30162 8424
rect 30156 8384 30604 8412
rect 30156 8372 30162 8384
rect 24673 8347 24731 8353
rect 24673 8344 24685 8347
rect 22195 8316 24685 8344
rect 24673 8313 24685 8316
rect 24719 8344 24731 8347
rect 25958 8344 25964 8356
rect 24719 8316 25964 8344
rect 24719 8313 24731 8316
rect 24673 8307 24731 8313
rect 25958 8304 25964 8316
rect 26016 8344 26022 8356
rect 29917 8347 29975 8353
rect 29917 8344 29929 8347
rect 26016 8316 29929 8344
rect 26016 8304 26022 8316
rect 29917 8313 29929 8316
rect 29963 8344 29975 8347
rect 30466 8344 30472 8356
rect 29963 8316 30472 8344
rect 29963 8313 29975 8316
rect 29917 8307 29975 8313
rect 30466 8304 30472 8316
rect 30524 8304 30530 8356
rect 30576 8344 30604 8384
rect 30650 8372 30656 8424
rect 30708 8372 30714 8424
rect 31386 8372 31392 8424
rect 31444 8372 31450 8424
rect 31757 8347 31815 8353
rect 31757 8344 31769 8347
rect 30576 8316 31769 8344
rect 31757 8313 31769 8316
rect 31803 8344 31815 8347
rect 31938 8344 31944 8356
rect 31803 8316 31944 8344
rect 31803 8313 31815 8316
rect 31757 8307 31815 8313
rect 31938 8304 31944 8316
rect 31996 8304 32002 8356
rect 10928 8248 11008 8276
rect 10928 8236 10934 8248
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 16356 8248 16405 8276
rect 16356 8236 16362 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16393 8239 16451 8245
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 21818 8276 21824 8288
rect 17644 8248 21824 8276
rect 17644 8236 17650 8248
rect 21818 8236 21824 8248
rect 21876 8236 21882 8288
rect 22370 8236 22376 8288
rect 22428 8276 22434 8288
rect 22833 8279 22891 8285
rect 22833 8276 22845 8279
rect 22428 8248 22845 8276
rect 22428 8236 22434 8248
rect 22833 8245 22845 8248
rect 22879 8245 22891 8279
rect 22833 8239 22891 8245
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 26142 8276 26148 8288
rect 24820 8248 26148 8276
rect 24820 8236 24826 8248
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 27430 8236 27436 8288
rect 27488 8276 27494 8288
rect 28169 8279 28227 8285
rect 28169 8276 28181 8279
rect 27488 8248 28181 8276
rect 27488 8236 27494 8248
rect 28169 8245 28181 8248
rect 28215 8245 28227 8279
rect 28169 8239 28227 8245
rect 28718 8236 28724 8288
rect 28776 8276 28782 8288
rect 28813 8279 28871 8285
rect 28813 8276 28825 8279
rect 28776 8248 28825 8276
rect 28776 8236 28782 8248
rect 28813 8245 28825 8248
rect 28859 8245 28871 8279
rect 28813 8239 28871 8245
rect 30101 8279 30159 8285
rect 30101 8245 30113 8279
rect 30147 8276 30159 8279
rect 30282 8276 30288 8288
rect 30147 8248 30288 8276
rect 30147 8245 30159 8248
rect 30101 8239 30159 8245
rect 30282 8236 30288 8248
rect 30340 8236 30346 8288
rect 30837 8279 30895 8285
rect 30837 8245 30849 8279
rect 30883 8276 30895 8279
rect 30926 8276 30932 8288
rect 30883 8248 30932 8276
rect 30883 8245 30895 8248
rect 30837 8239 30895 8245
rect 30926 8236 30932 8248
rect 30984 8236 30990 8288
rect 32674 8236 32680 8288
rect 32732 8276 32738 8288
rect 32784 8276 32812 8443
rect 34330 8440 34336 8492
rect 34388 8440 34394 8492
rect 34514 8440 34520 8492
rect 34572 8440 34578 8492
rect 34900 8480 34928 8508
rect 35713 8483 35771 8489
rect 34900 8452 35388 8480
rect 33226 8372 33232 8424
rect 33284 8372 33290 8424
rect 33410 8372 33416 8424
rect 33468 8412 33474 8424
rect 33505 8415 33563 8421
rect 33505 8412 33517 8415
rect 33468 8384 33517 8412
rect 33468 8372 33474 8384
rect 33505 8381 33517 8384
rect 33551 8381 33563 8415
rect 33505 8375 33563 8381
rect 33244 8344 33272 8372
rect 33870 8344 33876 8356
rect 33244 8316 33876 8344
rect 33870 8304 33876 8316
rect 33928 8344 33934 8356
rect 33965 8347 34023 8353
rect 33965 8344 33977 8347
rect 33928 8316 33977 8344
rect 33928 8304 33934 8316
rect 33965 8313 33977 8316
rect 34011 8313 34023 8347
rect 33965 8307 34023 8313
rect 35158 8304 35164 8356
rect 35216 8304 35222 8356
rect 35360 8353 35388 8452
rect 35713 8449 35725 8483
rect 35759 8480 35771 8483
rect 36004 8480 36032 8508
rect 36280 8489 36308 8520
rect 36464 8520 38117 8548
rect 36464 8492 36492 8520
rect 38105 8517 38117 8520
rect 38151 8548 38163 8551
rect 38565 8551 38623 8557
rect 38565 8548 38577 8551
rect 38151 8520 38577 8548
rect 38151 8517 38163 8520
rect 38105 8511 38163 8517
rect 38565 8517 38577 8520
rect 38611 8517 38623 8551
rect 44910 8548 44916 8560
rect 38565 8511 38623 8517
rect 38672 8520 44916 8548
rect 35759 8452 36032 8480
rect 36265 8483 36323 8489
rect 35759 8449 35771 8452
rect 35713 8443 35771 8449
rect 36265 8449 36277 8483
rect 36311 8449 36323 8483
rect 36265 8443 36323 8449
rect 36446 8440 36452 8492
rect 36504 8440 36510 8492
rect 36998 8440 37004 8492
rect 37056 8480 37062 8492
rect 38672 8480 38700 8520
rect 44910 8508 44916 8520
rect 44968 8508 44974 8560
rect 37056 8452 38700 8480
rect 37056 8440 37062 8452
rect 40402 8440 40408 8492
rect 40460 8440 40466 8492
rect 42978 8440 42984 8492
rect 43036 8480 43042 8492
rect 44821 8483 44879 8489
rect 44821 8480 44833 8483
rect 43036 8452 44833 8480
rect 43036 8440 43042 8452
rect 44821 8449 44833 8452
rect 44867 8449 44879 8483
rect 45020 8480 45048 8588
rect 45370 8576 45376 8628
rect 45428 8576 45434 8628
rect 47581 8619 47639 8625
rect 47581 8585 47593 8619
rect 47627 8616 47639 8619
rect 48130 8616 48136 8628
rect 47627 8588 48136 8616
rect 47627 8585 47639 8588
rect 47581 8579 47639 8585
rect 48130 8576 48136 8588
rect 48188 8576 48194 8628
rect 49142 8576 49148 8628
rect 49200 8576 49206 8628
rect 51077 8619 51135 8625
rect 51077 8585 51089 8619
rect 51123 8616 51135 8619
rect 51258 8616 51264 8628
rect 51123 8588 51264 8616
rect 51123 8585 51135 8588
rect 51077 8579 51135 8585
rect 51258 8576 51264 8588
rect 51316 8576 51322 8628
rect 51721 8619 51779 8625
rect 51721 8585 51733 8619
rect 51767 8616 51779 8619
rect 52178 8616 52184 8628
rect 51767 8588 52184 8616
rect 51767 8585 51779 8588
rect 51721 8579 51779 8585
rect 52178 8576 52184 8588
rect 52236 8576 52242 8628
rect 54754 8576 54760 8628
rect 54812 8576 54818 8628
rect 54941 8619 54999 8625
rect 54941 8585 54953 8619
rect 54987 8616 54999 8619
rect 55490 8616 55496 8628
rect 54987 8588 55496 8616
rect 54987 8585 54999 8588
rect 54941 8579 54999 8585
rect 55490 8576 55496 8588
rect 55548 8576 55554 8628
rect 56778 8616 56784 8628
rect 55600 8588 56784 8616
rect 45088 8551 45146 8557
rect 45088 8517 45100 8551
rect 45134 8548 45146 8551
rect 45388 8548 45416 8576
rect 47213 8551 47271 8557
rect 45134 8520 45416 8548
rect 45480 8520 46520 8548
rect 45134 8517 45146 8520
rect 45088 8511 45146 8517
rect 45480 8480 45508 8520
rect 46290 8480 46296 8492
rect 45020 8452 45508 8480
rect 45848 8452 46296 8480
rect 44821 8443 44879 8449
rect 35434 8372 35440 8424
rect 35492 8412 35498 8424
rect 35897 8415 35955 8421
rect 35897 8412 35909 8415
rect 35492 8384 35909 8412
rect 35492 8372 35498 8384
rect 35897 8381 35909 8384
rect 35943 8412 35955 8415
rect 37090 8412 37096 8424
rect 35943 8384 37096 8412
rect 35943 8381 35955 8384
rect 35897 8375 35955 8381
rect 37090 8372 37096 8384
rect 37148 8372 37154 8424
rect 37550 8372 37556 8424
rect 37608 8412 37614 8424
rect 37829 8415 37887 8421
rect 37829 8412 37841 8415
rect 37608 8384 37841 8412
rect 37608 8372 37614 8384
rect 37829 8381 37841 8384
rect 37875 8381 37887 8415
rect 37829 8375 37887 8381
rect 37918 8372 37924 8424
rect 37976 8412 37982 8424
rect 38013 8415 38071 8421
rect 38013 8412 38025 8415
rect 37976 8384 38025 8412
rect 37976 8372 37982 8384
rect 38013 8381 38025 8384
rect 38059 8381 38071 8415
rect 38930 8412 38936 8424
rect 38013 8375 38071 8381
rect 38396 8384 38936 8412
rect 35345 8347 35403 8353
rect 35345 8313 35357 8347
rect 35391 8313 35403 8347
rect 35345 8307 35403 8313
rect 36817 8347 36875 8353
rect 36817 8313 36829 8347
rect 36863 8344 36875 8347
rect 36906 8344 36912 8356
rect 36863 8316 36912 8344
rect 36863 8313 36875 8316
rect 36817 8307 36875 8313
rect 36906 8304 36912 8316
rect 36964 8304 36970 8356
rect 36998 8304 37004 8356
rect 37056 8304 37062 8356
rect 37016 8276 37044 8304
rect 32732 8248 37044 8276
rect 32732 8236 32738 8248
rect 37090 8236 37096 8288
rect 37148 8276 37154 8288
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37148 8248 37473 8276
rect 37148 8236 37154 8248
rect 37461 8245 37473 8248
rect 37507 8276 37519 8279
rect 38396 8276 38424 8384
rect 38930 8372 38936 8384
rect 38988 8372 38994 8424
rect 39114 8372 39120 8424
rect 39172 8372 39178 8424
rect 39853 8415 39911 8421
rect 39853 8381 39865 8415
rect 39899 8381 39911 8415
rect 39853 8375 39911 8381
rect 38473 8347 38531 8353
rect 38473 8313 38485 8347
rect 38519 8344 38531 8347
rect 39868 8344 39896 8375
rect 43070 8372 43076 8424
rect 43128 8372 43134 8424
rect 44726 8372 44732 8424
rect 44784 8372 44790 8424
rect 38519 8316 39896 8344
rect 38519 8313 38531 8316
rect 38473 8307 38531 8313
rect 40218 8304 40224 8356
rect 40276 8344 40282 8356
rect 40494 8344 40500 8356
rect 40276 8316 40500 8344
rect 40276 8304 40282 8316
rect 40494 8304 40500 8316
rect 40552 8344 40558 8356
rect 41049 8347 41107 8353
rect 41049 8344 41061 8347
rect 40552 8316 41061 8344
rect 40552 8304 40558 8316
rect 41049 8313 41061 8316
rect 41095 8313 41107 8347
rect 44085 8347 44143 8353
rect 41049 8307 41107 8313
rect 42352 8316 42564 8344
rect 37507 8248 38424 8276
rect 37507 8245 37519 8248
rect 37461 8239 37519 8245
rect 39298 8236 39304 8288
rect 39356 8236 39362 8288
rect 42058 8236 42064 8288
rect 42116 8276 42122 8288
rect 42352 8276 42380 8316
rect 42116 8248 42380 8276
rect 42116 8236 42122 8248
rect 42426 8236 42432 8288
rect 42484 8236 42490 8288
rect 42536 8276 42564 8316
rect 43364 8316 44036 8344
rect 43364 8276 43392 8316
rect 42536 8248 43392 8276
rect 43441 8279 43499 8285
rect 43441 8245 43453 8279
rect 43487 8276 43499 8279
rect 43898 8276 43904 8288
rect 43487 8248 43904 8276
rect 43487 8245 43499 8248
rect 43441 8239 43499 8245
rect 43898 8236 43904 8248
rect 43956 8236 43962 8288
rect 44008 8276 44036 8316
rect 44085 8313 44097 8347
rect 44131 8344 44143 8347
rect 44174 8344 44180 8356
rect 44131 8316 44180 8344
rect 44131 8313 44143 8316
rect 44085 8307 44143 8313
rect 44174 8304 44180 8316
rect 44232 8304 44238 8356
rect 45848 8276 45876 8452
rect 46290 8440 46296 8452
rect 46348 8480 46354 8492
rect 46385 8483 46443 8489
rect 46385 8480 46397 8483
rect 46348 8452 46397 8480
rect 46348 8440 46354 8452
rect 46385 8449 46397 8452
rect 46431 8449 46443 8483
rect 46492 8480 46520 8520
rect 47213 8517 47225 8551
rect 47259 8548 47271 8551
rect 47670 8548 47676 8560
rect 47259 8520 47676 8548
rect 47259 8517 47271 8520
rect 47213 8511 47271 8517
rect 47670 8508 47676 8520
rect 47728 8508 47734 8560
rect 48716 8551 48774 8557
rect 48716 8517 48728 8551
rect 48762 8548 48774 8551
rect 49160 8548 49188 8576
rect 53828 8551 53886 8557
rect 48762 8520 49188 8548
rect 53576 8520 53788 8548
rect 48762 8517 48774 8520
rect 48716 8511 48774 8517
rect 51813 8483 51871 8489
rect 46492 8452 51074 8480
rect 46385 8443 46443 8449
rect 48961 8415 49019 8421
rect 48961 8381 48973 8415
rect 49007 8412 49019 8415
rect 50154 8412 50160 8424
rect 49007 8384 50160 8412
rect 49007 8381 49019 8384
rect 48961 8375 49019 8381
rect 50154 8372 50160 8384
rect 50212 8372 50218 8424
rect 50430 8372 50436 8424
rect 50488 8372 50494 8424
rect 51046 8344 51074 8452
rect 51813 8449 51825 8483
rect 51859 8480 51871 8483
rect 51902 8480 51908 8492
rect 51859 8452 51908 8480
rect 51859 8449 51871 8452
rect 51813 8443 51871 8449
rect 51902 8440 51908 8452
rect 51960 8440 51966 8492
rect 53576 8489 53604 8520
rect 53561 8483 53619 8489
rect 53561 8449 53573 8483
rect 53607 8449 53619 8483
rect 53561 8443 53619 8449
rect 53650 8440 53656 8492
rect 53708 8440 53714 8492
rect 53760 8480 53788 8520
rect 53828 8517 53840 8551
rect 53874 8548 53886 8551
rect 54772 8548 54800 8576
rect 53874 8520 54800 8548
rect 55401 8551 55459 8557
rect 53874 8517 53886 8520
rect 53828 8511 53886 8517
rect 55401 8517 55413 8551
rect 55447 8548 55459 8551
rect 55600 8548 55628 8588
rect 56778 8576 56784 8588
rect 56836 8576 56842 8628
rect 57146 8576 57152 8628
rect 57204 8576 57210 8628
rect 57238 8576 57244 8628
rect 57296 8616 57302 8628
rect 57885 8619 57943 8625
rect 57885 8616 57897 8619
rect 57296 8588 57897 8616
rect 57296 8576 57302 8588
rect 57885 8585 57897 8588
rect 57931 8585 57943 8619
rect 57885 8579 57943 8585
rect 55447 8520 55628 8548
rect 55447 8517 55459 8520
rect 55401 8511 55459 8517
rect 54294 8480 54300 8492
rect 53760 8452 54300 8480
rect 54294 8440 54300 8452
rect 54352 8440 54358 8492
rect 56134 8440 56140 8492
rect 56192 8489 56198 8492
rect 56192 8483 56241 8489
rect 56192 8449 56195 8483
rect 56229 8449 56241 8483
rect 57164 8480 57192 8576
rect 57241 8483 57299 8489
rect 57241 8480 57253 8483
rect 57164 8452 57253 8480
rect 56192 8443 56241 8449
rect 57241 8449 57253 8452
rect 57287 8449 57299 8483
rect 57241 8443 57299 8449
rect 56192 8440 56198 8443
rect 53374 8372 53380 8424
rect 53432 8372 53438 8424
rect 53668 8412 53696 8440
rect 53484 8384 53696 8412
rect 53484 8344 53512 8384
rect 55674 8372 55680 8424
rect 55732 8412 55738 8424
rect 56045 8415 56103 8421
rect 56045 8412 56057 8415
rect 55732 8384 56057 8412
rect 55732 8372 55738 8384
rect 56045 8381 56057 8384
rect 56091 8381 56103 8415
rect 56045 8375 56103 8381
rect 56321 8415 56379 8421
rect 56321 8381 56333 8415
rect 56367 8412 56379 8415
rect 56502 8412 56508 8424
rect 56367 8384 56508 8412
rect 56367 8381 56379 8384
rect 56321 8375 56379 8381
rect 56502 8372 56508 8384
rect 56560 8372 56566 8424
rect 57057 8415 57115 8421
rect 57057 8381 57069 8415
rect 57103 8381 57115 8415
rect 57057 8375 57115 8381
rect 51046 8316 53512 8344
rect 55306 8304 55312 8356
rect 55364 8344 55370 8356
rect 56597 8347 56655 8353
rect 56597 8344 56609 8347
rect 55364 8316 55720 8344
rect 55364 8304 55370 8316
rect 44008 8248 45876 8276
rect 46201 8279 46259 8285
rect 46201 8245 46213 8279
rect 46247 8276 46259 8279
rect 46474 8276 46480 8288
rect 46247 8248 46480 8276
rect 46247 8245 46259 8248
rect 46201 8239 46259 8245
rect 46474 8236 46480 8248
rect 46532 8236 46538 8288
rect 49878 8236 49884 8288
rect 49936 8236 49942 8288
rect 50062 8236 50068 8288
rect 50120 8276 50126 8288
rect 52365 8279 52423 8285
rect 52365 8276 52377 8279
rect 50120 8248 52377 8276
rect 50120 8236 50126 8248
rect 52365 8245 52377 8248
rect 52411 8276 52423 8279
rect 52638 8276 52644 8288
rect 52411 8248 52644 8276
rect 52411 8245 52423 8248
rect 52365 8239 52423 8245
rect 52638 8236 52644 8248
rect 52696 8236 52702 8288
rect 52822 8236 52828 8288
rect 52880 8236 52886 8288
rect 55692 8276 55720 8316
rect 56520 8316 56609 8344
rect 56520 8276 56548 8316
rect 56597 8313 56609 8316
rect 56643 8344 56655 8347
rect 56870 8344 56876 8356
rect 56643 8316 56876 8344
rect 56643 8313 56655 8316
rect 56597 8307 56655 8313
rect 56870 8304 56876 8316
rect 56928 8304 56934 8356
rect 57072 8344 57100 8375
rect 57882 8372 57888 8424
rect 57940 8412 57946 8424
rect 58437 8415 58495 8421
rect 58437 8412 58449 8415
rect 57940 8384 58449 8412
rect 57940 8372 57946 8384
rect 58437 8381 58449 8384
rect 58483 8381 58495 8415
rect 58437 8375 58495 8381
rect 58158 8344 58164 8356
rect 57072 8316 58164 8344
rect 58158 8304 58164 8316
rect 58216 8304 58222 8356
rect 55692 8248 56548 8276
rect 1104 8186 58880 8208
rect 1104 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 22616 8186
rect 22668 8134 22680 8186
rect 22732 8134 22744 8186
rect 22796 8134 22808 8186
rect 22860 8134 22872 8186
rect 22924 8134 37060 8186
rect 37112 8134 37124 8186
rect 37176 8134 37188 8186
rect 37240 8134 37252 8186
rect 37304 8134 37316 8186
rect 37368 8134 51504 8186
rect 51556 8134 51568 8186
rect 51620 8134 51632 8186
rect 51684 8134 51696 8186
rect 51748 8134 51760 8186
rect 51812 8134 58880 8186
rect 1104 8112 58880 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3510 8072 3516 8084
rect 3467 8044 3516 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8628 8044 8953 8072
rect 8628 8032 8634 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 13262 8072 13268 8084
rect 8941 8035 8999 8041
rect 9416 8044 13268 8072
rect 3786 7964 3792 8016
rect 3844 7964 3850 8016
rect 9416 8004 9444 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 15473 8075 15531 8081
rect 15473 8041 15485 8075
rect 15519 8072 15531 8075
rect 15746 8072 15752 8084
rect 15519 8044 15752 8072
rect 15519 8041 15531 8044
rect 15473 8035 15531 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19889 8075 19947 8081
rect 19889 8072 19901 8075
rect 19484 8044 19901 8072
rect 19484 8032 19490 8044
rect 19889 8041 19901 8044
rect 19935 8041 19947 8075
rect 19889 8035 19947 8041
rect 20990 8032 20996 8084
rect 21048 8032 21054 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 21876 8044 22131 8072
rect 21876 8032 21882 8044
rect 6840 7976 9444 8004
rect 6840 7945 6868 7976
rect 10502 7964 10508 8016
rect 10560 8004 10566 8016
rect 22103 8004 22131 8044
rect 22462 8032 22468 8084
rect 22520 8072 22526 8084
rect 22741 8075 22799 8081
rect 22741 8072 22753 8075
rect 22520 8044 22753 8072
rect 22520 8032 22526 8044
rect 22741 8041 22753 8044
rect 22787 8041 22799 8075
rect 22741 8035 22799 8041
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23474 8072 23480 8084
rect 23072 8044 23480 8072
rect 23072 8032 23078 8044
rect 23474 8032 23480 8044
rect 23532 8072 23538 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 23532 8044 24685 8072
rect 23532 8032 23538 8044
rect 24673 8041 24685 8044
rect 24719 8072 24731 8075
rect 24762 8072 24768 8084
rect 24719 8044 24768 8072
rect 24719 8041 24731 8044
rect 24673 8035 24731 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 25130 8032 25136 8084
rect 25188 8072 25194 8084
rect 25225 8075 25283 8081
rect 25225 8072 25237 8075
rect 25188 8044 25237 8072
rect 25188 8032 25194 8044
rect 25225 8041 25237 8044
rect 25271 8041 25283 8075
rect 25225 8035 25283 8041
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 28813 8075 28871 8081
rect 25924 8044 26004 8072
rect 25924 8032 25930 8044
rect 10560 7976 11100 8004
rect 10560 7964 10566 7976
rect 6825 7939 6883 7945
rect 4080 7908 4568 7936
rect 3512 7871 3570 7877
rect 3512 7837 3524 7871
rect 3558 7837 3570 7871
rect 3512 7831 3570 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 3694 7868 3700 7880
rect 3651 7840 3700 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3527 7800 3555 7831
rect 3694 7828 3700 7840
rect 3752 7868 3758 7880
rect 4080 7877 4108 7908
rect 4064 7871 4122 7877
rect 4064 7868 4076 7871
rect 3752 7840 4076 7868
rect 3752 7828 3758 7840
rect 4064 7837 4076 7840
rect 4110 7837 4122 7871
rect 4064 7831 4122 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4172 7800 4200 7831
rect 3527 7772 4200 7800
rect 3804 7744 3832 7772
rect 3786 7692 3792 7744
rect 3844 7692 3850 7744
rect 4540 7741 4568 7908
rect 6825 7905 6837 7939
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 7892 7908 8585 7936
rect 7892 7896 7898 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7936 10379 7939
rect 10962 7936 10968 7948
rect 10367 7908 10968 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11072 7945 11100 7976
rect 15488 7976 16160 8004
rect 15488 7948 15516 7976
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7905 11115 7939
rect 12115 7939 12173 7945
rect 12115 7936 12127 7939
rect 11057 7899 11115 7905
rect 11440 7908 12127 7936
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5316 7840 6101 7868
rect 5316 7828 5322 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 6236 7840 6285 7868
rect 6236 7828 6242 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6972 7840 7205 7868
rect 6972 7828 6978 7840
rect 7193 7837 7205 7840
rect 7239 7868 7251 7871
rect 7282 7868 7288 7880
rect 7239 7840 7288 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7282 7828 7288 7840
rect 7340 7868 7346 7880
rect 8662 7868 8668 7880
rect 7340 7840 8668 7868
rect 7340 7828 7346 7840
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10468 7840 10885 7868
rect 10468 7828 10474 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 7837 7803 7895 7809
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 8110 7800 8116 7812
rect 7883 7772 8116 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 10054 7803 10112 7809
rect 10054 7800 10066 7803
rect 8956 7772 10066 7800
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 6086 7732 6092 7744
rect 4571 7704 6092 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7732 7619 7735
rect 7650 7732 7656 7744
rect 7607 7704 7656 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 7745 7735 7803 7741
rect 7745 7701 7757 7735
rect 7791 7732 7803 7735
rect 8956 7732 8984 7772
rect 10054 7769 10066 7772
rect 10100 7769 10112 7803
rect 10054 7763 10112 7769
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11440 7800 11468 7908
rect 12115 7905 12127 7908
rect 12161 7905 12173 7939
rect 12115 7899 12173 7905
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 13814 7896 13820 7948
rect 13872 7896 13878 7948
rect 15470 7896 15476 7948
rect 15528 7896 15534 7948
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 16132 7945 16160 7976
rect 18064 7976 22048 8004
rect 18064 7948 18092 7976
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17678 7936 17684 7948
rect 17635 7908 17684 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18046 7936 18052 7948
rect 17911 7908 18052 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 18564 7908 19257 7936
rect 18564 7896 18570 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7868 13231 7871
rect 13998 7868 14004 7880
rect 13219 7840 14004 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 11112 7772 11468 7800
rect 11112 7760 11118 7772
rect 13004 7744 13032 7831
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14182 7868 14188 7880
rect 14139 7840 14188 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15252 7840 17071 7868
rect 15252 7828 15258 7840
rect 14360 7803 14418 7809
rect 14360 7769 14372 7803
rect 14406 7800 14418 7803
rect 15010 7800 15016 7812
rect 14406 7772 15016 7800
rect 14406 7769 14418 7772
rect 14360 7763 14418 7769
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 15979 7772 16344 7800
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 16316 7744 16344 7772
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 16761 7803 16819 7809
rect 16761 7800 16773 7803
rect 16724 7772 16773 7800
rect 16724 7760 16730 7772
rect 16761 7769 16773 7772
rect 16807 7800 16819 7803
rect 16942 7800 16948 7812
rect 16807 7772 16948 7800
rect 16807 7769 16819 7772
rect 16761 7763 16819 7769
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 17043 7800 17071 7840
rect 17954 7828 17960 7880
rect 18012 7868 18018 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 18012 7840 18153 7868
rect 18012 7828 18018 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 20714 7828 20720 7880
rect 20772 7828 20778 7880
rect 17043 7772 20760 7800
rect 7791 7704 8984 7732
rect 7791 7701 7803 7704
rect 7745 7695 7803 7701
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7732 11023 7735
rect 11333 7735 11391 7741
rect 11333 7732 11345 7735
rect 11011 7704 11345 7732
rect 11011 7701 11023 7704
rect 10965 7695 11023 7701
rect 11333 7701 11345 7704
rect 11379 7701 11391 7735
rect 11333 7695 11391 7701
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 13044 7704 13277 7732
rect 13044 7692 13050 7704
rect 13265 7701 13277 7704
rect 13311 7701 13323 7735
rect 13265 7695 13323 7701
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 15746 7732 15752 7744
rect 15611 7704 15752 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 18506 7692 18512 7744
rect 18564 7692 18570 7744
rect 20073 7735 20131 7741
rect 20073 7701 20085 7735
rect 20119 7732 20131 7735
rect 20162 7732 20168 7744
rect 20119 7704 20168 7732
rect 20119 7701 20131 7704
rect 20073 7695 20131 7701
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 20732 7732 20760 7772
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 20864 7772 20913 7800
rect 20864 7760 20870 7772
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 22020 7800 22048 7976
rect 22103 7976 24256 8004
rect 22103 7945 22131 7976
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7905 22155 7939
rect 24228 7936 24256 7976
rect 24854 7964 24860 8016
rect 24912 7964 24918 8016
rect 25976 8004 26004 8044
rect 28813 8041 28825 8075
rect 28859 8072 28871 8075
rect 28902 8072 28908 8084
rect 28859 8044 28908 8072
rect 28859 8041 28871 8044
rect 28813 8035 28871 8041
rect 28902 8032 28908 8044
rect 28960 8032 28966 8084
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 29825 8075 29883 8081
rect 29825 8072 29837 8075
rect 29696 8044 29837 8072
rect 29696 8032 29702 8044
rect 29825 8041 29837 8044
rect 29871 8041 29883 8075
rect 29825 8035 29883 8041
rect 30009 8075 30067 8081
rect 30009 8041 30021 8075
rect 30055 8072 30067 8075
rect 30650 8072 30656 8084
rect 30055 8044 30656 8072
rect 30055 8041 30067 8044
rect 30009 8035 30067 8041
rect 30650 8032 30656 8044
rect 30708 8032 30714 8084
rect 35434 8072 35440 8084
rect 31220 8044 35440 8072
rect 27157 8007 27215 8013
rect 27157 8004 27169 8007
rect 25976 7976 27169 8004
rect 27157 7973 27169 7976
rect 27203 8004 27215 8007
rect 30742 8004 30748 8016
rect 27203 7976 30748 8004
rect 27203 7973 27215 7976
rect 27157 7967 27215 7973
rect 25774 7936 25780 7948
rect 24228 7908 25780 7936
rect 22097 7899 22155 7905
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 25869 7939 25927 7945
rect 25869 7905 25881 7939
rect 25915 7936 25927 7939
rect 25958 7936 25964 7948
rect 25915 7908 25964 7936
rect 25915 7905 25927 7908
rect 25869 7899 25927 7905
rect 25958 7896 25964 7908
rect 26016 7896 26022 7948
rect 26142 7896 26148 7948
rect 26200 7936 26206 7948
rect 26200 7908 27927 7936
rect 26200 7896 26206 7908
rect 22370 7828 22376 7880
rect 22428 7828 22434 7880
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 25590 7828 25596 7880
rect 25648 7868 25654 7880
rect 26970 7868 26976 7880
rect 25648 7840 26976 7868
rect 25648 7828 25654 7840
rect 26970 7828 26976 7840
rect 27028 7828 27034 7880
rect 27899 7868 27927 7908
rect 27982 7896 27988 7948
rect 28040 7896 28046 7948
rect 28184 7945 28212 7976
rect 30742 7964 30748 7976
rect 30800 7964 30806 8016
rect 28169 7939 28227 7945
rect 28169 7905 28181 7939
rect 28215 7905 28227 7939
rect 28169 7899 28227 7905
rect 28353 7939 28411 7945
rect 28353 7905 28365 7939
rect 28399 7936 28411 7939
rect 28399 7908 28672 7936
rect 28399 7905 28411 7908
rect 28353 7899 28411 7905
rect 28534 7868 28540 7880
rect 27899 7840 28540 7868
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 28644 7812 28672 7908
rect 29638 7896 29644 7948
rect 29696 7936 29702 7948
rect 31220 7945 31248 8044
rect 35434 8032 35440 8044
rect 35492 8032 35498 8084
rect 36170 8032 36176 8084
rect 36228 8032 36234 8084
rect 36265 8075 36323 8081
rect 36265 8041 36277 8075
rect 36311 8072 36323 8075
rect 36354 8072 36360 8084
rect 36311 8044 36360 8072
rect 36311 8041 36323 8044
rect 36265 8035 36323 8041
rect 36354 8032 36360 8044
rect 36412 8032 36418 8084
rect 37737 8075 37795 8081
rect 37737 8041 37749 8075
rect 37783 8072 37795 8075
rect 39114 8072 39120 8084
rect 37783 8044 39120 8072
rect 37783 8041 37795 8044
rect 37737 8035 37795 8041
rect 39114 8032 39120 8044
rect 39172 8032 39178 8084
rect 44637 8075 44695 8081
rect 44637 8041 44649 8075
rect 44683 8041 44695 8075
rect 44637 8035 44695 8041
rect 33226 7964 33232 8016
rect 33284 7964 33290 8016
rect 43349 8007 43407 8013
rect 43349 7973 43361 8007
rect 43395 8004 43407 8007
rect 44652 8004 44680 8035
rect 44726 8032 44732 8084
rect 44784 8072 44790 8084
rect 45005 8075 45063 8081
rect 45005 8072 45017 8075
rect 44784 8044 45017 8072
rect 44784 8032 44790 8044
rect 45005 8041 45017 8044
rect 45051 8041 45063 8075
rect 49881 8075 49939 8081
rect 49881 8072 49893 8075
rect 45005 8035 45063 8041
rect 45572 8044 49893 8072
rect 45278 8004 45284 8016
rect 43395 7976 44036 8004
rect 44652 7976 45284 8004
rect 43395 7973 43407 7976
rect 43349 7967 43407 7973
rect 30561 7939 30619 7945
rect 30561 7936 30573 7939
rect 29696 7908 30573 7936
rect 29696 7896 29702 7908
rect 30561 7905 30573 7908
rect 30607 7936 30619 7939
rect 31205 7939 31263 7945
rect 31205 7936 31217 7939
rect 30607 7908 31217 7936
rect 30607 7905 30619 7908
rect 30561 7899 30619 7905
rect 31205 7905 31217 7908
rect 31251 7905 31263 7939
rect 31205 7899 31263 7905
rect 31754 7896 31760 7948
rect 31812 7936 31818 7948
rect 32306 7936 32312 7948
rect 31812 7908 32312 7936
rect 31812 7896 31818 7908
rect 32306 7896 32312 7908
rect 32364 7896 32370 7948
rect 33244 7936 33272 7964
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 33244 7908 33425 7936
rect 33413 7905 33425 7908
rect 33459 7905 33471 7939
rect 33413 7899 33471 7905
rect 42978 7896 42984 7948
rect 43036 7896 43042 7948
rect 44008 7945 44036 7976
rect 45278 7964 45284 7976
rect 45336 7964 45342 8016
rect 45572 7945 45600 8044
rect 49881 8041 49893 8044
rect 49927 8041 49939 8075
rect 49881 8035 49939 8041
rect 50157 8075 50215 8081
rect 50157 8041 50169 8075
rect 50203 8072 50215 8075
rect 50430 8072 50436 8084
rect 50203 8044 50436 8072
rect 50203 8041 50215 8044
rect 50157 8035 50215 8041
rect 47305 8007 47363 8013
rect 47305 7973 47317 8007
rect 47351 8004 47363 8007
rect 47670 8004 47676 8016
rect 47351 7976 47676 8004
rect 47351 7973 47363 7976
rect 47305 7967 47363 7973
rect 47670 7964 47676 7976
rect 47728 8004 47734 8016
rect 49053 8007 49111 8013
rect 49053 8004 49065 8007
rect 47728 7976 49065 8004
rect 47728 7964 47734 7976
rect 49053 7973 49065 7976
rect 49099 8004 49111 8007
rect 49786 8004 49792 8016
rect 49099 7976 49792 8004
rect 49099 7973 49111 7976
rect 49053 7967 49111 7973
rect 49786 7964 49792 7976
rect 49844 7964 49850 8016
rect 43993 7939 44051 7945
rect 43993 7905 44005 7939
rect 44039 7905 44051 7939
rect 45557 7939 45615 7945
rect 45557 7936 45569 7939
rect 43993 7899 44051 7905
rect 44652 7908 45569 7936
rect 30466 7828 30472 7880
rect 30524 7868 30530 7880
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 30524 7840 30849 7868
rect 30524 7828 30530 7840
rect 30837 7837 30849 7840
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 31148 7840 31708 7868
rect 23109 7803 23167 7809
rect 23109 7800 23121 7803
rect 22020 7772 23121 7800
rect 20901 7763 20959 7769
rect 23109 7769 23121 7772
rect 23155 7800 23167 7803
rect 23934 7800 23940 7812
rect 23155 7772 23940 7800
rect 23155 7769 23167 7772
rect 23109 7763 23167 7769
rect 23934 7760 23940 7772
rect 23992 7760 23998 7812
rect 25038 7760 25044 7812
rect 25096 7760 25102 7812
rect 26418 7800 26424 7812
rect 26252 7772 26424 7800
rect 22002 7732 22008 7744
rect 20732 7704 22008 7732
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 23198 7692 23204 7744
rect 23256 7732 23262 7744
rect 23293 7735 23351 7741
rect 23293 7732 23305 7735
rect 23256 7704 23305 7732
rect 23256 7692 23262 7704
rect 23293 7701 23305 7704
rect 23339 7701 23351 7735
rect 23293 7695 23351 7701
rect 25685 7735 25743 7741
rect 25685 7701 25697 7735
rect 25731 7732 25743 7735
rect 26252 7732 26280 7772
rect 26418 7760 26424 7772
rect 26476 7760 26482 7812
rect 27341 7803 27399 7809
rect 27341 7800 27353 7803
rect 26620 7772 27353 7800
rect 26620 7744 26648 7772
rect 27341 7769 27353 7772
rect 27387 7800 27399 7803
rect 28445 7803 28503 7809
rect 28445 7800 28457 7803
rect 27387 7772 28457 7800
rect 27387 7769 27399 7772
rect 27341 7763 27399 7769
rect 28445 7769 28457 7772
rect 28491 7769 28503 7803
rect 28445 7763 28503 7769
rect 28626 7760 28632 7812
rect 28684 7760 28690 7812
rect 30377 7803 30435 7809
rect 30377 7769 30389 7803
rect 30423 7800 30435 7803
rect 30926 7800 30932 7812
rect 30423 7772 30932 7800
rect 30423 7769 30435 7772
rect 30377 7763 30435 7769
rect 30926 7760 30932 7772
rect 30984 7800 30990 7812
rect 31148 7800 31176 7840
rect 30984 7772 31176 7800
rect 31680 7800 31708 7840
rect 31938 7828 31944 7880
rect 31996 7828 32002 7880
rect 33045 7871 33103 7877
rect 33045 7837 33057 7871
rect 33091 7868 33103 7871
rect 34333 7871 34391 7877
rect 34333 7868 34345 7871
rect 33091 7840 34345 7868
rect 33091 7837 33103 7840
rect 33045 7831 33103 7837
rect 34333 7837 34345 7840
rect 34379 7837 34391 7871
rect 34333 7831 34391 7837
rect 34793 7871 34851 7877
rect 34793 7837 34805 7871
rect 34839 7868 34851 7871
rect 34882 7868 34888 7880
rect 34839 7840 34888 7868
rect 34839 7837 34851 7840
rect 34793 7831 34851 7837
rect 32306 7800 32312 7812
rect 31680 7772 32312 7800
rect 30984 7760 30990 7772
rect 32306 7760 32312 7772
rect 32364 7760 32370 7812
rect 25731 7704 26280 7732
rect 25731 7701 25743 7704
rect 25685 7695 25743 7701
rect 26326 7692 26332 7744
rect 26384 7692 26390 7744
rect 26602 7692 26608 7744
rect 26660 7692 26666 7744
rect 26786 7692 26792 7744
rect 26844 7692 26850 7744
rect 26878 7692 26884 7744
rect 26936 7732 26942 7744
rect 30098 7732 30104 7744
rect 26936 7704 30104 7732
rect 26936 7692 26942 7704
rect 30098 7692 30104 7704
rect 30156 7692 30162 7744
rect 30469 7735 30527 7741
rect 30469 7701 30481 7735
rect 30515 7732 30527 7735
rect 30558 7732 30564 7744
rect 30515 7704 30564 7732
rect 30515 7701 30527 7704
rect 30469 7695 30527 7701
rect 30558 7692 30564 7704
rect 30616 7692 30622 7744
rect 30742 7692 30748 7744
rect 30800 7732 30806 7744
rect 33060 7732 33088 7831
rect 34882 7828 34888 7840
rect 34940 7868 34946 7880
rect 37645 7871 37703 7877
rect 37645 7868 37657 7871
rect 34940 7840 37657 7868
rect 34940 7828 34946 7840
rect 37645 7837 37657 7840
rect 37691 7868 37703 7871
rect 39114 7868 39120 7880
rect 37691 7840 39120 7868
rect 37691 7837 37703 7840
rect 37645 7831 37703 7837
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39298 7828 39304 7880
rect 39356 7828 39362 7880
rect 41046 7828 41052 7880
rect 41104 7828 41110 7880
rect 41233 7871 41291 7877
rect 41233 7837 41245 7871
rect 41279 7837 41291 7871
rect 41233 7831 41291 7837
rect 35060 7803 35118 7809
rect 35060 7769 35072 7803
rect 35106 7800 35118 7803
rect 35250 7800 35256 7812
rect 35106 7772 35256 7800
rect 35106 7769 35118 7772
rect 35060 7763 35118 7769
rect 35250 7760 35256 7772
rect 35308 7760 35314 7812
rect 36354 7760 36360 7812
rect 36412 7800 36418 7812
rect 36538 7800 36544 7812
rect 36412 7772 36544 7800
rect 36412 7760 36418 7772
rect 36538 7760 36544 7772
rect 36596 7760 36602 7812
rect 37400 7803 37458 7809
rect 37400 7769 37412 7803
rect 37446 7800 37458 7803
rect 37826 7800 37832 7812
rect 37446 7772 37832 7800
rect 37446 7769 37458 7772
rect 37400 7763 37458 7769
rect 37826 7760 37832 7772
rect 37884 7760 37890 7812
rect 38872 7803 38930 7809
rect 38872 7769 38884 7803
rect 38918 7800 38930 7803
rect 39316 7800 39344 7828
rect 38918 7772 39344 7800
rect 38918 7769 38930 7772
rect 38872 7763 38930 7769
rect 40954 7760 40960 7812
rect 41012 7800 41018 7812
rect 41248 7800 41276 7831
rect 41506 7828 41512 7880
rect 41564 7868 41570 7880
rect 41969 7871 42027 7877
rect 41969 7868 41981 7871
rect 41564 7840 41981 7868
rect 41564 7828 41570 7840
rect 41969 7837 41981 7840
rect 42015 7868 42027 7871
rect 42996 7868 43024 7896
rect 42015 7840 43024 7868
rect 42015 7837 42027 7840
rect 41969 7831 42027 7837
rect 41012 7772 41276 7800
rect 42236 7803 42294 7809
rect 41012 7760 41018 7772
rect 42236 7769 42248 7803
rect 42282 7800 42294 7803
rect 42426 7800 42432 7812
rect 42282 7772 42432 7800
rect 42282 7769 42294 7772
rect 42236 7763 42294 7769
rect 42426 7760 42432 7772
rect 42484 7760 42490 7812
rect 44652 7744 44680 7908
rect 45557 7905 45569 7908
rect 45603 7905 45615 7939
rect 45557 7899 45615 7905
rect 47762 7896 47768 7948
rect 47820 7896 47826 7948
rect 48593 7939 48651 7945
rect 48593 7905 48605 7939
rect 48639 7905 48651 7939
rect 49896 7936 49924 8035
rect 50430 8032 50436 8044
rect 50488 8032 50494 8084
rect 51074 8032 51080 8084
rect 51132 8072 51138 8084
rect 51350 8072 51356 8084
rect 51132 8044 51356 8072
rect 51132 8032 51138 8044
rect 51350 8032 51356 8044
rect 51408 8072 51414 8084
rect 51721 8075 51779 8081
rect 51721 8072 51733 8075
rect 51408 8044 51733 8072
rect 51408 8032 51414 8044
rect 51721 8041 51733 8044
rect 51767 8041 51779 8075
rect 57793 8075 57851 8081
rect 51721 8035 51779 8041
rect 53668 8044 57376 8072
rect 50709 7939 50767 7945
rect 50709 7936 50721 7939
rect 49896 7908 50721 7936
rect 48593 7899 48651 7905
rect 50709 7905 50721 7908
rect 50755 7936 50767 7939
rect 50755 7908 52224 7936
rect 50755 7905 50767 7908
rect 50709 7899 50767 7905
rect 45370 7828 45376 7880
rect 45428 7828 45434 7880
rect 46750 7828 46756 7880
rect 46808 7828 46814 7880
rect 46842 7828 46848 7880
rect 46900 7877 46906 7880
rect 46900 7871 46949 7877
rect 46900 7837 46903 7871
rect 46937 7837 46949 7871
rect 46900 7831 46949 7837
rect 46900 7828 46906 7831
rect 47026 7828 47032 7880
rect 47084 7828 47090 7880
rect 47946 7828 47952 7880
rect 48004 7828 48010 7880
rect 48406 7828 48412 7880
rect 48464 7828 48470 7880
rect 44729 7803 44787 7809
rect 44729 7769 44741 7803
rect 44775 7800 44787 7803
rect 45830 7800 45836 7812
rect 44775 7772 45836 7800
rect 44775 7769 44787 7772
rect 44729 7763 44787 7769
rect 45830 7760 45836 7772
rect 45888 7760 45894 7812
rect 48501 7803 48559 7809
rect 48501 7800 48513 7803
rect 47780 7772 48513 7800
rect 30800 7704 33088 7732
rect 30800 7692 30806 7704
rect 36170 7692 36176 7744
rect 36228 7732 36234 7744
rect 38746 7732 38752 7744
rect 36228 7704 38752 7732
rect 36228 7692 36234 7704
rect 38746 7692 38752 7704
rect 38804 7692 38810 7744
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 40494 7692 40500 7744
rect 40552 7692 40558 7744
rect 41782 7692 41788 7744
rect 41840 7732 41846 7744
rect 41877 7735 41935 7741
rect 41877 7732 41889 7735
rect 41840 7704 41889 7732
rect 41840 7692 41846 7704
rect 41877 7701 41889 7704
rect 41923 7732 41935 7735
rect 42334 7732 42340 7744
rect 41923 7704 42340 7732
rect 41923 7701 41935 7704
rect 41877 7695 41935 7701
rect 42334 7692 42340 7704
rect 42392 7692 42398 7744
rect 42978 7692 42984 7744
rect 43036 7732 43042 7744
rect 43441 7735 43499 7741
rect 43441 7732 43453 7735
rect 43036 7704 43453 7732
rect 43036 7692 43042 7704
rect 43441 7701 43453 7704
rect 43487 7701 43499 7735
rect 43441 7695 43499 7701
rect 44453 7735 44511 7741
rect 44453 7701 44465 7735
rect 44499 7732 44511 7735
rect 44634 7732 44640 7744
rect 44499 7704 44640 7732
rect 44499 7701 44511 7704
rect 44453 7695 44511 7701
rect 44634 7692 44640 7704
rect 44692 7692 44698 7744
rect 45465 7735 45523 7741
rect 45465 7701 45477 7735
rect 45511 7732 45523 7735
rect 45554 7732 45560 7744
rect 45511 7704 45560 7732
rect 45511 7701 45523 7704
rect 45465 7695 45523 7701
rect 45554 7692 45560 7704
rect 45612 7692 45618 7744
rect 46109 7735 46167 7741
rect 46109 7701 46121 7735
rect 46155 7732 46167 7735
rect 47780 7732 47808 7772
rect 48501 7769 48513 7772
rect 48547 7769 48559 7803
rect 48501 7763 48559 7769
rect 48608 7744 48636 7899
rect 50982 7828 50988 7880
rect 51040 7828 51046 7880
rect 50525 7803 50583 7809
rect 50525 7769 50537 7803
rect 50571 7800 50583 7803
rect 51350 7800 51356 7812
rect 50571 7772 51356 7800
rect 50571 7769 50583 7772
rect 50525 7763 50583 7769
rect 51350 7760 51356 7772
rect 51408 7800 51414 7812
rect 51629 7803 51687 7809
rect 51629 7800 51641 7803
rect 51408 7772 51641 7800
rect 51408 7760 51414 7772
rect 51629 7769 51641 7772
rect 51675 7769 51687 7803
rect 52196 7800 52224 7908
rect 52270 7896 52276 7948
rect 52328 7896 52334 7948
rect 52638 7896 52644 7948
rect 52696 7936 52702 7948
rect 52696 7908 52960 7936
rect 52696 7896 52702 7908
rect 52822 7828 52828 7880
rect 52880 7828 52886 7880
rect 52932 7868 52960 7908
rect 53668 7868 53696 8044
rect 53745 7939 53803 7945
rect 53745 7905 53757 7939
rect 53791 7905 53803 7939
rect 57348 7936 57376 8044
rect 57793 8041 57805 8075
rect 57839 8072 57851 8075
rect 57882 8072 57888 8084
rect 57839 8044 57888 8072
rect 57839 8041 57851 8044
rect 57793 8035 57851 8041
rect 57882 8032 57888 8044
rect 57940 8032 57946 8084
rect 58434 8032 58440 8084
rect 58492 8032 58498 8084
rect 57701 8007 57759 8013
rect 57701 7973 57713 8007
rect 57747 8004 57759 8007
rect 58452 8004 58480 8032
rect 57747 7976 58480 8004
rect 57747 7973 57759 7976
rect 57701 7967 57759 7973
rect 57882 7936 57888 7948
rect 57348 7908 57888 7936
rect 53745 7899 53803 7905
rect 52932 7840 53696 7868
rect 53760 7868 53788 7899
rect 57882 7896 57888 7908
rect 57940 7936 57946 7948
rect 58345 7939 58403 7945
rect 58345 7936 58357 7939
rect 57940 7908 58357 7936
rect 57940 7896 57946 7908
rect 58345 7905 58357 7908
rect 58391 7905 58403 7939
rect 58345 7899 58403 7905
rect 54294 7868 54300 7880
rect 53760 7840 54300 7868
rect 54294 7828 54300 7840
rect 54352 7828 54358 7880
rect 55861 7871 55919 7877
rect 55861 7868 55873 7871
rect 54956 7840 55873 7868
rect 53742 7800 53748 7812
rect 52196 7772 53748 7800
rect 51629 7763 51687 7769
rect 53742 7760 53748 7772
rect 53800 7760 53806 7812
rect 54012 7803 54070 7809
rect 54012 7769 54024 7803
rect 54058 7800 54070 7803
rect 54202 7800 54208 7812
rect 54058 7772 54208 7800
rect 54058 7769 54070 7772
rect 54012 7763 54070 7769
rect 54202 7760 54208 7772
rect 54260 7760 54266 7812
rect 46155 7704 47808 7732
rect 46155 7701 46167 7704
rect 46109 7695 46167 7701
rect 48038 7692 48044 7744
rect 48096 7692 48102 7744
rect 48590 7692 48596 7744
rect 48648 7692 48654 7744
rect 50614 7692 50620 7744
rect 50672 7692 50678 7744
rect 52730 7692 52736 7744
rect 52788 7692 52794 7744
rect 53193 7735 53251 7741
rect 53193 7701 53205 7735
rect 53239 7732 53251 7735
rect 54956 7732 54984 7840
rect 55861 7837 55873 7840
rect 55907 7837 55919 7871
rect 55861 7831 55919 7837
rect 56226 7828 56232 7880
rect 56284 7868 56290 7880
rect 56594 7877 56600 7880
rect 56321 7871 56379 7877
rect 56321 7868 56333 7871
rect 56284 7840 56333 7868
rect 56284 7828 56290 7840
rect 56321 7837 56333 7840
rect 56367 7837 56379 7871
rect 56588 7868 56600 7877
rect 56555 7840 56600 7868
rect 56321 7831 56379 7837
rect 56588 7831 56600 7840
rect 56594 7828 56600 7831
rect 56652 7828 56658 7880
rect 58158 7828 58164 7880
rect 58216 7828 58222 7880
rect 55030 7760 55036 7812
rect 55088 7800 55094 7812
rect 55309 7803 55367 7809
rect 55309 7800 55321 7803
rect 55088 7772 55321 7800
rect 55088 7760 55094 7772
rect 55309 7769 55321 7772
rect 55355 7769 55367 7803
rect 55309 7763 55367 7769
rect 53239 7704 54984 7732
rect 53239 7701 53251 7704
rect 53193 7695 53251 7701
rect 55122 7692 55128 7744
rect 55180 7692 55186 7744
rect 57054 7692 57060 7744
rect 57112 7732 57118 7744
rect 58253 7735 58311 7741
rect 58253 7732 58265 7735
rect 57112 7704 58265 7732
rect 57112 7692 57118 7704
rect 58253 7701 58265 7704
rect 58299 7701 58311 7735
rect 58253 7695 58311 7701
rect 1104 7642 59040 7664
rect 1104 7590 15394 7642
rect 15446 7590 15458 7642
rect 15510 7590 15522 7642
rect 15574 7590 15586 7642
rect 15638 7590 15650 7642
rect 15702 7590 29838 7642
rect 29890 7590 29902 7642
rect 29954 7590 29966 7642
rect 30018 7590 30030 7642
rect 30082 7590 30094 7642
rect 30146 7590 44282 7642
rect 44334 7590 44346 7642
rect 44398 7590 44410 7642
rect 44462 7590 44474 7642
rect 44526 7590 44538 7642
rect 44590 7590 58726 7642
rect 58778 7590 58790 7642
rect 58842 7590 58854 7642
rect 58906 7590 58918 7642
rect 58970 7590 58982 7642
rect 59034 7590 59040 7642
rect 1104 7568 59040 7590
rect 3694 7488 3700 7540
rect 3752 7488 3758 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6362 7528 6368 7540
rect 6043 7500 6368 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 7616 7500 7941 7528
rect 7616 7488 7622 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9398 7528 9404 7540
rect 9079 7500 9404 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 9950 7528 9956 7540
rect 9824 7500 9956 7528
rect 9824 7488 9830 7500
rect 9950 7488 9956 7500
rect 10008 7528 10014 7540
rect 10008 7500 11192 7528
rect 10008 7488 10014 7500
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7429 5319 7463
rect 5261 7423 5319 7429
rect 7193 7463 7251 7469
rect 7193 7429 7205 7463
rect 7239 7460 7251 7463
rect 7239 7432 8156 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 5276 7392 5304 7423
rect 8128 7404 8156 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 10560 7432 11100 7460
rect 10560 7420 10566 7432
rect 5442 7392 5448 7404
rect 5276 7364 5448 7392
rect 5442 7352 5448 7364
rect 5500 7392 5506 7404
rect 7282 7392 7288 7404
rect 5500 7364 7288 7392
rect 5500 7352 5506 7364
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7432 7364 7481 7392
rect 7432 7352 7438 7364
rect 7469 7361 7481 7364
rect 7515 7392 7527 7395
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 7515 7364 7573 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 7834 7392 7840 7404
rect 7791 7364 7840 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5592 7296 5733 7324
rect 5592 7284 5598 7296
rect 5721 7293 5733 7296
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7760 7324 7788 7355
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8168 7364 8892 7392
rect 8168 7352 8174 7364
rect 6871 7296 7788 7324
rect 8205 7327 8263 7333
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 8754 7324 8760 7336
rect 8251 7296 8760 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 8864 7324 8892 7364
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 11072 7401 11100 7432
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 10413 7327 10471 7333
rect 8864 7296 9536 7324
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 5261 7259 5319 7265
rect 5261 7256 5273 7259
rect 3844 7228 5273 7256
rect 3844 7216 3850 7228
rect 5261 7225 5273 7228
rect 5307 7225 5319 7259
rect 5261 7219 5319 7225
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 9401 7259 9459 7265
rect 9401 7256 9413 7259
rect 7708 7228 9413 7256
rect 7708 7216 7714 7228
rect 9401 7225 9413 7228
rect 9447 7225 9459 7259
rect 9508 7256 9536 7296
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 10870 7324 10876 7336
rect 10459 7296 10876 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11164 7256 11192 7500
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11296 7500 11805 7528
rect 11296 7488 11302 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 12345 7531 12403 7537
rect 12345 7497 12357 7531
rect 12391 7528 12403 7531
rect 12986 7528 12992 7540
rect 12391 7500 12992 7528
rect 12391 7497 12403 7500
rect 12345 7491 12403 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 14056 7500 14197 7528
rect 14056 7488 14062 7500
rect 14185 7497 14197 7500
rect 14231 7528 14243 7531
rect 14550 7528 14556 7540
rect 14231 7500 14556 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 15010 7488 15016 7540
rect 15068 7488 15074 7540
rect 15746 7488 15752 7540
rect 15804 7488 15810 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 15988 7500 16313 7528
rect 15988 7488 15994 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 18932 7500 19334 7528
rect 18932 7488 18938 7500
rect 12526 7420 12532 7472
rect 12584 7420 12590 7472
rect 12802 7420 12808 7472
rect 12860 7420 12866 7472
rect 12544 7392 12572 7420
rect 15378 7392 15384 7404
rect 12084 7364 12434 7392
rect 12084 7336 12112 7364
rect 12406 7336 12434 7364
rect 12544 7364 15384 7392
rect 12066 7284 12072 7336
rect 12124 7284 12130 7336
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12253 7327 12311 7333
rect 12253 7324 12265 7327
rect 12216 7296 12265 7324
rect 12216 7284 12222 7296
rect 12253 7293 12265 7296
rect 12299 7293 12311 7327
rect 12406 7296 12440 7336
rect 12253 7287 12311 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12544 7256 12572 7364
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 15764 7392 15792 7488
rect 15703 7364 15792 7392
rect 16393 7395 16451 7401
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 16393 7361 16405 7395
rect 16439 7392 16451 7395
rect 16942 7392 16948 7404
rect 16439 7364 16948 7392
rect 16439 7361 16451 7364
rect 16393 7355 16451 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 18069 7395 18127 7401
rect 18069 7361 18081 7395
rect 18115 7392 18127 7395
rect 18230 7392 18236 7404
rect 18115 7364 18236 7392
rect 18115 7361 18127 7364
rect 18069 7355 18127 7361
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 19306 7392 19334 7500
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 21910 7528 21916 7540
rect 20220 7500 21916 7528
rect 20220 7488 20226 7500
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 23201 7531 23259 7537
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 23842 7528 23848 7540
rect 23247 7500 23848 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 24949 7531 25007 7537
rect 24949 7497 24961 7531
rect 24995 7528 25007 7531
rect 25590 7528 25596 7540
rect 24995 7500 25596 7528
rect 24995 7497 25007 7500
rect 24949 7491 25007 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 26418 7488 26424 7540
rect 26476 7528 26482 7540
rect 31205 7531 31263 7537
rect 26476 7500 29776 7528
rect 26476 7488 26482 7500
rect 20257 7463 20315 7469
rect 20257 7429 20269 7463
rect 20303 7460 20315 7463
rect 20530 7460 20536 7472
rect 20303 7432 20536 7460
rect 20303 7429 20315 7432
rect 20257 7423 20315 7429
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 24670 7460 24676 7472
rect 21836 7432 24676 7460
rect 19306 7364 20392 7392
rect 20364 7336 20392 7364
rect 21266 7352 21272 7404
rect 21324 7392 21330 7404
rect 21836 7401 21864 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 26786 7420 26792 7472
rect 26844 7460 26850 7472
rect 26844 7432 27660 7460
rect 26844 7420 26850 7432
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21324 7364 21833 7392
rect 21324 7352 21330 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 22077 7395 22135 7401
rect 22077 7392 22089 7395
rect 21821 7355 21879 7361
rect 21928 7364 22089 7392
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 9508 7228 10640 7256
rect 11164 7228 12572 7256
rect 12713 7259 12771 7265
rect 9401 7219 9459 7225
rect 7469 7191 7527 7197
rect 7469 7157 7481 7191
rect 7515 7188 7527 7191
rect 8846 7188 8852 7200
rect 7515 7160 8852 7188
rect 7515 7157 7527 7160
rect 7469 7151 7527 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 10502 7148 10508 7200
rect 10560 7148 10566 7200
rect 10612 7188 10640 7228
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 13372 7256 13400 7287
rect 13538 7284 13544 7336
rect 13596 7284 13602 7336
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15286 7324 15292 7336
rect 14967 7296 15292 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 18322 7284 18328 7336
rect 18380 7284 18386 7336
rect 19705 7327 19763 7333
rect 19705 7293 19717 7327
rect 19751 7324 19763 7327
rect 19751 7296 19840 7324
rect 19751 7293 19763 7296
rect 19705 7287 19763 7293
rect 19812 7265 19840 7296
rect 20346 7284 20352 7336
rect 20404 7284 20410 7336
rect 21085 7327 21143 7333
rect 21085 7293 21097 7327
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21637 7327 21695 7333
rect 21637 7293 21649 7327
rect 21683 7324 21695 7327
rect 21928 7324 21956 7364
rect 22077 7361 22089 7364
rect 22123 7361 22135 7395
rect 22077 7355 22135 7361
rect 23658 7352 23664 7404
rect 23716 7352 23722 7404
rect 24946 7352 24952 7404
rect 25004 7392 25010 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 25004 7364 25053 7392
rect 25004 7352 25010 7364
rect 25041 7361 25053 7364
rect 25087 7392 25099 7395
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 25087 7364 27169 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 27157 7361 27169 7364
rect 27203 7392 27215 7395
rect 27522 7392 27528 7404
rect 27203 7364 27528 7392
rect 27203 7361 27215 7364
rect 27157 7355 27215 7361
rect 27522 7352 27528 7364
rect 27580 7352 27586 7404
rect 27632 7392 27660 7432
rect 27899 7432 29684 7460
rect 27899 7392 27927 7432
rect 27632 7364 27927 7392
rect 27982 7352 27988 7404
rect 28040 7352 28046 7404
rect 28718 7352 28724 7404
rect 28776 7401 28782 7404
rect 29656 7401 29684 7432
rect 28776 7392 28788 7401
rect 29641 7395 29699 7401
rect 28776 7364 28821 7392
rect 28776 7355 28788 7364
rect 29641 7361 29653 7395
rect 29687 7361 29699 7395
rect 29748 7392 29776 7500
rect 31205 7497 31217 7531
rect 31251 7528 31263 7531
rect 31386 7528 31392 7540
rect 31251 7500 31392 7528
rect 31251 7497 31263 7500
rect 31205 7491 31263 7497
rect 31386 7488 31392 7500
rect 31444 7488 31450 7540
rect 36262 7488 36268 7540
rect 36320 7488 36326 7540
rect 36354 7488 36360 7540
rect 36412 7488 36418 7540
rect 36449 7531 36507 7537
rect 36449 7497 36461 7531
rect 36495 7528 36507 7531
rect 37918 7528 37924 7540
rect 36495 7500 37924 7528
rect 36495 7497 36507 7500
rect 36449 7491 36507 7497
rect 37918 7488 37924 7500
rect 37976 7488 37982 7540
rect 39114 7488 39120 7540
rect 39172 7488 39178 7540
rect 40494 7488 40500 7540
rect 40552 7488 40558 7540
rect 40954 7488 40960 7540
rect 41012 7488 41018 7540
rect 41046 7488 41052 7540
rect 41104 7488 41110 7540
rect 41414 7488 41420 7540
rect 41472 7528 41478 7540
rect 41509 7531 41567 7537
rect 41509 7528 41521 7531
rect 41472 7500 41521 7528
rect 41472 7488 41478 7500
rect 41509 7497 41521 7500
rect 41555 7528 41567 7531
rect 42705 7531 42763 7537
rect 42705 7528 42717 7531
rect 41555 7500 42717 7528
rect 41555 7497 41567 7500
rect 41509 7491 41567 7497
rect 42705 7497 42717 7500
rect 42751 7497 42763 7531
rect 42705 7491 42763 7497
rect 42797 7531 42855 7537
rect 42797 7497 42809 7531
rect 42843 7528 42855 7531
rect 42978 7528 42984 7540
rect 42843 7500 42984 7528
rect 42843 7497 42855 7500
rect 42797 7491 42855 7497
rect 42978 7488 42984 7500
rect 43036 7488 43042 7540
rect 43070 7488 43076 7540
rect 43128 7528 43134 7540
rect 43165 7531 43223 7537
rect 43165 7528 43177 7531
rect 43128 7500 43177 7528
rect 43128 7488 43134 7500
rect 43165 7497 43177 7500
rect 43211 7497 43223 7531
rect 43165 7491 43223 7497
rect 45646 7488 45652 7540
rect 45704 7488 45710 7540
rect 45830 7488 45836 7540
rect 45888 7528 45894 7540
rect 47210 7528 47216 7540
rect 45888 7500 47216 7528
rect 45888 7488 45894 7500
rect 47210 7488 47216 7500
rect 47268 7488 47274 7540
rect 47854 7488 47860 7540
rect 47912 7528 47918 7540
rect 48317 7531 48375 7537
rect 48317 7528 48329 7531
rect 47912 7500 48329 7528
rect 47912 7488 47918 7500
rect 48317 7497 48329 7500
rect 48363 7497 48375 7531
rect 48317 7491 48375 7497
rect 50617 7531 50675 7537
rect 50617 7497 50629 7531
rect 50663 7528 50675 7531
rect 50982 7528 50988 7540
rect 50663 7500 50988 7528
rect 50663 7497 50675 7500
rect 50617 7491 50675 7497
rect 50982 7488 50988 7500
rect 51040 7488 51046 7540
rect 51994 7488 52000 7540
rect 52052 7528 52058 7540
rect 52181 7531 52239 7537
rect 52181 7528 52193 7531
rect 52052 7500 52193 7528
rect 52052 7488 52058 7500
rect 52181 7497 52193 7500
rect 52227 7497 52239 7531
rect 52181 7491 52239 7497
rect 52733 7531 52791 7537
rect 52733 7497 52745 7531
rect 52779 7528 52791 7531
rect 53374 7528 53380 7540
rect 52779 7500 53380 7528
rect 52779 7497 52791 7500
rect 52733 7491 52791 7497
rect 53374 7488 53380 7500
rect 53432 7488 53438 7540
rect 54294 7528 54300 7540
rect 54128 7500 54300 7528
rect 30092 7463 30150 7469
rect 30092 7429 30104 7463
rect 30138 7460 30150 7463
rect 30282 7460 30288 7472
rect 30138 7432 30288 7460
rect 30138 7429 30150 7432
rect 30092 7423 30150 7429
rect 30282 7420 30288 7432
rect 30340 7420 30346 7472
rect 36280 7460 36308 7488
rect 38013 7463 38071 7469
rect 38013 7460 38025 7463
rect 32048 7432 34928 7460
rect 36280 7432 38025 7460
rect 32048 7392 32076 7432
rect 29748 7364 32076 7392
rect 32125 7395 32183 7401
rect 29641 7355 29699 7361
rect 32125 7361 32137 7395
rect 32171 7392 32183 7395
rect 32214 7392 32220 7404
rect 32171 7364 32220 7392
rect 32171 7361 32183 7364
rect 32125 7355 32183 7361
rect 28776 7352 28782 7355
rect 32214 7352 32220 7364
rect 32272 7352 32278 7404
rect 32392 7395 32450 7401
rect 32392 7361 32404 7395
rect 32438 7392 32450 7395
rect 32438 7364 33548 7392
rect 32438 7361 32450 7364
rect 32392 7355 32450 7361
rect 21683 7296 21956 7324
rect 21683 7293 21695 7296
rect 21637 7287 21695 7293
rect 19797 7259 19855 7265
rect 12759 7228 13400 7256
rect 14200 7228 16712 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 14200 7188 14228 7228
rect 16684 7200 16712 7228
rect 18800 7228 19472 7256
rect 10612 7160 14228 7188
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 16666 7148 16672 7200
rect 16724 7148 16730 7200
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 17402 7188 17408 7200
rect 16991 7160 17408 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 18800 7188 18828 7228
rect 17736 7160 18828 7188
rect 19061 7191 19119 7197
rect 17736 7148 17742 7160
rect 19061 7157 19073 7191
rect 19107 7188 19119 7191
rect 19334 7188 19340 7200
rect 19107 7160 19340 7188
rect 19107 7157 19119 7160
rect 19061 7151 19119 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19444 7188 19472 7228
rect 19797 7225 19809 7259
rect 19843 7225 19855 7259
rect 19797 7219 19855 7225
rect 20809 7191 20867 7197
rect 20809 7188 20821 7191
rect 19444 7160 20821 7188
rect 20809 7157 20821 7160
rect 20855 7188 20867 7191
rect 20990 7188 20996 7200
rect 20855 7160 20996 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21100 7188 21128 7287
rect 23014 7284 23020 7336
rect 23072 7324 23078 7336
rect 23753 7327 23811 7333
rect 23753 7324 23765 7327
rect 23072 7296 23765 7324
rect 23072 7284 23078 7296
rect 23753 7293 23765 7296
rect 23799 7293 23811 7327
rect 23753 7287 23811 7293
rect 23934 7284 23940 7336
rect 23992 7284 23998 7336
rect 24394 7284 24400 7336
rect 24452 7284 24458 7336
rect 27617 7259 27675 7265
rect 27617 7225 27629 7259
rect 27663 7256 27675 7259
rect 28000 7256 28028 7352
rect 28997 7327 29055 7333
rect 28997 7293 29009 7327
rect 29043 7324 29055 7327
rect 29825 7327 29883 7333
rect 29825 7324 29837 7327
rect 29043 7296 29837 7324
rect 29043 7293 29055 7296
rect 28997 7287 29055 7293
rect 29825 7293 29837 7296
rect 29871 7293 29883 7327
rect 29825 7287 29883 7293
rect 27663 7228 28028 7256
rect 27663 7225 27675 7228
rect 27617 7219 27675 7225
rect 22462 7188 22468 7200
rect 21100 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 23290 7148 23296 7200
rect 23348 7148 23354 7200
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 25924 7160 26341 7188
rect 25924 7148 25930 7160
rect 26329 7157 26341 7160
rect 26375 7188 26387 7191
rect 29012 7188 29040 7287
rect 31846 7284 31852 7336
rect 31904 7284 31910 7336
rect 33520 7324 33548 7364
rect 33594 7352 33600 7404
rect 33652 7352 33658 7404
rect 33870 7352 33876 7404
rect 33928 7352 33934 7404
rect 34900 7401 34928 7432
rect 38013 7429 38025 7432
rect 38059 7429 38071 7463
rect 38013 7423 38071 7429
rect 34885 7395 34943 7401
rect 34885 7361 34897 7395
rect 34931 7392 34943 7395
rect 37553 7395 37611 7401
rect 34931 7364 36308 7392
rect 34931 7361 34943 7364
rect 34885 7355 34943 7361
rect 33686 7324 33692 7336
rect 33520 7296 33692 7324
rect 33686 7284 33692 7296
rect 33744 7284 33750 7336
rect 33888 7324 33916 7352
rect 33965 7327 34023 7333
rect 33965 7324 33977 7327
rect 33888 7296 33977 7324
rect 33965 7293 33977 7296
rect 34011 7293 34023 7327
rect 33965 7287 34023 7293
rect 26375 7160 29040 7188
rect 26375 7157 26387 7160
rect 26329 7151 26387 7157
rect 29086 7148 29092 7200
rect 29144 7148 29150 7200
rect 31294 7148 31300 7200
rect 31352 7148 31358 7200
rect 33502 7148 33508 7200
rect 33560 7148 33566 7200
rect 33980 7188 34008 7287
rect 35066 7284 35072 7336
rect 35124 7284 35130 7336
rect 36170 7284 36176 7336
rect 36228 7284 36234 7336
rect 36280 7324 36308 7364
rect 37553 7361 37565 7395
rect 37599 7392 37611 7395
rect 39132 7392 39160 7488
rect 39844 7463 39902 7469
rect 39844 7429 39856 7463
rect 39890 7460 39902 7463
rect 40512 7460 40540 7488
rect 42058 7460 42064 7472
rect 39890 7432 40540 7460
rect 40604 7432 42064 7460
rect 39890 7429 39902 7432
rect 39844 7423 39902 7429
rect 39577 7395 39635 7401
rect 39577 7392 39589 7395
rect 37599 7364 38056 7392
rect 39132 7364 39589 7392
rect 37599 7361 37611 7364
rect 37553 7355 37611 7361
rect 37568 7324 37596 7355
rect 36280 7296 37596 7324
rect 37737 7327 37795 7333
rect 37737 7293 37749 7327
rect 37783 7293 37795 7327
rect 37737 7287 37795 7293
rect 36814 7216 36820 7268
rect 36872 7216 36878 7268
rect 37752 7188 37780 7287
rect 37918 7284 37924 7336
rect 37976 7284 37982 7336
rect 38028 7324 38056 7364
rect 39577 7361 39589 7364
rect 39623 7361 39635 7395
rect 40604 7392 40632 7432
rect 42058 7420 42064 7432
rect 42116 7420 42122 7472
rect 42242 7420 42248 7472
rect 42300 7420 42306 7472
rect 42518 7420 42524 7472
rect 42576 7460 42582 7472
rect 43717 7463 43775 7469
rect 43717 7460 43729 7463
rect 42576 7432 43729 7460
rect 42576 7420 42582 7432
rect 43717 7429 43729 7432
rect 43763 7429 43775 7463
rect 45922 7460 45928 7472
rect 43717 7423 43775 7429
rect 44192 7432 45928 7460
rect 39577 7355 39635 7361
rect 39684 7364 40632 7392
rect 41417 7395 41475 7401
rect 39684 7324 39712 7364
rect 41417 7361 41429 7395
rect 41463 7392 41475 7395
rect 41782 7392 41788 7404
rect 41463 7364 41788 7392
rect 41463 7361 41475 7364
rect 41417 7355 41475 7361
rect 41782 7352 41788 7364
rect 41840 7352 41846 7404
rect 38028 7296 39712 7324
rect 41046 7284 41052 7336
rect 41104 7324 41110 7336
rect 41690 7324 41696 7336
rect 41104 7296 41696 7324
rect 41104 7284 41110 7296
rect 41690 7284 41696 7296
rect 41748 7284 41754 7336
rect 42260 7324 42288 7420
rect 42886 7352 42892 7404
rect 42944 7392 42950 7404
rect 44192 7401 44220 7432
rect 45922 7420 45928 7432
rect 45980 7420 45986 7472
rect 46017 7463 46075 7469
rect 46017 7429 46029 7463
rect 46063 7460 46075 7463
rect 47026 7460 47032 7472
rect 46063 7432 47032 7460
rect 46063 7429 46075 7432
rect 46017 7423 46075 7429
rect 47026 7420 47032 7432
rect 47084 7460 47090 7472
rect 47121 7463 47179 7469
rect 47121 7460 47133 7463
rect 47084 7432 47133 7460
rect 47084 7420 47090 7432
rect 47121 7429 47133 7432
rect 47167 7429 47179 7463
rect 47121 7423 47179 7429
rect 43625 7395 43683 7401
rect 43625 7392 43637 7395
rect 42944 7364 43637 7392
rect 42944 7352 42950 7364
rect 43625 7361 43637 7364
rect 43671 7361 43683 7395
rect 43625 7355 43683 7361
rect 44177 7395 44235 7401
rect 44177 7361 44189 7395
rect 44223 7361 44235 7395
rect 44177 7355 44235 7361
rect 44266 7352 44272 7404
rect 44324 7392 44330 7404
rect 44433 7395 44491 7401
rect 44433 7392 44445 7395
rect 44324 7364 44445 7392
rect 44324 7352 44330 7364
rect 44433 7361 44445 7364
rect 44479 7361 44491 7395
rect 44433 7355 44491 7361
rect 45554 7352 45560 7404
rect 45612 7392 45618 7404
rect 46109 7395 46167 7401
rect 46109 7392 46121 7395
rect 45612 7364 46121 7392
rect 45612 7352 45618 7364
rect 46109 7361 46121 7364
rect 46155 7392 46167 7395
rect 46382 7392 46388 7404
rect 46155 7364 46388 7392
rect 46155 7361 46167 7364
rect 46109 7355 46167 7361
rect 46382 7352 46388 7364
rect 46440 7352 46446 7404
rect 46750 7352 46756 7404
rect 46808 7392 46814 7404
rect 47872 7392 47900 7488
rect 49504 7463 49562 7469
rect 49504 7429 49516 7463
rect 49550 7460 49562 7463
rect 49878 7460 49884 7472
rect 49550 7432 49884 7460
rect 49550 7429 49562 7432
rect 49504 7423 49562 7429
rect 49878 7420 49884 7432
rect 49936 7420 49942 7472
rect 54128 7404 54156 7500
rect 54294 7488 54300 7500
rect 54352 7488 54358 7540
rect 54662 7488 54668 7540
rect 54720 7528 54726 7540
rect 54757 7531 54815 7537
rect 54757 7528 54769 7531
rect 54720 7500 54769 7528
rect 54720 7488 54726 7500
rect 54757 7497 54769 7500
rect 54803 7497 54815 7531
rect 54757 7491 54815 7497
rect 55030 7488 55036 7540
rect 55088 7488 55094 7540
rect 55122 7488 55128 7540
rect 55180 7488 55186 7540
rect 55769 7531 55827 7537
rect 55769 7497 55781 7531
rect 55815 7528 55827 7531
rect 56502 7528 56508 7540
rect 55815 7500 56508 7528
rect 55815 7497 55827 7500
rect 55769 7491 55827 7497
rect 55048 7460 55076 7488
rect 54220 7432 55076 7460
rect 46808 7364 47900 7392
rect 47949 7395 48007 7401
rect 46808 7352 46814 7364
rect 47949 7361 47961 7395
rect 47995 7392 48007 7395
rect 48590 7392 48596 7404
rect 47995 7364 48596 7392
rect 47995 7361 48007 7364
rect 47949 7355 48007 7361
rect 42521 7327 42579 7333
rect 42521 7324 42533 7327
rect 42260 7296 42533 7324
rect 42521 7293 42533 7296
rect 42567 7293 42579 7327
rect 42521 7287 42579 7293
rect 43898 7284 43904 7336
rect 43956 7324 43962 7336
rect 43956 7296 44220 7324
rect 43956 7284 43962 7296
rect 38381 7259 38439 7265
rect 38381 7225 38393 7259
rect 38427 7256 38439 7259
rect 38838 7256 38844 7268
rect 38427 7228 38844 7256
rect 38427 7225 38439 7228
rect 38381 7219 38439 7225
rect 38838 7216 38844 7228
rect 38896 7216 38902 7268
rect 43916 7256 43944 7284
rect 39224 7228 39436 7256
rect 39224 7200 39252 7228
rect 38657 7191 38715 7197
rect 38657 7188 38669 7191
rect 33980 7160 38669 7188
rect 38657 7157 38669 7160
rect 38703 7188 38715 7191
rect 39206 7188 39212 7200
rect 38703 7160 39212 7188
rect 38703 7157 38715 7160
rect 38657 7151 38715 7157
rect 39206 7148 39212 7160
rect 39264 7148 39270 7200
rect 39298 7148 39304 7200
rect 39356 7148 39362 7200
rect 39408 7188 39436 7228
rect 41386 7228 43944 7256
rect 41386 7188 41414 7228
rect 39408 7160 41414 7188
rect 41690 7148 41696 7200
rect 41748 7188 41754 7200
rect 42058 7188 42064 7200
rect 41748 7160 42064 7188
rect 41748 7148 41754 7160
rect 42058 7148 42064 7160
rect 42116 7188 42122 7200
rect 43162 7188 43168 7200
rect 42116 7160 43168 7188
rect 42116 7148 42122 7160
rect 43162 7148 43168 7160
rect 43220 7148 43226 7200
rect 43254 7148 43260 7200
rect 43312 7148 43318 7200
rect 44192 7188 44220 7296
rect 46290 7284 46296 7336
rect 46348 7284 46354 7336
rect 46474 7284 46480 7336
rect 46532 7284 46538 7336
rect 47964 7256 47992 7355
rect 48590 7352 48596 7364
rect 48648 7392 48654 7404
rect 53857 7395 53915 7401
rect 48648 7364 51948 7392
rect 48648 7352 48654 7364
rect 49237 7327 49295 7333
rect 49237 7293 49249 7327
rect 49283 7293 49295 7327
rect 49237 7287 49295 7293
rect 45112 7228 47992 7256
rect 45112 7188 45140 7228
rect 44192 7160 45140 7188
rect 45554 7148 45560 7200
rect 45612 7148 45618 7200
rect 49252 7188 49280 7287
rect 51258 7284 51264 7336
rect 51316 7324 51322 7336
rect 51920 7333 51948 7364
rect 53857 7361 53869 7395
rect 53903 7392 53915 7395
rect 53903 7364 54064 7392
rect 53903 7361 53915 7364
rect 53857 7355 53915 7361
rect 51445 7327 51503 7333
rect 51445 7324 51457 7327
rect 51316 7296 51457 7324
rect 51316 7284 51322 7296
rect 51445 7293 51457 7296
rect 51491 7293 51503 7327
rect 51445 7287 51503 7293
rect 51905 7327 51963 7333
rect 51905 7293 51917 7327
rect 51951 7293 51963 7327
rect 51905 7287 51963 7293
rect 50154 7188 50160 7200
rect 49252 7160 50160 7188
rect 50154 7148 50160 7160
rect 50212 7148 50218 7200
rect 50890 7148 50896 7200
rect 50948 7148 50954 7200
rect 51920 7188 51948 7287
rect 51994 7284 52000 7336
rect 52052 7324 52058 7336
rect 52089 7327 52147 7333
rect 52089 7324 52101 7327
rect 52052 7296 52101 7324
rect 52052 7284 52058 7296
rect 52089 7293 52101 7296
rect 52135 7293 52147 7327
rect 54036 7324 54064 7364
rect 54110 7352 54116 7404
rect 54168 7352 54174 7404
rect 54220 7324 54248 7432
rect 55140 7401 55168 7488
rect 54665 7395 54723 7401
rect 54665 7361 54677 7395
rect 54711 7392 54723 7395
rect 55125 7395 55183 7401
rect 54711 7364 55076 7392
rect 54711 7361 54723 7364
rect 54665 7355 54723 7361
rect 54036 7296 54248 7324
rect 52089 7287 52147 7293
rect 54846 7284 54852 7336
rect 54904 7284 54910 7336
rect 55048 7324 55076 7364
rect 55125 7361 55137 7395
rect 55171 7361 55183 7395
rect 55125 7355 55183 7361
rect 55784 7324 55812 7491
rect 56502 7488 56508 7500
rect 56560 7488 56566 7540
rect 56686 7488 56692 7540
rect 56744 7488 56750 7540
rect 56778 7488 56784 7540
rect 56836 7488 56842 7540
rect 57701 7531 57759 7537
rect 57701 7497 57713 7531
rect 57747 7528 57759 7531
rect 57882 7528 57888 7540
rect 57747 7500 57888 7528
rect 57747 7497 57759 7500
rect 57701 7491 57759 7497
rect 57882 7488 57888 7500
rect 57940 7488 57946 7540
rect 58158 7488 58164 7540
rect 58216 7528 58222 7540
rect 58529 7531 58587 7537
rect 58529 7528 58541 7531
rect 58216 7500 58541 7528
rect 58216 7488 58222 7500
rect 58529 7497 58541 7500
rect 58575 7497 58587 7531
rect 58529 7491 58587 7497
rect 57790 7352 57796 7404
rect 57848 7392 57854 7404
rect 57885 7395 57943 7401
rect 57885 7392 57897 7395
rect 57848 7364 57897 7392
rect 57848 7352 57854 7364
rect 57885 7361 57897 7364
rect 57931 7361 57943 7395
rect 57885 7355 57943 7361
rect 55048 7296 55812 7324
rect 56229 7327 56287 7333
rect 56229 7293 56241 7327
rect 56275 7324 56287 7327
rect 56965 7327 57023 7333
rect 56965 7324 56977 7327
rect 56275 7296 56977 7324
rect 56275 7293 56287 7296
rect 56229 7287 56287 7293
rect 56965 7293 56977 7296
rect 57011 7324 57023 7327
rect 57698 7324 57704 7336
rect 57011 7296 57704 7324
rect 57011 7293 57023 7296
rect 56965 7287 57023 7293
rect 57698 7284 57704 7296
rect 57756 7284 57762 7336
rect 52549 7259 52607 7265
rect 52549 7225 52561 7259
rect 52595 7256 52607 7259
rect 52595 7228 53236 7256
rect 52595 7225 52607 7228
rect 52549 7219 52607 7225
rect 52270 7188 52276 7200
rect 51920 7160 52276 7188
rect 52270 7148 52276 7160
rect 52328 7148 52334 7200
rect 53208 7188 53236 7228
rect 53926 7188 53932 7200
rect 53208 7160 53932 7188
rect 53926 7148 53932 7160
rect 53984 7148 53990 7200
rect 54294 7148 54300 7200
rect 54352 7148 54358 7200
rect 56318 7148 56324 7200
rect 56376 7148 56382 7200
rect 1104 7098 58880 7120
rect 1104 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 22616 7098
rect 22668 7046 22680 7098
rect 22732 7046 22744 7098
rect 22796 7046 22808 7098
rect 22860 7046 22872 7098
rect 22924 7046 37060 7098
rect 37112 7046 37124 7098
rect 37176 7046 37188 7098
rect 37240 7046 37252 7098
rect 37304 7046 37316 7098
rect 37368 7046 51504 7098
rect 51556 7046 51568 7098
rect 51620 7046 51632 7098
rect 51684 7046 51696 7098
rect 51748 7046 51760 7098
rect 51812 7046 58880 7098
rect 1104 7024 58880 7046
rect 4893 6987 4951 6993
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4939 6956 5181 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 6273 6987 6331 6993
rect 6273 6953 6285 6987
rect 6319 6984 6331 6987
rect 7374 6984 7380 6996
rect 6319 6956 7380 6984
rect 6319 6953 6331 6956
rect 6273 6947 6331 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 9677 6987 9735 6993
rect 9677 6953 9689 6987
rect 9723 6984 9735 6987
rect 10594 6984 10600 6996
rect 9723 6956 10600 6984
rect 9723 6953 9735 6956
rect 9677 6947 9735 6953
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10796 6956 10885 6984
rect 9876 6888 10640 6916
rect 3050 6848 3056 6860
rect 2700 6820 3056 6848
rect 2700 6789 2728 6820
rect 3050 6808 3056 6820
rect 3108 6848 3114 6860
rect 5442 6848 5448 6860
rect 3108 6820 5448 6848
rect 3108 6808 3114 6820
rect 3528 6792 3556 6820
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5500 6820 5549 6848
rect 5500 6808 5506 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5810 6848 5816 6860
rect 5675 6820 5816 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 5994 6808 6000 6860
rect 6052 6808 6058 6860
rect 6086 6808 6092 6860
rect 6144 6857 6150 6860
rect 6144 6851 6172 6857
rect 6160 6848 6172 6851
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 6160 6820 7573 6848
rect 6160 6817 6172 6820
rect 6144 6811 6172 6817
rect 7561 6817 7573 6820
rect 7607 6848 7619 6851
rect 7650 6848 7656 6860
rect 7607 6820 7656 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 6144 6808 6150 6811
rect 7650 6808 7656 6820
rect 7708 6848 7714 6860
rect 9766 6848 9772 6860
rect 7708 6820 9772 6848
rect 7708 6808 7714 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 2884 6712 2912 6743
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3234 6780 3240 6792
rect 3191 6752 3240 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3510 6740 3516 6792
rect 3568 6740 3574 6792
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 6825 6783 6883 6789
rect 4396 6752 6776 6780
rect 4396 6740 4402 6752
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 2884 6684 3341 6712
rect 3329 6681 3341 6684
rect 3375 6712 3387 6715
rect 3418 6712 3424 6724
rect 3375 6684 3424 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 3418 6672 3424 6684
rect 3476 6712 3482 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3476 6684 3801 6712
rect 3476 6672 3482 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 3973 6715 4031 6721
rect 3973 6712 3985 6715
rect 3936 6684 3985 6712
rect 3936 6672 3942 6684
rect 3973 6681 3985 6684
rect 4019 6681 4031 6715
rect 3973 6675 4031 6681
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 4203 6684 5181 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 6546 6712 6552 6724
rect 5684 6684 6552 6712
rect 5684 6672 5690 6684
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2004 6616 2789 6644
rect 2004 6604 2010 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 4982 6604 4988 6656
rect 5040 6604 5046 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5592 6616 5917 6644
rect 5592 6604 5598 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 6748 6644 6776 6752
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6871 6752 7021 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 7098 6780 7104 6792
rect 7055 6752 7104 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7098 6740 7104 6752
rect 7156 6780 7162 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7156 6752 7941 6780
rect 7156 6740 7162 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9876 6780 9904 6888
rect 8812 6752 9904 6780
rect 8812 6740 8818 6752
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10612 6780 10640 6888
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 10796 6848 10824 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 12250 6984 12256 6996
rect 11296 6956 12256 6984
rect 11296 6944 11302 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 15194 6984 15200 6996
rect 12406 6956 15200 6984
rect 12406 6916 12434 6956
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15436 6956 16252 6984
rect 15436 6944 15442 6956
rect 10735 6820 10824 6848
rect 10888 6888 12434 6916
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10888 6780 10916 6888
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11020 6820 11529 6848
rect 11020 6808 11026 6820
rect 11517 6817 11529 6820
rect 11563 6848 11575 6851
rect 11563 6820 12112 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 10612 6752 10916 6780
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 12084 6780 12112 6820
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12216 6820 14504 6848
rect 12216 6808 12222 6820
rect 12084 6752 12572 6780
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 9033 6715 9091 6721
rect 9033 6712 9045 6715
rect 8076 6684 9045 6712
rect 8076 6672 8082 6684
rect 9033 6681 9045 6684
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 9217 6715 9275 6721
rect 9217 6681 9229 6715
rect 9263 6712 9275 6715
rect 10594 6712 10600 6724
rect 9263 6684 10600 6712
rect 9263 6681 9275 6684
rect 9217 6675 9275 6681
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 10962 6672 10968 6724
rect 11020 6672 11026 6724
rect 11330 6672 11336 6724
rect 11388 6672 11394 6724
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 12544 6721 12572 6752
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 14366 6780 14372 6792
rect 13924 6752 14372 6780
rect 12529 6715 12587 6721
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 13924 6712 13952 6752
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14476 6789 14504 6820
rect 14550 6808 14556 6860
rect 14608 6808 14614 6860
rect 14645 6851 14703 6857
rect 14645 6817 14657 6851
rect 14691 6848 14703 6851
rect 15470 6848 15476 6860
rect 14691 6820 15476 6848
rect 14691 6817 14703 6820
rect 14645 6811 14703 6817
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14660 6712 14688 6811
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 16114 6848 16120 6860
rect 15611 6820 16120 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16224 6857 16252 6956
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18325 6987 18383 6993
rect 18325 6984 18337 6987
rect 18288 6956 18337 6984
rect 18288 6944 18294 6956
rect 18325 6953 18337 6956
rect 18371 6953 18383 6987
rect 18325 6947 18383 6953
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 20714 6984 20720 6996
rect 20671 6956 20720 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 20990 6944 20996 6996
rect 21048 6984 21054 6996
rect 21634 6984 21640 6996
rect 21048 6956 21640 6984
rect 21048 6944 21054 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22462 6944 22468 6996
rect 22520 6984 22526 6996
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22520 6956 22937 6984
rect 22520 6944 22526 6956
rect 22925 6953 22937 6956
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 23014 6944 23020 6996
rect 23072 6944 23078 6996
rect 24394 6944 24400 6996
rect 24452 6984 24458 6996
rect 24489 6987 24547 6993
rect 24489 6984 24501 6987
rect 24452 6956 24501 6984
rect 24452 6944 24458 6956
rect 24489 6953 24501 6956
rect 24535 6953 24547 6987
rect 24489 6947 24547 6953
rect 24964 6956 27844 6984
rect 23032 6916 23060 6944
rect 24964 6916 24992 6956
rect 17512 6888 17724 6916
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16602 6851 16660 6857
rect 16602 6848 16614 6851
rect 16356 6820 16614 6848
rect 16356 6808 16362 6820
rect 16602 6817 16614 6820
rect 16648 6817 16660 6851
rect 16602 6811 16660 6817
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17512 6848 17540 6888
rect 17696 6860 17724 6888
rect 22112 6888 23060 6916
rect 23952 6888 24992 6916
rect 16807 6820 17540 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17586 6808 17592 6860
rect 17644 6808 17650 6860
rect 17678 6808 17684 6860
rect 17736 6808 17742 6860
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 19058 6848 19064 6860
rect 18380 6820 19064 6848
rect 18380 6808 18386 6820
rect 19058 6808 19064 6820
rect 19116 6848 19122 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19116 6820 19257 6848
rect 19116 6808 19122 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 22112 6848 22140 6888
rect 23952 6860 23980 6888
rect 21039 6820 22140 6848
rect 22189 6851 22247 6857
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 22189 6817 22201 6851
rect 22235 6848 22247 6851
rect 22235 6820 22508 6848
rect 22235 6817 22247 6820
rect 22189 6811 22247 6817
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 12575 6684 13952 6712
rect 14016 6684 14688 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 6748 6616 10057 6644
rect 5905 6607 5963 6613
rect 10045 6613 10057 6616
rect 10091 6644 10103 6647
rect 10980 6644 11008 6672
rect 10091 6616 11008 6644
rect 11348 6644 11376 6672
rect 11790 6644 11796 6656
rect 11348 6616 11796 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 11790 6604 11796 6616
rect 11848 6644 11854 6656
rect 12176 6644 12204 6672
rect 14016 6656 14044 6684
rect 11848 6616 12204 6644
rect 11848 6604 11854 6616
rect 12986 6604 12992 6656
rect 13044 6604 13050 6656
rect 13906 6604 13912 6656
rect 13964 6604 13970 6656
rect 13998 6604 14004 6656
rect 14056 6604 14062 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 15764 6644 15792 6743
rect 16482 6740 16488 6792
rect 16540 6740 16546 6792
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 18046 6780 18052 6792
rect 17451 6752 18052 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 18248 6752 18889 6780
rect 17862 6712 17868 6724
rect 17236 6684 17868 6712
rect 17236 6644 17264 6684
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 15764 6616 17264 6644
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 18248 6653 18276 6752
rect 18877 6749 18889 6752
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19501 6783 19559 6789
rect 19501 6780 19513 6783
rect 19392 6752 19513 6780
rect 19392 6740 19398 6752
rect 19501 6749 19513 6752
rect 19547 6749 19559 6783
rect 19501 6743 19559 6749
rect 21634 6740 21640 6792
rect 21692 6740 21698 6792
rect 21726 6740 21732 6792
rect 21784 6789 21790 6792
rect 21784 6783 21833 6789
rect 21784 6749 21787 6783
rect 21821 6749 21833 6783
rect 21784 6743 21833 6749
rect 21784 6740 21790 6743
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22480 6780 22508 6820
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 22612 6820 22661 6848
rect 22612 6808 22618 6820
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 22833 6851 22891 6857
rect 22833 6817 22845 6851
rect 22879 6848 22891 6851
rect 23198 6848 23204 6860
rect 22879 6820 23204 6848
rect 22879 6817 22891 6820
rect 22833 6811 22891 6817
rect 23198 6808 23204 6820
rect 23256 6848 23262 6860
rect 23385 6851 23443 6857
rect 23385 6848 23397 6851
rect 23256 6820 23397 6848
rect 23256 6808 23262 6820
rect 23385 6817 23397 6820
rect 23431 6817 23443 6851
rect 23385 6811 23443 6817
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 23934 6808 23940 6860
rect 23992 6808 23998 6860
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26326 6848 26332 6860
rect 26283 6820 26332 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26326 6808 26332 6820
rect 26384 6808 26390 6860
rect 26421 6851 26479 6857
rect 26421 6817 26433 6851
rect 26467 6848 26479 6851
rect 26602 6848 26608 6860
rect 26467 6820 26608 6848
rect 26467 6817 26479 6820
rect 26421 6811 26479 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 26881 6851 26939 6857
rect 26881 6848 26893 6851
rect 26844 6820 26893 6848
rect 26844 6808 26850 6820
rect 26881 6817 26893 6820
rect 26927 6817 26939 6851
rect 26881 6811 26939 6817
rect 26970 6808 26976 6860
rect 27028 6848 27034 6860
rect 27274 6851 27332 6857
rect 27274 6848 27286 6851
rect 27028 6820 27286 6848
rect 27028 6808 27034 6820
rect 27274 6817 27286 6820
rect 27320 6817 27332 6851
rect 27274 6811 27332 6817
rect 27433 6851 27491 6857
rect 27433 6817 27445 6851
rect 27479 6848 27491 6851
rect 27614 6848 27620 6860
rect 27479 6820 27620 6848
rect 27479 6817 27491 6820
rect 27433 6811 27491 6817
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 27816 6848 27844 6956
rect 28534 6944 28540 6996
rect 28592 6984 28598 6996
rect 32582 6984 32588 6996
rect 28592 6956 32588 6984
rect 28592 6944 28598 6956
rect 32582 6944 32588 6956
rect 32640 6944 32646 6996
rect 33594 6944 33600 6996
rect 33652 6984 33658 6996
rect 35621 6987 35679 6993
rect 35621 6984 35633 6987
rect 33652 6956 35633 6984
rect 33652 6944 33658 6956
rect 35621 6953 35633 6956
rect 35667 6953 35679 6987
rect 35621 6947 35679 6953
rect 36924 6956 37872 6984
rect 33318 6916 33324 6928
rect 32600 6888 33324 6916
rect 27982 6848 27988 6860
rect 27816 6820 27988 6848
rect 27982 6808 27988 6820
rect 28040 6848 28046 6860
rect 28261 6851 28319 6857
rect 28261 6848 28273 6851
rect 28040 6820 28273 6848
rect 28040 6808 28046 6820
rect 28261 6817 28273 6820
rect 28307 6817 28319 6851
rect 31938 6848 31944 6860
rect 28261 6811 28319 6817
rect 31496 6820 31944 6848
rect 31496 6792 31524 6820
rect 31938 6808 31944 6820
rect 31996 6808 32002 6860
rect 32125 6851 32183 6857
rect 32125 6817 32137 6851
rect 32171 6848 32183 6851
rect 32600 6848 32628 6888
rect 33318 6876 33324 6888
rect 33376 6876 33382 6928
rect 34146 6916 34152 6928
rect 33612 6888 34152 6916
rect 32171 6820 32628 6848
rect 32677 6851 32735 6857
rect 32171 6817 32183 6820
rect 32125 6811 32183 6817
rect 32677 6817 32689 6851
rect 32723 6848 32735 6851
rect 33612 6848 33640 6888
rect 34146 6876 34152 6888
rect 34204 6916 34210 6928
rect 35066 6916 35072 6928
rect 34204 6888 35072 6916
rect 34204 6876 34210 6888
rect 35066 6876 35072 6888
rect 35124 6916 35130 6928
rect 36722 6916 36728 6928
rect 35124 6888 36728 6916
rect 35124 6876 35130 6888
rect 36722 6876 36728 6888
rect 36780 6916 36786 6928
rect 36924 6925 36952 6956
rect 36909 6919 36967 6925
rect 36909 6916 36921 6919
rect 36780 6888 36921 6916
rect 36780 6876 36786 6888
rect 36909 6885 36921 6888
rect 36955 6885 36967 6919
rect 37844 6916 37872 6956
rect 37918 6944 37924 6996
rect 37976 6984 37982 6996
rect 38105 6987 38163 6993
rect 38105 6984 38117 6987
rect 37976 6956 38117 6984
rect 37976 6944 37982 6956
rect 38105 6953 38117 6956
rect 38151 6953 38163 6987
rect 38105 6947 38163 6953
rect 41046 6944 41052 6996
rect 41104 6944 41110 6996
rect 41156 6956 43116 6984
rect 38381 6919 38439 6925
rect 38381 6916 38393 6919
rect 37844 6888 38393 6916
rect 36909 6879 36967 6885
rect 38381 6885 38393 6888
rect 38427 6916 38439 6919
rect 38427 6888 38516 6916
rect 38427 6885 38439 6888
rect 38381 6879 38439 6885
rect 32723 6820 33640 6848
rect 32723 6817 32735 6820
rect 32677 6811 32735 6817
rect 33686 6808 33692 6860
rect 33744 6848 33750 6860
rect 34701 6851 34759 6857
rect 34701 6848 34713 6851
rect 33744 6820 34713 6848
rect 33744 6808 33750 6820
rect 34701 6817 34713 6820
rect 34747 6817 34759 6851
rect 35805 6851 35863 6857
rect 35805 6848 35817 6851
rect 34701 6811 34759 6817
rect 34808 6820 35817 6848
rect 25613 6783 25671 6789
rect 22480 6752 23152 6780
rect 23124 6724 23152 6752
rect 25613 6749 25625 6783
rect 25659 6780 25671 6783
rect 25774 6780 25780 6792
rect 25659 6752 25780 6780
rect 25659 6749 25671 6752
rect 25613 6743 25671 6749
rect 25774 6740 25780 6752
rect 25832 6740 25838 6792
rect 25866 6740 25872 6792
rect 25924 6740 25930 6792
rect 27154 6740 27160 6792
rect 27212 6740 27218 6792
rect 28074 6740 28080 6792
rect 28132 6780 28138 6792
rect 28537 6783 28595 6789
rect 28537 6780 28549 6783
rect 28132 6752 28549 6780
rect 28132 6740 28138 6752
rect 28537 6749 28549 6752
rect 28583 6749 28595 6783
rect 28537 6743 28595 6749
rect 31133 6783 31191 6789
rect 31133 6749 31145 6783
rect 31179 6780 31191 6783
rect 31294 6780 31300 6792
rect 31179 6752 31300 6780
rect 31179 6749 31191 6752
rect 31133 6743 31191 6749
rect 31294 6740 31300 6752
rect 31352 6740 31358 6792
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6780 31447 6783
rect 31478 6780 31484 6792
rect 31435 6752 31484 6780
rect 31435 6749 31447 6752
rect 31389 6743 31447 6749
rect 31478 6740 31484 6752
rect 31536 6740 31542 6792
rect 32306 6789 32312 6792
rect 32284 6783 32312 6789
rect 32284 6749 32296 6783
rect 32284 6743 32312 6749
rect 32306 6740 32312 6743
rect 32364 6740 32370 6792
rect 32398 6740 32404 6792
rect 32456 6740 32462 6792
rect 33134 6740 33140 6792
rect 33192 6740 33198 6792
rect 33318 6740 33324 6792
rect 33376 6740 33382 6792
rect 33505 6783 33563 6789
rect 33505 6749 33517 6783
rect 33551 6749 33563 6783
rect 33505 6743 33563 6749
rect 23106 6672 23112 6724
rect 23164 6712 23170 6724
rect 23164 6684 24256 6712
rect 23164 6672 23170 6684
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 20990 6604 20996 6656
rect 21048 6644 21054 6656
rect 22278 6644 22284 6656
rect 21048 6616 22284 6644
rect 21048 6604 21054 6616
rect 22278 6604 22284 6616
rect 22336 6644 22342 6656
rect 23198 6644 23204 6656
rect 22336 6616 23204 6644
rect 22336 6604 22342 6616
rect 23198 6604 23204 6616
rect 23256 6644 23262 6656
rect 24228 6653 24256 6684
rect 24670 6672 24676 6724
rect 24728 6712 24734 6724
rect 25884 6712 25912 6740
rect 24728 6684 25912 6712
rect 24728 6672 24734 6684
rect 23293 6647 23351 6653
rect 23293 6644 23305 6647
rect 23256 6616 23305 6644
rect 23256 6604 23262 6616
rect 23293 6613 23305 6616
rect 23339 6613 23351 6647
rect 23293 6607 23351 6613
rect 24213 6647 24271 6653
rect 24213 6613 24225 6647
rect 24259 6644 24271 6647
rect 26786 6644 26792 6656
rect 24259 6616 26792 6644
rect 24259 6613 24271 6616
rect 24213 6607 24271 6613
rect 26786 6604 26792 6616
rect 26844 6644 26850 6656
rect 27062 6644 27068 6656
rect 26844 6616 27068 6644
rect 26844 6604 26850 6616
rect 27062 6604 27068 6616
rect 27120 6604 27126 6656
rect 28077 6647 28135 6653
rect 28077 6613 28089 6647
rect 28123 6644 28135 6647
rect 28445 6647 28503 6653
rect 28445 6644 28457 6647
rect 28123 6616 28457 6644
rect 28123 6613 28135 6616
rect 28077 6607 28135 6613
rect 28445 6613 28457 6616
rect 28491 6613 28503 6647
rect 28445 6607 28503 6613
rect 28902 6604 28908 6656
rect 28960 6604 28966 6656
rect 30009 6647 30067 6653
rect 30009 6613 30021 6647
rect 30055 6644 30067 6647
rect 30558 6644 30564 6656
rect 30055 6616 30564 6644
rect 30055 6613 30067 6616
rect 30009 6607 30067 6613
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31481 6647 31539 6653
rect 31481 6613 31493 6647
rect 31527 6644 31539 6647
rect 31662 6644 31668 6656
rect 31527 6616 31668 6644
rect 31527 6613 31539 6616
rect 31481 6607 31539 6613
rect 31662 6604 31668 6616
rect 31720 6604 31726 6656
rect 32582 6604 32588 6656
rect 32640 6644 32646 6656
rect 33520 6644 33548 6743
rect 33962 6740 33968 6792
rect 34020 6780 34026 6792
rect 34808 6780 34836 6820
rect 35805 6817 35817 6820
rect 35851 6817 35863 6851
rect 35805 6811 35863 6817
rect 36170 6808 36176 6860
rect 36228 6808 36234 6860
rect 36265 6851 36323 6857
rect 36265 6817 36277 6851
rect 36311 6848 36323 6851
rect 36354 6848 36360 6860
rect 36311 6820 36360 6848
rect 36311 6817 36323 6820
rect 36265 6811 36323 6817
rect 36354 6808 36360 6820
rect 36412 6808 36418 6860
rect 36446 6808 36452 6860
rect 36504 6808 36510 6860
rect 36998 6808 37004 6860
rect 37056 6848 37062 6860
rect 37302 6851 37360 6857
rect 37302 6848 37314 6851
rect 37056 6820 37314 6848
rect 37056 6808 37062 6820
rect 37302 6817 37314 6820
rect 37348 6817 37360 6851
rect 37302 6811 37360 6817
rect 37461 6851 37519 6857
rect 37461 6817 37473 6851
rect 37507 6848 37519 6851
rect 37642 6848 37648 6860
rect 37507 6820 37648 6848
rect 37507 6817 37519 6820
rect 37461 6811 37519 6817
rect 37642 6808 37648 6820
rect 37700 6808 37706 6860
rect 34020 6752 34836 6780
rect 34020 6740 34026 6752
rect 35250 6740 35256 6792
rect 35308 6740 35314 6792
rect 36188 6780 36216 6808
rect 35912 6752 36216 6780
rect 34241 6715 34299 6721
rect 34241 6681 34253 6715
rect 34287 6712 34299 6715
rect 34698 6712 34704 6724
rect 34287 6684 34704 6712
rect 34287 6681 34299 6684
rect 34241 6675 34299 6681
rect 34698 6672 34704 6684
rect 34756 6712 34762 6724
rect 35912 6712 35940 6752
rect 37182 6740 37188 6792
rect 37240 6740 37246 6792
rect 34756 6684 35940 6712
rect 34756 6672 34762 6684
rect 35986 6672 35992 6724
rect 36044 6672 36050 6724
rect 32640 6616 33548 6644
rect 38488 6644 38516 6888
rect 38608 6808 38614 6860
rect 38666 6848 38672 6860
rect 38749 6851 38807 6857
rect 38749 6848 38761 6851
rect 38666 6820 38761 6848
rect 38666 6808 38672 6820
rect 38749 6817 38761 6820
rect 38795 6817 38807 6851
rect 38749 6811 38807 6817
rect 38930 6808 38936 6860
rect 38988 6848 38994 6860
rect 39577 6851 39635 6857
rect 39577 6848 39589 6851
rect 38988 6820 39589 6848
rect 38988 6808 38994 6820
rect 39577 6817 39589 6820
rect 39623 6848 39635 6851
rect 40589 6851 40647 6857
rect 40589 6848 40601 6851
rect 39623 6820 40601 6848
rect 39623 6817 39635 6820
rect 39577 6811 39635 6817
rect 40589 6817 40601 6820
rect 40635 6848 40647 6851
rect 41156 6848 41184 6956
rect 40635 6820 41184 6848
rect 40635 6817 40647 6820
rect 40589 6811 40647 6817
rect 41966 6808 41972 6860
rect 42024 6857 42030 6860
rect 42024 6851 42073 6857
rect 42024 6817 42027 6851
rect 42061 6817 42073 6851
rect 42024 6811 42073 6817
rect 42024 6808 42030 6811
rect 42426 6808 42432 6860
rect 42484 6808 42490 6860
rect 42889 6851 42947 6857
rect 42889 6817 42901 6851
rect 42935 6848 42947 6851
rect 42978 6848 42984 6860
rect 42935 6820 42984 6848
rect 42935 6817 42947 6820
rect 42889 6811 42947 6817
rect 42978 6808 42984 6820
rect 43036 6808 43042 6860
rect 43088 6848 43116 6956
rect 46198 6944 46204 6996
rect 46256 6944 46262 6996
rect 46382 6944 46388 6996
rect 46440 6984 46446 6996
rect 46477 6987 46535 6993
rect 46477 6984 46489 6987
rect 46440 6956 46489 6984
rect 46440 6944 46446 6956
rect 46477 6953 46489 6956
rect 46523 6984 46535 6987
rect 47302 6984 47308 6996
rect 46523 6956 47308 6984
rect 46523 6953 46535 6956
rect 46477 6947 46535 6953
rect 47302 6944 47308 6956
rect 47360 6944 47366 6996
rect 49786 6944 49792 6996
rect 49844 6984 49850 6996
rect 50341 6987 50399 6993
rect 50341 6984 50353 6987
rect 49844 6956 50353 6984
rect 49844 6944 49850 6956
rect 50341 6953 50353 6956
rect 50387 6984 50399 6987
rect 50387 6956 51856 6984
rect 50387 6953 50399 6956
rect 50341 6947 50399 6953
rect 47854 6876 47860 6928
rect 47912 6916 47918 6928
rect 47912 6888 49924 6916
rect 47912 6876 47918 6888
rect 43088 6820 43208 6848
rect 41874 6740 41880 6792
rect 41932 6740 41938 6792
rect 42150 6740 42156 6792
rect 42208 6740 42214 6792
rect 43073 6783 43131 6789
rect 43073 6749 43085 6783
rect 43119 6749 43131 6783
rect 43180 6780 43208 6820
rect 43254 6808 43260 6860
rect 43312 6848 43318 6860
rect 43717 6851 43775 6857
rect 43717 6848 43729 6851
rect 43312 6820 43729 6848
rect 43312 6808 43318 6820
rect 43717 6817 43729 6820
rect 43763 6817 43775 6851
rect 43717 6811 43775 6817
rect 45554 6808 45560 6860
rect 45612 6808 45618 6860
rect 47765 6851 47823 6857
rect 47765 6817 47777 6851
rect 47811 6848 47823 6851
rect 48038 6848 48044 6860
rect 47811 6820 48044 6848
rect 47811 6817 47823 6820
rect 47765 6811 47823 6817
rect 48038 6808 48044 6820
rect 48096 6808 48102 6860
rect 49896 6857 49924 6888
rect 49881 6851 49939 6857
rect 49881 6817 49893 6851
rect 49927 6848 49939 6851
rect 51353 6851 51411 6857
rect 51353 6848 51365 6851
rect 49927 6820 51365 6848
rect 49927 6817 49939 6820
rect 49881 6811 49939 6817
rect 51353 6817 51365 6820
rect 51399 6817 51411 6851
rect 51353 6811 51411 6817
rect 51442 6808 51448 6860
rect 51500 6857 51506 6860
rect 51500 6851 51549 6857
rect 51500 6817 51503 6851
rect 51537 6817 51549 6851
rect 51828 6848 51856 6956
rect 54202 6944 54208 6996
rect 54260 6944 54266 6996
rect 56781 6987 56839 6993
rect 56781 6953 56793 6987
rect 56827 6984 56839 6987
rect 57054 6984 57060 6996
rect 56827 6956 57060 6984
rect 56827 6953 56839 6956
rect 56781 6947 56839 6953
rect 57054 6944 57060 6956
rect 57112 6944 57118 6996
rect 51905 6851 51963 6857
rect 51905 6848 51917 6851
rect 51828 6820 51917 6848
rect 51500 6811 51549 6817
rect 51905 6817 51917 6820
rect 51951 6817 51963 6851
rect 51905 6811 51963 6817
rect 52365 6851 52423 6857
rect 52365 6817 52377 6851
rect 52411 6848 52423 6851
rect 52822 6848 52828 6860
rect 52411 6820 52828 6848
rect 52411 6817 52423 6820
rect 52365 6811 52423 6817
rect 51500 6808 51506 6811
rect 52822 6808 52828 6820
rect 52880 6808 52886 6860
rect 53926 6808 53932 6860
rect 53984 6808 53990 6860
rect 54294 6808 54300 6860
rect 54352 6848 54358 6860
rect 54757 6851 54815 6857
rect 54757 6848 54769 6851
rect 54352 6820 54769 6848
rect 54352 6808 54358 6820
rect 54757 6817 54769 6820
rect 54803 6817 54815 6851
rect 54757 6811 54815 6817
rect 56229 6851 56287 6857
rect 56229 6817 56241 6851
rect 56275 6848 56287 6851
rect 56318 6848 56324 6860
rect 56275 6820 56324 6848
rect 56275 6817 56287 6820
rect 56229 6811 56287 6817
rect 56318 6808 56324 6820
rect 56376 6808 56382 6860
rect 57422 6808 57428 6860
rect 57480 6808 57486 6860
rect 58345 6851 58403 6857
rect 58345 6817 58357 6851
rect 58391 6848 58403 6851
rect 58434 6848 58440 6860
rect 58391 6820 58440 6848
rect 58391 6817 58403 6820
rect 58345 6811 58403 6817
rect 58434 6808 58440 6820
rect 58492 6808 58498 6860
rect 44634 6780 44640 6792
rect 43180 6752 44640 6780
rect 43073 6743 43131 6749
rect 38930 6672 38936 6724
rect 38988 6672 38994 6724
rect 40126 6712 40132 6724
rect 39960 6684 40132 6712
rect 39960 6644 39988 6684
rect 40126 6672 40132 6684
rect 40184 6672 40190 6724
rect 40497 6715 40555 6721
rect 40497 6681 40509 6715
rect 40543 6712 40555 6715
rect 41322 6712 41328 6724
rect 40543 6684 41328 6712
rect 40543 6681 40555 6684
rect 40497 6675 40555 6681
rect 41322 6672 41328 6684
rect 41380 6672 41386 6724
rect 38488 6616 39988 6644
rect 32640 6604 32646 6616
rect 40034 6604 40040 6656
rect 40092 6604 40098 6656
rect 40402 6604 40408 6656
rect 40460 6604 40466 6656
rect 41233 6647 41291 6653
rect 41233 6613 41245 6647
rect 41279 6644 41291 6647
rect 42518 6644 42524 6656
rect 41279 6616 42524 6644
rect 41279 6613 41291 6616
rect 41233 6607 41291 6613
rect 42518 6604 42524 6616
rect 42576 6604 42582 6656
rect 42610 6604 42616 6656
rect 42668 6644 42674 6656
rect 43088 6644 43116 6743
rect 44634 6740 44640 6752
rect 44692 6740 44698 6792
rect 46842 6740 46848 6792
rect 46900 6780 46906 6792
rect 47857 6783 47915 6789
rect 47857 6780 47869 6783
rect 46900 6752 47869 6780
rect 46900 6740 46906 6752
rect 47857 6749 47869 6752
rect 47903 6749 47915 6783
rect 47857 6743 47915 6749
rect 48406 6740 48412 6792
rect 48464 6740 48470 6792
rect 49145 6783 49203 6789
rect 49145 6749 49157 6783
rect 49191 6749 49203 6783
rect 49145 6743 49203 6749
rect 43254 6672 43260 6724
rect 43312 6712 43318 6724
rect 45465 6715 45523 6721
rect 45465 6712 45477 6715
rect 43312 6684 45477 6712
rect 43312 6672 43318 6684
rect 45465 6681 45477 6684
rect 45511 6712 45523 6715
rect 46290 6712 46296 6724
rect 45511 6684 46296 6712
rect 45511 6681 45523 6684
rect 45465 6675 45523 6681
rect 46290 6672 46296 6684
rect 46348 6672 46354 6724
rect 46382 6672 46388 6724
rect 46440 6672 46446 6724
rect 47394 6672 47400 6724
rect 47452 6712 47458 6724
rect 49160 6712 49188 6743
rect 51626 6740 51632 6792
rect 51684 6740 51690 6792
rect 52549 6783 52607 6789
rect 52549 6749 52561 6783
rect 52595 6749 52607 6783
rect 52549 6743 52607 6749
rect 47452 6684 49188 6712
rect 47452 6672 47458 6684
rect 42668 6616 43116 6644
rect 42668 6604 42674 6616
rect 43162 6604 43168 6656
rect 43220 6604 43226 6656
rect 47026 6604 47032 6656
rect 47084 6644 47090 6656
rect 47121 6647 47179 6653
rect 47121 6644 47133 6647
rect 47084 6616 47133 6644
rect 47084 6604 47090 6616
rect 47121 6613 47133 6616
rect 47167 6613 47179 6647
rect 47121 6607 47179 6613
rect 47946 6604 47952 6656
rect 48004 6644 48010 6656
rect 48593 6647 48651 6653
rect 48593 6644 48605 6647
rect 48004 6616 48605 6644
rect 48004 6604 48010 6616
rect 48593 6613 48605 6616
rect 48639 6613 48651 6647
rect 48593 6607 48651 6613
rect 50709 6647 50767 6653
rect 50709 6613 50721 6647
rect 50755 6644 50767 6647
rect 51994 6644 52000 6656
rect 50755 6616 52000 6644
rect 50755 6613 50767 6616
rect 50709 6607 50767 6613
rect 51994 6604 52000 6616
rect 52052 6604 52058 6656
rect 52178 6604 52184 6656
rect 52236 6644 52242 6656
rect 52564 6644 52592 6743
rect 52638 6740 52644 6792
rect 52696 6780 52702 6792
rect 53193 6783 53251 6789
rect 53193 6780 53205 6783
rect 52696 6752 53205 6780
rect 52696 6740 52702 6752
rect 53193 6749 53205 6752
rect 53239 6749 53251 6783
rect 53193 6743 53251 6749
rect 55122 6740 55128 6792
rect 55180 6780 55186 6792
rect 56594 6780 56600 6792
rect 55180 6752 56600 6780
rect 55180 6740 55186 6752
rect 56594 6740 56600 6752
rect 56652 6780 56658 6792
rect 57333 6783 57391 6789
rect 57333 6780 57345 6783
rect 56652 6752 57345 6780
rect 56652 6740 56658 6752
rect 57333 6749 57345 6752
rect 57379 6780 57391 6783
rect 57941 6783 57999 6789
rect 57941 6780 57953 6783
rect 57379 6752 57953 6780
rect 57379 6749 57391 6752
rect 57333 6743 57391 6749
rect 57941 6749 57953 6752
rect 57987 6749 57999 6783
rect 57941 6743 57999 6749
rect 56870 6672 56876 6724
rect 56928 6672 56934 6724
rect 57606 6672 57612 6724
rect 57664 6672 57670 6724
rect 57698 6672 57704 6724
rect 57756 6712 57762 6724
rect 58069 6715 58127 6721
rect 58069 6712 58081 6715
rect 57756 6684 58081 6712
rect 57756 6672 57762 6684
rect 58069 6681 58081 6684
rect 58115 6681 58127 6715
rect 58069 6675 58127 6681
rect 58161 6715 58219 6721
rect 58161 6681 58173 6715
rect 58207 6681 58219 6715
rect 58161 6675 58219 6681
rect 52641 6647 52699 6653
rect 52641 6644 52653 6647
rect 52236 6616 52653 6644
rect 52236 6604 52242 6616
rect 52641 6613 52653 6616
rect 52687 6613 52699 6647
rect 52641 6607 52699 6613
rect 53374 6604 53380 6656
rect 53432 6604 53438 6656
rect 55582 6604 55588 6656
rect 55640 6604 55646 6656
rect 56597 6647 56655 6653
rect 56597 6613 56609 6647
rect 56643 6644 56655 6647
rect 57238 6644 57244 6656
rect 56643 6616 57244 6644
rect 56643 6613 56655 6616
rect 56597 6607 56655 6613
rect 57238 6604 57244 6616
rect 57296 6644 57302 6656
rect 58176 6644 58204 6675
rect 58250 6672 58256 6724
rect 58308 6712 58314 6724
rect 58345 6715 58403 6721
rect 58345 6712 58357 6715
rect 58308 6684 58357 6712
rect 58308 6672 58314 6684
rect 58345 6681 58357 6684
rect 58391 6681 58403 6715
rect 58345 6675 58403 6681
rect 57296 6616 58204 6644
rect 57296 6604 57302 6616
rect 1104 6554 59040 6576
rect 1104 6502 15394 6554
rect 15446 6502 15458 6554
rect 15510 6502 15522 6554
rect 15574 6502 15586 6554
rect 15638 6502 15650 6554
rect 15702 6502 29838 6554
rect 29890 6502 29902 6554
rect 29954 6502 29966 6554
rect 30018 6502 30030 6554
rect 30082 6502 30094 6554
rect 30146 6502 44282 6554
rect 44334 6502 44346 6554
rect 44398 6502 44410 6554
rect 44462 6502 44474 6554
rect 44526 6502 44538 6554
rect 44590 6502 58726 6554
rect 58778 6502 58790 6554
rect 58842 6502 58854 6554
rect 58906 6502 58918 6554
rect 58970 6502 58982 6554
rect 59034 6502 59040 6554
rect 1104 6480 59040 6502
rect 3418 6400 3424 6452
rect 3476 6400 3482 6452
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 4246 6440 4252 6452
rect 3651 6412 4252 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6052 6412 6745 6440
rect 6052 6400 6058 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 8665 6443 8723 6449
rect 8665 6409 8677 6443
rect 8711 6440 8723 6443
rect 8938 6440 8944 6452
rect 8711 6412 8944 6440
rect 8711 6409 8723 6412
rect 8665 6403 8723 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 11241 6443 11299 6449
rect 11241 6409 11253 6443
rect 11287 6440 11299 6443
rect 11974 6440 11980 6452
rect 11287 6412 11980 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12066 6400 12072 6452
rect 12124 6400 12130 6452
rect 12986 6400 12992 6452
rect 13044 6400 13050 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 14093 6443 14151 6449
rect 14093 6440 14105 6443
rect 13412 6412 14105 6440
rect 13412 6400 13418 6412
rect 14093 6409 14105 6412
rect 14139 6409 14151 6443
rect 14093 6403 14151 6409
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 14332 6412 14473 6440
rect 14332 6400 14338 6412
rect 14461 6409 14473 6412
rect 14507 6440 14519 6443
rect 16482 6440 16488 6452
rect 14507 6412 16488 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 17770 6440 17776 6452
rect 17144 6412 17776 6440
rect 3436 6313 3464 6400
rect 3528 6344 3740 6372
rect 3528 6316 3556 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 3421 6307 3479 6313
rect 1627 6276 2774 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1854 6196 1860 6248
rect 1912 6196 1918 6248
rect 2746 6168 2774 6276
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3712 6313 3740 6344
rect 4264 6313 4292 6400
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 5000 6304 5028 6400
rect 11698 6372 11704 6384
rect 5644 6344 11704 6372
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 5000 6276 5089 6304
rect 4249 6267 4307 6273
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 3620 6236 3648 6267
rect 3878 6236 3884 6248
rect 3620 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 5644 6236 5672 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5960 6276 6377 6304
rect 5960 6264 5966 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7552 6307 7610 6313
rect 7552 6273 7564 6307
rect 7598 6304 7610 6307
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 7598 6276 8769 6304
rect 7598 6273 7610 6276
rect 7552 6267 7610 6273
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8904 6276 8953 6304
rect 8904 6264 8910 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9766 6304 9772 6316
rect 9263 6276 9772 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12434 6304 12440 6316
rect 12207 6276 12440 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12434 6264 12440 6276
rect 12492 6304 12498 6316
rect 12894 6304 12900 6316
rect 12492 6276 12900 6304
rect 12492 6264 12498 6276
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 4479 6208 5672 6236
rect 5813 6239 5871 6245
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5859 6208 5948 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5920 6180 5948 6208
rect 7282 6196 7288 6248
rect 7340 6196 7346 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10962 6236 10968 6248
rect 10652 6208 10968 6236
rect 10652 6196 10658 6208
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 2746 6140 4108 6168
rect 4080 6112 4108 6140
rect 5258 6128 5264 6180
rect 5316 6128 5322 6180
rect 5442 6128 5448 6180
rect 5500 6128 5506 6180
rect 5626 6128 5632 6180
rect 5684 6128 5690 6180
rect 5902 6128 5908 6180
rect 5960 6128 5966 6180
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 12342 6168 12348 6180
rect 9723 6140 12348 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 12342 6128 12348 6140
rect 12400 6168 12406 6180
rect 13004 6168 13032 6400
rect 14553 6375 14611 6381
rect 14553 6341 14565 6375
rect 14599 6372 14611 6375
rect 16022 6372 16028 6384
rect 14599 6344 16028 6372
rect 14599 6341 14611 6344
rect 14553 6335 14611 6341
rect 16022 6332 16028 6344
rect 16080 6372 16086 6384
rect 17144 6381 17172 6412
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18141 6443 18199 6449
rect 18141 6440 18153 6443
rect 17920 6412 18153 6440
rect 17920 6400 17926 6412
rect 18141 6409 18153 6412
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 20990 6400 20996 6452
rect 21048 6400 21054 6452
rect 21637 6443 21695 6449
rect 21637 6409 21649 6443
rect 21683 6440 21695 6443
rect 23106 6440 23112 6452
rect 21683 6412 23112 6440
rect 21683 6409 21695 6412
rect 21637 6403 21695 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23201 6443 23259 6449
rect 23201 6409 23213 6443
rect 23247 6440 23259 6443
rect 23382 6440 23388 6452
rect 23247 6412 23388 6440
rect 23247 6409 23259 6412
rect 23201 6403 23259 6409
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 26326 6400 26332 6452
rect 26384 6440 26390 6452
rect 26973 6443 27031 6449
rect 26973 6440 26985 6443
rect 26384 6412 26985 6440
rect 26384 6400 26390 6412
rect 26973 6409 26985 6412
rect 27019 6409 27031 6443
rect 26973 6403 27031 6409
rect 27982 6400 27988 6452
rect 28040 6400 28046 6452
rect 28626 6400 28632 6452
rect 28684 6440 28690 6452
rect 28721 6443 28779 6449
rect 28721 6440 28733 6443
rect 28684 6412 28733 6440
rect 28684 6400 28690 6412
rect 28721 6409 28733 6412
rect 28767 6409 28779 6443
rect 28721 6403 28779 6409
rect 30650 6400 30656 6452
rect 30708 6440 30714 6452
rect 31021 6443 31079 6449
rect 31021 6440 31033 6443
rect 30708 6412 31033 6440
rect 30708 6400 30714 6412
rect 31021 6409 31033 6412
rect 31067 6409 31079 6443
rect 31021 6403 31079 6409
rect 31481 6443 31539 6449
rect 31481 6409 31493 6443
rect 31527 6409 31539 6443
rect 31481 6403 31539 6409
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 16080 6344 17141 6372
rect 16080 6332 16086 6344
rect 17129 6341 17141 6344
rect 17175 6341 17187 6375
rect 17129 6335 17187 6341
rect 17313 6375 17371 6381
rect 17313 6341 17325 6375
rect 17359 6372 17371 6375
rect 18322 6372 18328 6384
rect 17359 6344 18328 6372
rect 17359 6341 17371 6344
rect 17313 6335 17371 6341
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 22094 6381 22100 6384
rect 19076 6344 21864 6372
rect 19076 6316 19104 6344
rect 15194 6313 15200 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14200 6276 14933 6304
rect 14200 6248 14228 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 15188 6267 15200 6313
rect 15194 6264 15200 6267
rect 15252 6264 15258 6316
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17460 6276 17509 6304
rect 17460 6264 17466 6276
rect 17497 6273 17509 6276
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17586 6264 17592 6316
rect 17644 6264 17650 6316
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18564 6276 18797 6304
rect 18564 6264 18570 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19058 6264 19064 6316
rect 19116 6264 19122 6316
rect 19328 6307 19386 6313
rect 19328 6273 19340 6307
rect 19374 6304 19386 6307
rect 19610 6304 19616 6316
rect 19374 6276 19616 6304
rect 19374 6273 19386 6276
rect 19328 6267 19386 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21726 6304 21732 6316
rect 20947 6276 21732 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 21836 6313 21864 6344
rect 22088 6335 22100 6381
rect 22152 6372 22158 6384
rect 25032 6375 25090 6381
rect 22152 6344 22188 6372
rect 22094 6332 22100 6335
rect 22152 6332 22158 6344
rect 25032 6341 25044 6375
rect 25078 6372 25090 6375
rect 29086 6372 29092 6384
rect 25078 6344 29092 6372
rect 25078 6341 25090 6344
rect 25032 6335 25090 6341
rect 29086 6332 29092 6344
rect 29144 6332 29150 6384
rect 31496 6372 31524 6403
rect 34882 6400 34888 6452
rect 34940 6440 34946 6452
rect 35069 6443 35127 6449
rect 35069 6440 35081 6443
rect 34940 6412 35081 6440
rect 34940 6400 34946 6412
rect 35069 6409 35081 6412
rect 35115 6409 35127 6443
rect 35069 6403 35127 6409
rect 36170 6400 36176 6452
rect 36228 6440 36234 6452
rect 36817 6443 36875 6449
rect 36817 6440 36829 6443
rect 36228 6412 36829 6440
rect 36228 6400 36234 6412
rect 36817 6409 36829 6412
rect 36863 6409 36875 6443
rect 36817 6403 36875 6409
rect 37737 6443 37795 6449
rect 37737 6409 37749 6443
rect 37783 6440 37795 6443
rect 37826 6440 37832 6452
rect 37783 6412 37832 6440
rect 37783 6409 37795 6412
rect 37737 6403 37795 6409
rect 31846 6372 31852 6384
rect 31496 6344 31852 6372
rect 31846 6332 31852 6344
rect 31904 6332 31910 6384
rect 32214 6332 32220 6384
rect 32272 6372 32278 6384
rect 34900 6372 34928 6400
rect 32272 6344 34928 6372
rect 36832 6372 36860 6403
rect 37826 6400 37832 6412
rect 37884 6440 37890 6452
rect 38470 6440 38476 6452
rect 37884 6412 38476 6440
rect 37884 6400 37890 6412
rect 38470 6400 38476 6412
rect 38528 6400 38534 6452
rect 38626 6412 40080 6440
rect 38626 6372 38654 6412
rect 36832 6344 38654 6372
rect 39408 6344 39988 6372
rect 32272 6332 32278 6344
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 14182 6196 14188 6248
rect 14240 6196 14246 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 14424 6208 14749 6236
rect 14424 6196 14430 6208
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 17037 6239 17095 6245
rect 17037 6205 17049 6239
rect 17083 6236 17095 6239
rect 17604 6236 17632 6264
rect 17083 6208 17632 6236
rect 17083 6205 17095 6208
rect 17037 6199 17095 6205
rect 12400 6140 13032 6168
rect 12400 6128 12406 6140
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 4062 6060 4068 6112
rect 4120 6060 4126 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4396 6072 4537 6100
rect 4396 6060 4402 6072
rect 4525 6069 4537 6072
rect 4571 6069 4583 6103
rect 5460 6100 5488 6128
rect 14752 6112 14780 6199
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 21174 6196 21180 6248
rect 21232 6196 21238 6248
rect 18892 6168 18920 6196
rect 15856 6140 18920 6168
rect 20441 6171 20499 6177
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5460 6072 5733 6100
rect 4525 6063 4583 6069
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6733 6103 6791 6109
rect 6733 6100 6745 6103
rect 6236 6072 6745 6100
rect 6236 6060 6242 6072
rect 6733 6069 6745 6072
rect 6779 6069 6791 6103
rect 6733 6063 6791 6069
rect 6917 6103 6975 6109
rect 6917 6069 6929 6103
rect 6963 6100 6975 6103
rect 9122 6100 9128 6112
rect 6963 6072 9128 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 13633 6103 13691 6109
rect 13633 6069 13645 6103
rect 13679 6100 13691 6103
rect 13998 6100 14004 6112
rect 13679 6072 14004 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 15856 6100 15884 6140
rect 20441 6137 20453 6171
rect 20487 6168 20499 6171
rect 20714 6168 20720 6180
rect 20487 6140 20720 6168
rect 20487 6137 20499 6140
rect 20441 6131 20499 6137
rect 20714 6128 20720 6140
rect 20772 6128 20778 6180
rect 14792 6072 15884 6100
rect 16301 6103 16359 6109
rect 14792 6060 14798 6072
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 17034 6100 17040 6112
rect 16347 6072 17040 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18230 6060 18236 6112
rect 18288 6060 18294 6112
rect 20530 6060 20536 6112
rect 20588 6060 20594 6112
rect 21836 6100 21864 6267
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 23845 6307 23903 6313
rect 23845 6304 23857 6307
rect 23348 6276 23857 6304
rect 23348 6264 23354 6276
rect 23845 6273 23857 6276
rect 23891 6273 23903 6307
rect 23845 6267 23903 6273
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 27522 6304 27528 6316
rect 26568 6276 27528 6304
rect 26568 6264 26574 6276
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 28813 6307 28871 6313
rect 28813 6273 28825 6307
rect 28859 6304 28871 6307
rect 30466 6304 30472 6316
rect 28859 6276 30472 6304
rect 28859 6273 28871 6276
rect 28813 6267 28871 6273
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31202 6304 31208 6316
rect 31159 6276 31208 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31202 6264 31208 6276
rect 31260 6304 31266 6316
rect 32306 6304 32312 6316
rect 31260 6276 32312 6304
rect 31260 6264 31266 6276
rect 32306 6264 32312 6276
rect 32364 6264 32370 6316
rect 32416 6313 32444 6344
rect 32401 6307 32459 6313
rect 32401 6273 32413 6307
rect 32447 6273 32459 6307
rect 32401 6267 32459 6273
rect 32490 6264 32496 6316
rect 32548 6304 32554 6316
rect 32657 6307 32715 6313
rect 32657 6304 32669 6307
rect 32548 6276 32669 6304
rect 32548 6264 32554 6276
rect 32657 6273 32669 6276
rect 32703 6273 32715 6307
rect 32657 6267 32715 6273
rect 34517 6307 34575 6313
rect 34517 6273 34529 6307
rect 34563 6304 34575 6307
rect 34606 6304 34612 6316
rect 34563 6276 34612 6304
rect 34563 6273 34575 6276
rect 34517 6267 34575 6273
rect 34606 6264 34612 6276
rect 34664 6264 34670 6316
rect 36541 6307 36599 6313
rect 36541 6273 36553 6307
rect 36587 6304 36599 6307
rect 36722 6304 36728 6316
rect 36587 6276 36728 6304
rect 36587 6273 36599 6276
rect 36541 6267 36599 6273
rect 36722 6264 36728 6276
rect 36780 6264 36786 6316
rect 37182 6264 37188 6316
rect 37240 6304 37246 6316
rect 37645 6307 37703 6313
rect 37645 6304 37657 6307
rect 37240 6276 37657 6304
rect 37240 6264 37246 6276
rect 37645 6273 37657 6276
rect 37691 6304 37703 6307
rect 38102 6304 38108 6316
rect 37691 6276 38108 6304
rect 37691 6273 37703 6276
rect 37645 6267 37703 6273
rect 38102 6264 38108 6276
rect 38160 6264 38166 6316
rect 38838 6264 38844 6316
rect 38896 6264 38902 6316
rect 39408 6313 39436 6344
rect 39960 6316 39988 6344
rect 39666 6313 39672 6316
rect 39393 6307 39451 6313
rect 39393 6273 39405 6307
rect 39439 6273 39451 6307
rect 39393 6267 39451 6273
rect 39660 6267 39672 6313
rect 39666 6264 39672 6267
rect 39724 6264 39730 6316
rect 39942 6264 39948 6316
rect 40000 6264 40006 6316
rect 40052 6304 40080 6412
rect 40402 6400 40408 6452
rect 40460 6440 40466 6452
rect 41509 6443 41567 6449
rect 41509 6440 41521 6443
rect 40460 6412 41521 6440
rect 40460 6400 40466 6412
rect 41509 6409 41521 6412
rect 41555 6440 41567 6443
rect 41966 6440 41972 6452
rect 41555 6412 41972 6440
rect 41555 6409 41567 6412
rect 41509 6403 41567 6409
rect 41966 6400 41972 6412
rect 42024 6400 42030 6452
rect 47394 6400 47400 6452
rect 47452 6400 47458 6452
rect 47581 6443 47639 6449
rect 47581 6409 47593 6443
rect 47627 6440 47639 6443
rect 48406 6440 48412 6452
rect 47627 6412 48412 6440
rect 47627 6409 47639 6412
rect 47581 6403 47639 6409
rect 48406 6400 48412 6412
rect 48464 6400 48470 6452
rect 51905 6443 51963 6449
rect 49160 6412 51856 6440
rect 40126 6332 40132 6384
rect 40184 6372 40190 6384
rect 42426 6372 42432 6384
rect 40184 6344 42432 6372
rect 40184 6332 40190 6344
rect 42426 6332 42432 6344
rect 42484 6332 42490 6384
rect 44542 6372 44548 6384
rect 42536 6344 44548 6372
rect 41693 6307 41751 6313
rect 40052 6276 41644 6304
rect 23198 6196 23204 6248
rect 23256 6236 23262 6248
rect 24397 6239 24455 6245
rect 24397 6236 24409 6239
rect 23256 6208 24409 6236
rect 23256 6196 23262 6208
rect 24397 6205 24409 6208
rect 24443 6205 24455 6239
rect 24397 6199 24455 6205
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 24765 6239 24823 6245
rect 24765 6236 24777 6239
rect 24728 6208 24777 6236
rect 24728 6196 24734 6208
rect 24765 6205 24777 6208
rect 24811 6205 24823 6239
rect 24765 6199 24823 6205
rect 27617 6239 27675 6245
rect 27617 6205 27629 6239
rect 27663 6205 27675 6239
rect 27617 6199 27675 6205
rect 30929 6239 30987 6245
rect 30929 6205 30941 6239
rect 30975 6205 30987 6239
rect 31754 6236 31760 6248
rect 30929 6199 30987 6205
rect 26145 6171 26203 6177
rect 26145 6137 26157 6171
rect 26191 6168 26203 6171
rect 27632 6168 27660 6199
rect 26191 6140 27660 6168
rect 30944 6168 30972 6199
rect 31726 6196 31760 6236
rect 31812 6196 31818 6248
rect 37829 6239 37887 6245
rect 37829 6236 37841 6239
rect 33704 6208 37841 6236
rect 31726 6168 31754 6196
rect 30944 6140 31754 6168
rect 26191 6137 26203 6140
rect 26145 6131 26203 6137
rect 22186 6100 22192 6112
rect 21836 6072 22192 6100
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 23290 6060 23296 6112
rect 23348 6060 23354 6112
rect 31726 6100 31754 6140
rect 33704 6100 33732 6208
rect 37829 6205 37841 6208
rect 37875 6236 37887 6239
rect 40865 6239 40923 6245
rect 40865 6236 40877 6239
rect 37875 6208 38654 6236
rect 37875 6205 37887 6208
rect 37829 6199 37887 6205
rect 33781 6171 33839 6177
rect 33781 6137 33793 6171
rect 33827 6168 33839 6171
rect 34514 6168 34520 6180
rect 33827 6140 34520 6168
rect 33827 6137 33839 6140
rect 33781 6131 33839 6137
rect 34514 6128 34520 6140
rect 34572 6128 34578 6180
rect 31726 6072 33732 6100
rect 33870 6060 33876 6112
rect 33928 6060 33934 6112
rect 37277 6103 37335 6109
rect 37277 6069 37289 6103
rect 37323 6100 37335 6103
rect 37458 6100 37464 6112
rect 37323 6072 37464 6100
rect 37323 6069 37335 6072
rect 37277 6063 37335 6069
rect 37458 6060 37464 6072
rect 37516 6060 37522 6112
rect 38286 6060 38292 6112
rect 38344 6060 38350 6112
rect 38626 6100 38654 6208
rect 40788 6208 40877 6236
rect 40788 6177 40816 6208
rect 40865 6205 40877 6208
rect 40911 6205 40923 6239
rect 41616 6236 41644 6276
rect 41693 6273 41705 6307
rect 41739 6304 41751 6307
rect 41782 6304 41788 6316
rect 41739 6276 41788 6304
rect 41739 6273 41751 6276
rect 41693 6267 41751 6273
rect 41782 6264 41788 6276
rect 41840 6264 41846 6316
rect 42536 6245 42564 6344
rect 44542 6332 44548 6344
rect 44600 6332 44606 6384
rect 46032 6344 49096 6372
rect 42797 6307 42855 6313
rect 42797 6273 42809 6307
rect 42843 6273 42855 6307
rect 42797 6267 42855 6273
rect 42153 6239 42211 6245
rect 42153 6236 42165 6239
rect 41616 6208 42165 6236
rect 40865 6199 40923 6205
rect 42153 6205 42165 6208
rect 42199 6236 42211 6239
rect 42521 6239 42579 6245
rect 42521 6236 42533 6239
rect 42199 6208 42533 6236
rect 42199 6205 42211 6208
rect 42153 6199 42211 6205
rect 42521 6205 42533 6208
rect 42567 6205 42579 6239
rect 42521 6199 42579 6205
rect 42610 6196 42616 6248
rect 42668 6236 42674 6248
rect 42705 6239 42763 6245
rect 42705 6236 42717 6239
rect 42668 6208 42717 6236
rect 42668 6196 42674 6208
rect 42705 6205 42717 6208
rect 42751 6205 42763 6239
rect 42705 6199 42763 6205
rect 40773 6171 40831 6177
rect 40773 6137 40785 6171
rect 40819 6137 40831 6171
rect 40773 6131 40831 6137
rect 41046 6128 41052 6180
rect 41104 6128 41110 6180
rect 41414 6128 41420 6180
rect 41472 6168 41478 6180
rect 41877 6171 41935 6177
rect 41877 6168 41889 6171
rect 41472 6140 41889 6168
rect 41472 6128 41478 6140
rect 41877 6137 41889 6140
rect 41923 6168 41935 6171
rect 42812 6168 42840 6267
rect 45922 6264 45928 6316
rect 45980 6304 45986 6316
rect 46032 6313 46060 6344
rect 46017 6307 46075 6313
rect 46017 6304 46029 6307
rect 45980 6276 46029 6304
rect 45980 6264 45986 6276
rect 46017 6273 46029 6276
rect 46063 6273 46075 6307
rect 46017 6267 46075 6273
rect 46284 6307 46342 6313
rect 46284 6273 46296 6307
rect 46330 6304 46342 6307
rect 46842 6304 46848 6316
rect 46330 6276 46848 6304
rect 46330 6273 46342 6276
rect 46284 6267 46342 6273
rect 46842 6264 46848 6276
rect 46900 6264 46906 6316
rect 47302 6264 47308 6316
rect 47360 6304 47366 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47360 6276 47961 6304
rect 47360 6264 47366 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 48038 6264 48044 6316
rect 48096 6264 48102 6316
rect 49068 6313 49096 6344
rect 49053 6307 49111 6313
rect 49053 6273 49065 6307
rect 49099 6273 49111 6307
rect 49053 6267 49111 6273
rect 43809 6239 43867 6245
rect 43809 6205 43821 6239
rect 43855 6205 43867 6239
rect 43809 6199 43867 6205
rect 41923 6140 42840 6168
rect 43165 6171 43223 6177
rect 41923 6137 41935 6140
rect 41877 6131 41935 6137
rect 43165 6137 43177 6171
rect 43211 6168 43223 6171
rect 43824 6168 43852 6199
rect 47394 6196 47400 6248
rect 47452 6236 47458 6248
rect 48133 6239 48191 6245
rect 48133 6236 48145 6239
rect 47452 6208 48145 6236
rect 47452 6196 47458 6208
rect 48133 6205 48145 6208
rect 48179 6236 48191 6239
rect 49160 6236 49188 6412
rect 50792 6375 50850 6381
rect 50792 6341 50804 6375
rect 50838 6372 50850 6375
rect 50890 6372 50896 6384
rect 50838 6344 50896 6372
rect 50838 6341 50850 6344
rect 50792 6335 50850 6341
rect 50890 6332 50896 6344
rect 50948 6332 50954 6384
rect 49326 6313 49332 6316
rect 49320 6267 49332 6313
rect 49326 6264 49332 6267
rect 49384 6264 49390 6316
rect 50154 6264 50160 6316
rect 50212 6304 50218 6316
rect 50525 6307 50583 6313
rect 50525 6304 50537 6307
rect 50212 6276 50537 6304
rect 50212 6264 50218 6276
rect 50525 6273 50537 6276
rect 50571 6304 50583 6307
rect 51828 6304 51856 6412
rect 51905 6409 51917 6443
rect 51951 6440 51963 6443
rect 52638 6440 52644 6452
rect 51951 6412 52644 6440
rect 51951 6409 51963 6412
rect 51905 6403 51963 6409
rect 52638 6400 52644 6412
rect 52696 6400 52702 6452
rect 55398 6400 55404 6452
rect 55456 6400 55462 6452
rect 56597 6443 56655 6449
rect 56597 6409 56609 6443
rect 56643 6440 56655 6443
rect 56962 6440 56968 6452
rect 56643 6412 56968 6440
rect 56643 6409 56655 6412
rect 56597 6403 56655 6409
rect 56962 6400 56968 6412
rect 57020 6400 57026 6452
rect 57885 6443 57943 6449
rect 57885 6409 57897 6443
rect 57931 6440 57943 6443
rect 58250 6440 58256 6452
rect 57931 6412 58256 6440
rect 57931 6409 57943 6412
rect 57885 6403 57943 6409
rect 52270 6332 52276 6384
rect 52328 6332 52334 6384
rect 51994 6304 52000 6316
rect 50571 6276 51764 6304
rect 51828 6276 52000 6304
rect 50571 6273 50583 6276
rect 50525 6267 50583 6273
rect 48179 6208 49188 6236
rect 51736 6236 51764 6276
rect 51994 6264 52000 6276
rect 52052 6304 52058 6316
rect 55416 6304 55444 6400
rect 56505 6375 56563 6381
rect 56505 6341 56517 6375
rect 56551 6372 56563 6375
rect 57900 6372 57928 6403
rect 58250 6400 58256 6412
rect 58308 6400 58314 6452
rect 56551 6344 57928 6372
rect 56551 6341 56563 6344
rect 56505 6335 56563 6341
rect 52052 6276 55444 6304
rect 52052 6264 52058 6276
rect 54110 6236 54116 6248
rect 51736 6208 54116 6236
rect 48179 6205 48191 6208
rect 48133 6199 48191 6205
rect 54110 6196 54116 6208
rect 54168 6196 54174 6248
rect 55490 6196 55496 6248
rect 55548 6196 55554 6248
rect 56321 6239 56379 6245
rect 56321 6205 56333 6239
rect 56367 6205 56379 6239
rect 56321 6199 56379 6205
rect 57609 6239 57667 6245
rect 57609 6205 57621 6239
rect 57655 6205 57667 6239
rect 57609 6199 57667 6205
rect 58529 6239 58587 6245
rect 58529 6205 58541 6239
rect 58575 6205 58587 6239
rect 58529 6199 58587 6205
rect 56336 6168 56364 6199
rect 43211 6140 43852 6168
rect 55416 6140 56364 6168
rect 56965 6171 57023 6177
rect 43211 6137 43223 6140
rect 43165 6131 43223 6137
rect 39301 6103 39359 6109
rect 39301 6100 39313 6103
rect 38626 6072 39313 6100
rect 39301 6069 39313 6072
rect 39347 6100 39359 6103
rect 41064 6100 41092 6128
rect 55416 6112 55444 6140
rect 56965 6137 56977 6171
rect 57011 6168 57023 6171
rect 57624 6168 57652 6199
rect 57011 6140 57652 6168
rect 57011 6137 57023 6140
rect 56965 6131 57023 6137
rect 39347 6072 41092 6100
rect 39347 6069 39359 6072
rect 39301 6063 39359 6069
rect 43254 6060 43260 6112
rect 43312 6060 43318 6112
rect 50430 6060 50436 6112
rect 50488 6060 50494 6112
rect 50798 6060 50804 6112
rect 50856 6100 50862 6112
rect 54113 6103 54171 6109
rect 54113 6100 54125 6103
rect 50856 6072 54125 6100
rect 50856 6060 50862 6072
rect 54113 6069 54125 6072
rect 54159 6100 54171 6103
rect 54846 6100 54852 6112
rect 54159 6072 54852 6100
rect 54159 6069 54171 6072
rect 54113 6063 54171 6069
rect 54846 6060 54852 6072
rect 54904 6060 54910 6112
rect 54938 6060 54944 6112
rect 54996 6060 55002 6112
rect 55398 6060 55404 6112
rect 55456 6060 55462 6112
rect 56134 6060 56140 6112
rect 56192 6060 56198 6112
rect 57054 6060 57060 6112
rect 57112 6060 57118 6112
rect 58544 6100 58572 6199
rect 58544 6072 58940 6100
rect 1104 6010 58880 6032
rect 1104 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 22616 6010
rect 22668 5958 22680 6010
rect 22732 5958 22744 6010
rect 22796 5958 22808 6010
rect 22860 5958 22872 6010
rect 22924 5958 37060 6010
rect 37112 5958 37124 6010
rect 37176 5958 37188 6010
rect 37240 5958 37252 6010
rect 37304 5958 37316 6010
rect 37368 5958 51504 6010
rect 51556 5958 51568 6010
rect 51620 5958 51632 6010
rect 51684 5958 51696 6010
rect 51748 5958 51760 6010
rect 51812 5958 58880 6010
rect 1104 5936 58880 5958
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 2133 5899 2191 5905
rect 2133 5896 2145 5899
rect 1912 5868 2145 5896
rect 1912 5856 1918 5868
rect 2133 5865 2145 5868
rect 2179 5865 2191 5899
rect 2958 5896 2964 5908
rect 2133 5859 2191 5865
rect 2357 5868 2964 5896
rect 1946 5788 1952 5840
rect 2004 5788 2010 5840
rect 1964 5760 1992 5788
rect 1872 5732 1992 5760
rect 2041 5763 2099 5769
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 1872 5692 1900 5732
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2357 5760 2385 5868
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 5902 5896 5908 5908
rect 3528 5868 5908 5896
rect 3234 5828 3240 5840
rect 3068 5800 3240 5828
rect 3068 5760 3096 5800
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 2087 5732 2385 5760
rect 2608 5732 3096 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 1811 5664 1900 5692
rect 1949 5695 2007 5701
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2608 5692 2636 5732
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 3528 5769 3556 5868
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6086 5856 6092 5908
rect 6144 5856 6150 5908
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 7650 5896 7656 5908
rect 6503 5868 7656 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8754 5896 8760 5908
rect 8435 5868 8760 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 12434 5896 12440 5908
rect 9232 5868 12440 5896
rect 6104 5828 6132 5856
rect 9232 5828 9260 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 13538 5896 13544 5908
rect 12759 5868 13544 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 15565 5899 15623 5905
rect 15565 5896 15577 5899
rect 15344 5868 15577 5896
rect 15344 5856 15350 5868
rect 15565 5865 15577 5868
rect 15611 5865 15623 5899
rect 15565 5859 15623 5865
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16485 5899 16543 5905
rect 16485 5896 16497 5899
rect 16172 5868 16497 5896
rect 16172 5856 16178 5868
rect 16485 5865 16497 5868
rect 16531 5865 16543 5899
rect 16485 5859 16543 5865
rect 17034 5856 17040 5908
rect 17092 5856 17098 5908
rect 17589 5899 17647 5905
rect 17589 5865 17601 5899
rect 17635 5896 17647 5899
rect 17678 5896 17684 5908
rect 17635 5868 17684 5896
rect 17635 5865 17647 5868
rect 17589 5859 17647 5865
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 19981 5899 20039 5905
rect 19981 5896 19993 5899
rect 19668 5868 19993 5896
rect 19668 5856 19674 5868
rect 19981 5865 19993 5868
rect 20027 5865 20039 5899
rect 19981 5859 20039 5865
rect 20530 5856 20536 5908
rect 20588 5856 20594 5908
rect 20714 5856 20720 5908
rect 20772 5856 20778 5908
rect 21361 5899 21419 5905
rect 21361 5865 21373 5899
rect 21407 5896 21419 5899
rect 21726 5896 21732 5908
rect 21407 5868 21732 5896
rect 21407 5865 21419 5868
rect 21361 5859 21419 5865
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 28902 5856 28908 5908
rect 28960 5856 28966 5908
rect 30558 5856 30564 5908
rect 30616 5856 30622 5908
rect 31202 5856 31208 5908
rect 31260 5856 31266 5908
rect 32401 5899 32459 5905
rect 32401 5865 32413 5899
rect 32447 5896 32459 5899
rect 32582 5896 32588 5908
rect 32447 5868 32588 5896
rect 32447 5865 32459 5868
rect 32401 5859 32459 5865
rect 32582 5856 32588 5868
rect 32640 5856 32646 5908
rect 33229 5899 33287 5905
rect 33229 5865 33241 5899
rect 33275 5896 33287 5899
rect 35250 5896 35256 5908
rect 33275 5868 35256 5896
rect 33275 5865 33287 5868
rect 33229 5859 33287 5865
rect 35250 5856 35256 5868
rect 35308 5856 35314 5908
rect 37458 5856 37464 5908
rect 37516 5856 37522 5908
rect 38102 5856 38108 5908
rect 38160 5856 38166 5908
rect 39298 5856 39304 5908
rect 39356 5896 39362 5908
rect 39577 5899 39635 5905
rect 39577 5896 39589 5899
rect 39356 5868 39589 5896
rect 39356 5856 39362 5868
rect 39577 5865 39589 5868
rect 39623 5865 39635 5899
rect 39577 5859 39635 5865
rect 39666 5856 39672 5908
rect 39724 5896 39730 5908
rect 39853 5899 39911 5905
rect 39853 5896 39865 5899
rect 39724 5868 39865 5896
rect 39724 5856 39730 5868
rect 39853 5865 39865 5868
rect 39899 5865 39911 5899
rect 39853 5859 39911 5865
rect 40126 5856 40132 5908
rect 40184 5896 40190 5908
rect 40865 5899 40923 5905
rect 40865 5896 40877 5899
rect 40184 5868 40877 5896
rect 40184 5856 40190 5868
rect 40865 5865 40877 5868
rect 40911 5865 40923 5899
rect 40865 5859 40923 5865
rect 42610 5856 42616 5908
rect 42668 5896 42674 5908
rect 43349 5899 43407 5905
rect 43349 5896 43361 5899
rect 42668 5868 43361 5896
rect 42668 5856 42674 5868
rect 43349 5865 43361 5868
rect 43395 5865 43407 5899
rect 43349 5859 43407 5865
rect 44542 5856 44548 5908
rect 44600 5896 44606 5908
rect 47394 5896 47400 5908
rect 44600 5868 47400 5896
rect 44600 5856 44606 5868
rect 47394 5856 47400 5868
rect 47452 5856 47458 5908
rect 49326 5856 49332 5908
rect 49384 5856 49390 5908
rect 50985 5899 51043 5905
rect 49712 5868 50660 5896
rect 6104 5800 9260 5828
rect 3513 5763 3571 5769
rect 3513 5760 3525 5763
rect 3200 5732 3525 5760
rect 3200 5720 3206 5732
rect 3513 5729 3525 5732
rect 3559 5729 3571 5763
rect 3513 5723 3571 5729
rect 9122 5720 9128 5772
rect 9180 5720 9186 5772
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 14182 5760 14188 5772
rect 12544 5732 14188 5760
rect 1995 5664 2636 5692
rect 2685 5695 2743 5701
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 2700 5624 2728 5655
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4338 5701 4344 5704
rect 4332 5692 4344 5701
rect 4299 5664 4344 5692
rect 4332 5655 4344 5664
rect 4338 5652 4344 5655
rect 4396 5652 4402 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6178 5692 6184 5704
rect 5592 5664 6184 5692
rect 5592 5652 5598 5664
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 9140 5692 9168 5720
rect 8067 5664 9168 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 1627 5596 2728 5624
rect 5460 5624 5488 5652
rect 7116 5624 7144 5655
rect 9214 5652 9220 5704
rect 9272 5652 9278 5704
rect 9876 5692 9904 5720
rect 12544 5704 12572 5732
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 16132 5769 16160 5856
rect 17052 5769 17080 5856
rect 20548 5769 20576 5856
rect 20732 5769 20760 5856
rect 26053 5831 26111 5837
rect 26053 5797 26065 5831
rect 26099 5828 26111 5831
rect 26099 5800 27016 5828
rect 26099 5797 26111 5800
rect 26053 5791 26111 5797
rect 16117 5763 16175 5769
rect 16117 5729 16129 5763
rect 16163 5729 16175 5763
rect 16117 5723 16175 5729
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 17037 5763 17095 5769
rect 16347 5732 16436 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 9876 5664 11345 5692
rect 11333 5661 11345 5664
rect 11379 5692 11391 5695
rect 12526 5692 12532 5704
rect 11379 5664 12532 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 7190 5624 7196 5636
rect 5460 5596 7196 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5624 7619 5627
rect 8757 5627 8815 5633
rect 8757 5624 8769 5627
rect 7607 5596 8769 5624
rect 7607 5593 7619 5596
rect 7561 5587 7619 5593
rect 8757 5593 8769 5596
rect 8803 5624 8815 5627
rect 9950 5624 9956 5636
rect 8803 5596 9956 5624
rect 8803 5593 8815 5596
rect 8757 5587 8815 5593
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 10134 5633 10140 5636
rect 10128 5624 10140 5633
rect 10095 5596 10140 5624
rect 10128 5587 10140 5596
rect 10134 5584 10140 5587
rect 10192 5584 10198 5636
rect 11600 5627 11658 5633
rect 11600 5593 11612 5627
rect 11646 5624 11658 5627
rect 12897 5627 12955 5633
rect 12897 5624 12909 5627
rect 11646 5596 12909 5624
rect 11646 5593 11658 5596
rect 11600 5587 11658 5593
rect 12897 5593 12909 5596
rect 12943 5593 12955 5627
rect 13556 5624 13584 5655
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14441 5695 14499 5701
rect 14441 5692 14453 5695
rect 13964 5664 14453 5692
rect 13964 5652 13970 5664
rect 14441 5661 14453 5664
rect 14487 5661 14499 5695
rect 14441 5655 14499 5661
rect 16022 5652 16028 5704
rect 16080 5652 16086 5704
rect 14090 5624 14096 5636
rect 13556 5596 14096 5624
rect 12897 5587 12955 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 15930 5624 15936 5636
rect 15580 5596 15936 5624
rect 4522 5516 4528 5568
rect 4580 5556 4586 5568
rect 5258 5556 5264 5568
rect 4580 5528 5264 5556
rect 4580 5516 4586 5528
rect 5258 5516 5264 5528
rect 5316 5556 5322 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 5316 5528 5457 5556
rect 5316 5516 5322 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 11238 5516 11244 5568
rect 11296 5516 11302 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 13998 5556 14004 5568
rect 13955 5528 14004 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 13998 5516 14004 5528
rect 14056 5556 14062 5568
rect 15580 5556 15608 5596
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 16408 5624 16436 5732
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 20533 5763 20591 5769
rect 20533 5729 20545 5763
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5729 20775 5763
rect 23201 5763 23259 5769
rect 23201 5760 23213 5763
rect 20717 5723 20775 5729
rect 22756 5732 23213 5760
rect 17954 5652 17960 5704
rect 18012 5692 18018 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 18012 5664 18245 5692
rect 18012 5652 18018 5664
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 22756 5692 22784 5732
rect 23201 5729 23213 5732
rect 23247 5760 23259 5763
rect 23474 5760 23480 5772
rect 23247 5732 23480 5760
rect 23247 5729 23259 5732
rect 23201 5723 23259 5729
rect 23474 5720 23480 5732
rect 23532 5720 23538 5772
rect 24670 5720 24676 5772
rect 24728 5720 24734 5772
rect 26602 5760 26608 5772
rect 25700 5732 26608 5760
rect 18233 5655 18291 5661
rect 19306 5664 22784 5692
rect 19306 5624 19334 5664
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 25700 5692 25728 5732
rect 26602 5720 26608 5732
rect 26660 5760 26666 5772
rect 26697 5763 26755 5769
rect 26697 5760 26709 5763
rect 26660 5732 26709 5760
rect 26660 5720 26666 5732
rect 26697 5729 26709 5732
rect 26743 5760 26755 5763
rect 26878 5760 26884 5772
rect 26743 5732 26884 5760
rect 26743 5729 26755 5732
rect 26697 5723 26755 5729
rect 26878 5720 26884 5732
rect 26936 5720 26942 5772
rect 26988 5769 27016 5800
rect 26973 5763 27031 5769
rect 26973 5729 26985 5763
rect 27019 5729 27031 5763
rect 26973 5723 27031 5729
rect 28626 5720 28632 5772
rect 28684 5720 28690 5772
rect 28920 5760 28948 5856
rect 30576 5769 30604 5856
rect 31110 5788 31116 5840
rect 31168 5828 31174 5840
rect 34977 5831 35035 5837
rect 31168 5800 33916 5828
rect 31168 5788 31174 5800
rect 30101 5763 30159 5769
rect 30101 5760 30113 5763
rect 28920 5732 30113 5760
rect 30101 5729 30113 5732
rect 30147 5729 30159 5763
rect 30101 5723 30159 5729
rect 30561 5763 30619 5769
rect 30561 5729 30573 5763
rect 30607 5729 30619 5763
rect 30561 5723 30619 5729
rect 32033 5763 32091 5769
rect 32033 5729 32045 5763
rect 32079 5760 32091 5763
rect 32585 5763 32643 5769
rect 32585 5760 32597 5763
rect 32079 5732 32597 5760
rect 32079 5729 32091 5732
rect 32033 5723 32091 5729
rect 32585 5729 32597 5732
rect 32631 5760 32643 5763
rect 33226 5760 33232 5772
rect 32631 5732 33232 5760
rect 32631 5729 32643 5732
rect 32585 5723 32643 5729
rect 33226 5720 33232 5732
rect 33284 5720 33290 5772
rect 33318 5720 33324 5772
rect 33376 5760 33382 5772
rect 33778 5760 33784 5772
rect 33376 5732 33784 5760
rect 33376 5720 33382 5732
rect 33778 5720 33784 5732
rect 33836 5720 33842 5772
rect 33888 5769 33916 5800
rect 34977 5797 34989 5831
rect 35023 5828 35035 5831
rect 35066 5828 35072 5840
rect 35023 5800 35072 5828
rect 35023 5797 35035 5800
rect 34977 5791 35035 5797
rect 35066 5788 35072 5800
rect 35124 5788 35130 5840
rect 36633 5831 36691 5837
rect 36633 5797 36645 5831
rect 36679 5797 36691 5831
rect 36633 5791 36691 5797
rect 33873 5763 33931 5769
rect 33873 5729 33885 5763
rect 33919 5760 33931 5763
rect 34698 5760 34704 5772
rect 33919 5732 34704 5760
rect 33919 5729 33931 5732
rect 33873 5723 33931 5729
rect 34698 5720 34704 5732
rect 34756 5720 34762 5772
rect 34882 5720 34888 5772
rect 34940 5760 34946 5772
rect 35253 5763 35311 5769
rect 35253 5760 35265 5763
rect 34940 5732 35265 5760
rect 34940 5720 34946 5732
rect 35253 5729 35265 5732
rect 35299 5729 35311 5763
rect 35253 5723 35311 5729
rect 24872 5664 25728 5692
rect 26513 5695 26571 5701
rect 24872 5624 24900 5664
rect 26513 5661 26525 5695
rect 26559 5692 26571 5695
rect 27154 5692 27160 5704
rect 26559 5664 27160 5692
rect 26559 5661 26571 5664
rect 26513 5655 26571 5661
rect 27154 5652 27160 5664
rect 27212 5692 27218 5704
rect 27617 5695 27675 5701
rect 27617 5692 27629 5695
rect 27212 5664 27629 5692
rect 27212 5652 27218 5664
rect 27617 5661 27629 5664
rect 27663 5661 27675 5695
rect 27617 5655 27675 5661
rect 15988 5596 19334 5624
rect 22112 5596 24900 5624
rect 24940 5627 24998 5633
rect 15988 5584 15994 5596
rect 14056 5528 15608 5556
rect 15657 5559 15715 5565
rect 14056 5516 14062 5528
rect 15657 5525 15669 5559
rect 15703 5556 15715 5559
rect 15838 5556 15844 5568
rect 15703 5528 15844 5556
rect 15703 5525 15715 5528
rect 15657 5519 15715 5525
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 17678 5516 17684 5568
rect 17736 5516 17742 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 19392 5528 19441 5556
rect 19392 5516 19398 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 22112 5556 22140 5596
rect 24940 5593 24952 5627
rect 24986 5624 24998 5627
rect 25590 5624 25596 5636
rect 24986 5596 25596 5624
rect 24986 5593 24998 5596
rect 24940 5587 24998 5593
rect 25590 5584 25596 5596
rect 25648 5584 25654 5636
rect 26605 5627 26663 5633
rect 26605 5593 26617 5627
rect 26651 5624 26663 5627
rect 28644 5624 28672 5720
rect 28810 5652 28816 5704
rect 28868 5652 28874 5704
rect 32861 5695 32919 5701
rect 32861 5661 32873 5695
rect 32907 5692 32919 5695
rect 33134 5692 33140 5704
rect 32907 5664 33140 5692
rect 32907 5661 32919 5664
rect 32861 5655 32919 5661
rect 33134 5652 33140 5664
rect 33192 5652 33198 5704
rect 33689 5695 33747 5701
rect 33689 5661 33701 5695
rect 33735 5692 33747 5695
rect 33962 5692 33968 5704
rect 33735 5664 33968 5692
rect 33735 5661 33747 5664
rect 33689 5655 33747 5661
rect 26651 5596 28672 5624
rect 26651 5593 26663 5596
rect 26605 5587 26663 5593
rect 30650 5584 30656 5636
rect 30708 5624 30714 5636
rect 32769 5627 32827 5633
rect 32769 5624 32781 5627
rect 30708 5596 32781 5624
rect 30708 5584 30714 5596
rect 32769 5593 32781 5596
rect 32815 5624 32827 5627
rect 33704 5624 33732 5655
rect 33962 5652 33968 5664
rect 34020 5652 34026 5704
rect 36648 5692 36676 5791
rect 37369 5763 37427 5769
rect 37369 5729 37381 5763
rect 37415 5760 37427 5763
rect 37476 5760 37504 5856
rect 49712 5840 49740 5868
rect 37642 5788 37648 5840
rect 37700 5828 37706 5840
rect 41233 5831 41291 5837
rect 41233 5828 41245 5831
rect 37700 5800 41245 5828
rect 37700 5788 37706 5800
rect 41233 5797 41245 5800
rect 41279 5828 41291 5831
rect 41690 5828 41696 5840
rect 41279 5800 41696 5828
rect 41279 5797 41291 5800
rect 41233 5791 41291 5797
rect 41690 5788 41696 5800
rect 41748 5788 41754 5840
rect 43257 5831 43315 5837
rect 43257 5797 43269 5831
rect 43303 5797 43315 5831
rect 43257 5791 43315 5797
rect 37415 5732 37504 5760
rect 37415 5729 37427 5732
rect 37369 5723 37427 5729
rect 37461 5695 37519 5701
rect 37461 5692 37473 5695
rect 36648 5664 37473 5692
rect 37461 5661 37473 5664
rect 37507 5661 37519 5695
rect 37461 5655 37519 5661
rect 32815 5596 33732 5624
rect 35520 5627 35578 5633
rect 32815 5593 32827 5596
rect 32769 5587 32827 5593
rect 35520 5593 35532 5627
rect 35566 5624 35578 5627
rect 36725 5627 36783 5633
rect 36725 5624 36737 5627
rect 35566 5596 36737 5624
rect 35566 5593 35578 5596
rect 35520 5587 35578 5593
rect 36725 5593 36737 5596
rect 36771 5593 36783 5627
rect 36725 5587 36783 5593
rect 36814 5584 36820 5636
rect 36872 5624 36878 5636
rect 37660 5624 37688 5788
rect 41506 5720 41512 5772
rect 41564 5720 41570 5772
rect 43272 5760 43300 5791
rect 46290 5788 46296 5840
rect 46348 5828 46354 5840
rect 49694 5828 49700 5840
rect 46348 5800 49700 5828
rect 46348 5788 46354 5800
rect 49694 5788 49700 5800
rect 49752 5788 49758 5840
rect 50157 5831 50215 5837
rect 50157 5828 50169 5831
rect 49988 5800 50169 5828
rect 49988 5769 50016 5800
rect 50157 5797 50169 5800
rect 50203 5797 50215 5831
rect 50632 5828 50660 5868
rect 50985 5865 50997 5899
rect 51031 5896 51043 5899
rect 51258 5896 51264 5908
rect 51031 5868 51264 5896
rect 51031 5865 51043 5868
rect 50985 5859 51043 5865
rect 51258 5856 51264 5868
rect 51316 5856 51322 5908
rect 55122 5856 55128 5908
rect 55180 5856 55186 5908
rect 58161 5899 58219 5905
rect 58161 5865 58173 5899
rect 58207 5896 58219 5899
rect 58912 5896 58940 6072
rect 58207 5868 58940 5896
rect 58207 5865 58219 5868
rect 58161 5859 58219 5865
rect 50798 5828 50804 5840
rect 50632 5800 50804 5828
rect 50157 5791 50215 5797
rect 43901 5763 43959 5769
rect 43901 5760 43913 5763
rect 43272 5732 43913 5760
rect 43901 5729 43913 5732
rect 43947 5729 43959 5763
rect 46845 5763 46903 5769
rect 46845 5760 46857 5763
rect 43901 5723 43959 5729
rect 45480 5732 46857 5760
rect 38654 5652 38660 5704
rect 38712 5692 38718 5704
rect 38749 5695 38807 5701
rect 38749 5692 38761 5695
rect 38712 5664 38761 5692
rect 38712 5652 38718 5664
rect 38749 5661 38761 5664
rect 38795 5661 38807 5695
rect 38749 5655 38807 5661
rect 40034 5652 40040 5704
rect 40092 5692 40098 5704
rect 40405 5695 40463 5701
rect 40405 5692 40417 5695
rect 40092 5664 40417 5692
rect 40092 5652 40098 5664
rect 40405 5661 40417 5664
rect 40451 5661 40463 5695
rect 41524 5692 41552 5720
rect 45480 5704 45508 5732
rect 46845 5729 46857 5732
rect 46891 5729 46903 5763
rect 46845 5723 46903 5729
rect 49973 5763 50031 5769
rect 49973 5729 49985 5763
rect 50019 5729 50031 5763
rect 50614 5760 50620 5772
rect 49973 5723 50031 5729
rect 50448 5732 50620 5760
rect 41877 5695 41935 5701
rect 41877 5692 41889 5695
rect 41524 5664 41889 5692
rect 40405 5655 40463 5661
rect 41877 5661 41889 5664
rect 41923 5661 41935 5695
rect 41877 5655 41935 5661
rect 43254 5652 43260 5704
rect 43312 5652 43318 5704
rect 45189 5695 45247 5701
rect 45189 5692 45201 5695
rect 43364 5664 45201 5692
rect 36872 5596 37688 5624
rect 42144 5627 42202 5633
rect 36872 5584 36878 5596
rect 42144 5593 42156 5627
rect 42190 5624 42202 5627
rect 43272 5624 43300 5652
rect 42190 5596 43300 5624
rect 42190 5593 42202 5596
rect 42144 5587 42202 5593
rect 20404 5528 22140 5556
rect 20404 5516 20410 5528
rect 22186 5516 22192 5568
rect 22244 5556 22250 5568
rect 22281 5559 22339 5565
rect 22281 5556 22293 5559
rect 22244 5528 22293 5556
rect 22244 5516 22250 5528
rect 22281 5525 22293 5528
rect 22327 5525 22339 5559
rect 22281 5519 22339 5525
rect 26145 5559 26203 5565
rect 26145 5525 26157 5559
rect 26191 5556 26203 5559
rect 26234 5556 26240 5568
rect 26191 5528 26240 5556
rect 26191 5525 26203 5528
rect 26145 5519 26203 5525
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 28258 5516 28264 5568
rect 28316 5516 28322 5568
rect 29546 5516 29552 5568
rect 29604 5516 29610 5568
rect 33318 5516 33324 5568
rect 33376 5516 33382 5568
rect 33410 5516 33416 5568
rect 33468 5556 33474 5568
rect 34425 5559 34483 5565
rect 34425 5556 34437 5559
rect 33468 5528 34437 5556
rect 33468 5516 33474 5528
rect 34425 5525 34437 5528
rect 34471 5556 34483 5559
rect 36832 5556 36860 5584
rect 34471 5528 36860 5556
rect 34471 5525 34483 5528
rect 34425 5519 34483 5525
rect 38194 5516 38200 5568
rect 38252 5516 38258 5568
rect 39114 5516 39120 5568
rect 39172 5516 39178 5568
rect 41690 5516 41696 5568
rect 41748 5556 41754 5568
rect 42702 5556 42708 5568
rect 41748 5528 42708 5556
rect 41748 5516 41754 5528
rect 42702 5516 42708 5528
rect 42760 5516 42766 5568
rect 42978 5516 42984 5568
rect 43036 5556 43042 5568
rect 43364 5556 43392 5664
rect 45189 5661 45201 5664
rect 45235 5692 45247 5695
rect 45462 5692 45468 5704
rect 45235 5664 45468 5692
rect 45235 5661 45247 5664
rect 45189 5655 45247 5661
rect 45462 5652 45468 5664
rect 45520 5652 45526 5704
rect 46106 5652 46112 5704
rect 46164 5652 46170 5704
rect 46198 5652 46204 5704
rect 46256 5692 46262 5704
rect 46477 5695 46535 5701
rect 46477 5692 46489 5695
rect 46256 5664 46489 5692
rect 46256 5652 46262 5664
rect 46477 5661 46489 5664
rect 46523 5661 46535 5695
rect 46477 5655 46535 5661
rect 44174 5584 44180 5636
rect 44232 5624 44238 5636
rect 44361 5627 44419 5633
rect 44361 5624 44373 5627
rect 44232 5596 44373 5624
rect 44232 5584 44238 5596
rect 44361 5593 44373 5596
rect 44407 5624 44419 5627
rect 50448 5624 50476 5732
rect 50614 5720 50620 5732
rect 50672 5720 50678 5772
rect 50724 5769 50752 5800
rect 50798 5788 50804 5800
rect 50856 5788 50862 5840
rect 52178 5828 52184 5840
rect 51460 5800 52184 5828
rect 51460 5769 51488 5800
rect 52178 5788 52184 5800
rect 52236 5788 52242 5840
rect 58342 5788 58348 5840
rect 58400 5788 58406 5840
rect 50709 5763 50767 5769
rect 50709 5729 50721 5763
rect 50755 5729 50767 5763
rect 50709 5723 50767 5729
rect 51445 5763 51503 5769
rect 51445 5729 51457 5763
rect 51491 5729 51503 5763
rect 51445 5723 51503 5729
rect 51626 5720 51632 5772
rect 51684 5760 51690 5772
rect 51994 5760 52000 5772
rect 51684 5732 52000 5760
rect 51684 5720 51690 5732
rect 51994 5720 52000 5732
rect 52052 5720 52058 5772
rect 50525 5695 50583 5701
rect 50525 5661 50537 5695
rect 50571 5692 50583 5695
rect 51350 5692 51356 5704
rect 50571 5664 51356 5692
rect 50571 5661 50583 5664
rect 50525 5655 50583 5661
rect 51350 5652 51356 5664
rect 51408 5652 51414 5704
rect 52730 5652 52736 5704
rect 52788 5692 52794 5704
rect 53193 5695 53251 5701
rect 53193 5692 53205 5695
rect 52788 5664 53205 5692
rect 52788 5652 52794 5664
rect 53193 5661 53205 5664
rect 53239 5661 53251 5695
rect 53193 5655 53251 5661
rect 55309 5695 55367 5701
rect 55309 5661 55321 5695
rect 55355 5692 55367 5695
rect 56318 5692 56324 5704
rect 55355 5664 56324 5692
rect 55355 5661 55367 5664
rect 55309 5655 55367 5661
rect 56318 5652 56324 5664
rect 56376 5692 56382 5704
rect 57054 5701 57060 5704
rect 56781 5695 56839 5701
rect 56781 5692 56793 5695
rect 56376 5664 56793 5692
rect 56376 5652 56382 5664
rect 56781 5661 56793 5664
rect 56827 5661 56839 5695
rect 57048 5692 57060 5701
rect 57015 5664 57060 5692
rect 56781 5655 56839 5661
rect 57048 5655 57060 5664
rect 57054 5652 57060 5655
rect 57112 5652 57118 5704
rect 58526 5652 58532 5704
rect 58584 5652 58590 5704
rect 55576 5627 55634 5633
rect 44407 5596 46336 5624
rect 50448 5596 52868 5624
rect 44407 5593 44419 5596
rect 44361 5587 44419 5593
rect 46308 5568 46336 5596
rect 43036 5528 43392 5556
rect 43036 5516 43042 5528
rect 44634 5516 44640 5568
rect 44692 5516 44698 5568
rect 45554 5516 45560 5568
rect 45612 5516 45618 5568
rect 46290 5516 46296 5568
rect 46348 5516 46354 5568
rect 51368 5565 51396 5596
rect 52840 5568 52868 5596
rect 55576 5593 55588 5627
rect 55622 5624 55634 5627
rect 56134 5624 56140 5636
rect 55622 5596 56140 5624
rect 55622 5593 55634 5596
rect 55576 5587 55634 5593
rect 56134 5584 56140 5596
rect 56192 5584 56198 5636
rect 56244 5596 57284 5624
rect 51353 5559 51411 5565
rect 51353 5525 51365 5559
rect 51399 5525 51411 5559
rect 51353 5519 51411 5525
rect 51994 5516 52000 5568
rect 52052 5556 52058 5568
rect 52181 5559 52239 5565
rect 52181 5556 52193 5559
rect 52052 5528 52193 5556
rect 52052 5516 52058 5528
rect 52181 5525 52193 5528
rect 52227 5525 52239 5559
rect 52181 5519 52239 5525
rect 52638 5516 52644 5568
rect 52696 5516 52702 5568
rect 52822 5516 52828 5568
rect 52880 5516 52886 5568
rect 54662 5516 54668 5568
rect 54720 5556 54726 5568
rect 54757 5559 54815 5565
rect 54757 5556 54769 5559
rect 54720 5528 54769 5556
rect 54720 5516 54726 5528
rect 54757 5525 54769 5528
rect 54803 5556 54815 5559
rect 56244 5556 56272 5596
rect 57256 5568 57284 5596
rect 54803 5528 56272 5556
rect 54803 5525 54815 5528
rect 54757 5519 54815 5525
rect 56686 5516 56692 5568
rect 56744 5516 56750 5568
rect 57238 5516 57244 5568
rect 57296 5516 57302 5568
rect 1104 5466 59040 5488
rect 1104 5414 15394 5466
rect 15446 5414 15458 5466
rect 15510 5414 15522 5466
rect 15574 5414 15586 5466
rect 15638 5414 15650 5466
rect 15702 5414 29838 5466
rect 29890 5414 29902 5466
rect 29954 5414 29966 5466
rect 30018 5414 30030 5466
rect 30082 5414 30094 5466
rect 30146 5414 44282 5466
rect 44334 5414 44346 5466
rect 44398 5414 44410 5466
rect 44462 5414 44474 5466
rect 44526 5414 44538 5466
rect 44590 5414 58726 5466
rect 58778 5414 58790 5466
rect 58842 5414 58854 5466
rect 58906 5414 58918 5466
rect 58970 5414 58982 5466
rect 59034 5414 59040 5466
rect 1104 5392 59040 5414
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3421 5355 3479 5361
rect 3421 5352 3433 5355
rect 3292 5324 3433 5352
rect 3292 5312 3298 5324
rect 3421 5321 3433 5324
rect 3467 5321 3479 5355
rect 3584 5355 3642 5361
rect 3584 5352 3596 5355
rect 3421 5315 3479 5321
rect 3528 5324 3596 5352
rect 2958 5244 2964 5296
rect 3016 5244 3022 5296
rect 3528 5228 3556 5324
rect 3584 5321 3596 5324
rect 3630 5321 3642 5355
rect 3584 5315 3642 5321
rect 3878 5312 3884 5364
rect 3936 5312 3942 5364
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 5626 5352 5632 5364
rect 4488 5324 5632 5352
rect 4488 5312 4494 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 12250 5352 12256 5364
rect 12207 5324 12256 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 22002 5352 22008 5364
rect 12406 5324 22008 5352
rect 3786 5244 3792 5296
rect 3844 5244 3850 5296
rect 5534 5284 5540 5296
rect 4448 5256 5540 5284
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 4448 5216 4476 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 7650 5244 7656 5296
rect 7708 5244 7714 5296
rect 9309 5287 9367 5293
rect 7852 5256 9260 5284
rect 3568 5188 4476 5216
rect 3568 5176 3574 5188
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7852 5225 7880 5256
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7340 5188 7849 5216
rect 7340 5176 7346 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8104 5219 8162 5225
rect 8104 5185 8116 5219
rect 8150 5216 8162 5219
rect 9122 5216 9128 5228
rect 8150 5188 9128 5216
rect 8150 5185 8162 5188
rect 8104 5179 8162 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9232 5216 9260 5256
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 11146 5284 11152 5296
rect 9355 5256 11152 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 12406 5284 12434 5324
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 22373 5355 22431 5361
rect 22373 5321 22385 5355
rect 22419 5352 22431 5355
rect 22830 5352 22836 5364
rect 22419 5324 22836 5352
rect 22419 5321 22431 5324
rect 22373 5315 22431 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 23290 5312 23296 5364
rect 23348 5312 23354 5364
rect 25590 5312 25596 5364
rect 25648 5312 25654 5364
rect 26602 5312 26608 5364
rect 26660 5312 26666 5364
rect 32490 5312 32496 5364
rect 32548 5312 32554 5364
rect 33134 5312 33140 5364
rect 33192 5352 33198 5364
rect 33229 5355 33287 5361
rect 33229 5352 33241 5355
rect 33192 5324 33241 5352
rect 33192 5312 33198 5324
rect 33229 5321 33241 5324
rect 33275 5321 33287 5355
rect 33229 5315 33287 5321
rect 33778 5312 33784 5364
rect 33836 5352 33842 5364
rect 33965 5355 34023 5361
rect 33965 5352 33977 5355
rect 33836 5324 33977 5352
rect 33836 5312 33842 5324
rect 33965 5321 33977 5324
rect 34011 5321 34023 5355
rect 33965 5315 34023 5321
rect 34698 5312 34704 5364
rect 34756 5352 34762 5364
rect 35161 5355 35219 5361
rect 35161 5352 35173 5355
rect 34756 5324 35173 5352
rect 34756 5312 34762 5324
rect 35161 5321 35173 5324
rect 35207 5321 35219 5355
rect 35161 5315 35219 5321
rect 36173 5355 36231 5361
rect 36173 5321 36185 5355
rect 36219 5352 36231 5355
rect 36814 5352 36820 5364
rect 36219 5324 36820 5352
rect 36219 5321 36231 5324
rect 36173 5315 36231 5321
rect 36814 5312 36820 5324
rect 36872 5312 36878 5364
rect 37550 5312 37556 5364
rect 37608 5352 37614 5364
rect 42797 5355 42855 5361
rect 37608 5324 42748 5352
rect 37608 5312 37614 5324
rect 11624 5256 12434 5284
rect 14001 5287 14059 5293
rect 9858 5216 9864 5228
rect 9232 5188 9864 5216
rect 9858 5176 9864 5188
rect 9916 5216 9922 5228
rect 10042 5216 10048 5228
rect 9916 5188 10048 5216
rect 9916 5176 9922 5188
rect 10042 5176 10048 5188
rect 10100 5216 10106 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10100 5188 10885 5216
rect 10100 5176 10106 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11296 5188 11529 5216
rect 11296 5176 11302 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5031 5120 5304 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5276 5092 5304 5120
rect 1854 5040 1860 5092
rect 1912 5080 1918 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 1912 5052 3341 5080
rect 1912 5040 1918 5052
rect 3329 5049 3341 5052
rect 3375 5080 3387 5083
rect 3418 5080 3424 5092
rect 3375 5052 3424 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3418 5040 3424 5052
rect 3476 5040 3482 5092
rect 3970 5080 3976 5092
rect 3620 5052 3976 5080
rect 2774 4972 2780 5024
rect 2832 4972 2838 5024
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 3234 5012 3240 5024
rect 3007 4984 3240 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3620 5021 3648 5052
rect 3970 5040 3976 5052
rect 4028 5080 4034 5092
rect 4028 5052 5028 5080
rect 4028 5040 4034 5052
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 4981 3663 5015
rect 5000 5012 5028 5052
rect 5258 5040 5264 5092
rect 5316 5040 5322 5092
rect 5350 5040 5356 5092
rect 5408 5080 5414 5092
rect 5408 5052 7788 5080
rect 5408 5040 5414 5052
rect 5810 5012 5816 5024
rect 5000 4984 5816 5012
rect 3605 4975 3663 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 7006 4972 7012 5024
rect 7064 4972 7070 5024
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 7760 5012 7788 5052
rect 9214 5040 9220 5092
rect 9272 5040 9278 5092
rect 11624 5012 11652 5256
rect 14001 5253 14013 5287
rect 14047 5284 14059 5287
rect 14734 5284 14740 5296
rect 14047 5256 14740 5284
rect 14047 5253 14059 5256
rect 14001 5247 14059 5253
rect 14734 5244 14740 5256
rect 14792 5244 14798 5296
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 15473 5287 15531 5293
rect 15473 5284 15485 5287
rect 15252 5256 15485 5284
rect 15252 5244 15258 5256
rect 15473 5253 15485 5256
rect 15519 5253 15531 5287
rect 15930 5284 15936 5296
rect 15473 5247 15531 5253
rect 15764 5256 15936 5284
rect 12434 5176 12440 5228
rect 12492 5176 12498 5228
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15764 5216 15792 5256
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 17678 5293 17684 5296
rect 17672 5284 17684 5293
rect 17639 5256 17684 5284
rect 17672 5247 17684 5256
rect 17678 5244 17684 5247
rect 17736 5244 17742 5296
rect 18414 5244 18420 5296
rect 18472 5284 18478 5296
rect 18966 5284 18972 5296
rect 18472 5256 18972 5284
rect 18472 5244 18478 5256
rect 18966 5244 18972 5256
rect 19024 5284 19030 5296
rect 22189 5287 22247 5293
rect 22189 5284 22201 5287
rect 19024 5256 22201 5284
rect 19024 5244 19030 5256
rect 22189 5253 22201 5256
rect 22235 5253 22247 5287
rect 22189 5247 22247 5253
rect 22741 5287 22799 5293
rect 22741 5253 22753 5287
rect 22787 5284 22799 5287
rect 23308 5284 23336 5312
rect 22787 5256 23336 5284
rect 28160 5287 28218 5293
rect 22787 5253 22799 5256
rect 22741 5247 22799 5253
rect 28160 5253 28172 5287
rect 28206 5284 28218 5287
rect 28258 5284 28264 5296
rect 28206 5256 28264 5284
rect 28206 5253 28218 5256
rect 28160 5247 28218 5253
rect 15427 5188 15792 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15896 5188 16037 5216
rect 15896 5176 15902 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 19334 5216 19340 5228
rect 16540 5188 19340 5216
rect 16540 5176 16546 5188
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 21174 5216 21180 5228
rect 20487 5188 21180 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 17402 5108 17408 5160
rect 17460 5108 17466 5160
rect 19429 5151 19487 5157
rect 19429 5148 19441 5151
rect 18800 5120 19441 5148
rect 16114 5040 16120 5092
rect 16172 5080 16178 5092
rect 18800 5089 18828 5120
rect 19429 5117 19441 5120
rect 19475 5117 19487 5151
rect 22204 5148 22232 5247
rect 28258 5244 28264 5256
rect 28316 5244 28322 5296
rect 31941 5287 31999 5293
rect 31941 5253 31953 5287
rect 31987 5284 31999 5287
rect 35894 5284 35900 5296
rect 31987 5256 35900 5284
rect 31987 5253 31999 5256
rect 31941 5247 31999 5253
rect 35894 5244 35900 5256
rect 35952 5244 35958 5296
rect 36722 5244 36728 5296
rect 36780 5284 36786 5296
rect 39301 5287 39359 5293
rect 39301 5284 39313 5287
rect 36780 5256 39313 5284
rect 36780 5244 36786 5256
rect 39301 5253 39313 5256
rect 39347 5284 39359 5287
rect 41690 5284 41696 5296
rect 39347 5256 41696 5284
rect 39347 5253 39359 5256
rect 39301 5247 39359 5253
rect 41690 5244 41696 5256
rect 41748 5244 41754 5296
rect 42720 5284 42748 5324
rect 42797 5321 42809 5355
rect 42843 5352 42855 5355
rect 43162 5352 43168 5364
rect 42843 5324 43168 5352
rect 42843 5321 42855 5324
rect 42797 5315 42855 5321
rect 43162 5312 43168 5324
rect 43220 5312 43226 5364
rect 45554 5312 45560 5364
rect 45612 5312 45618 5364
rect 45649 5355 45707 5361
rect 45649 5321 45661 5355
rect 45695 5352 45707 5355
rect 46106 5352 46112 5364
rect 45695 5324 46112 5352
rect 45695 5321 45707 5324
rect 45649 5315 45707 5321
rect 46106 5312 46112 5324
rect 46164 5312 46170 5364
rect 47026 5352 47032 5364
rect 46584 5324 47032 5352
rect 43070 5284 43076 5296
rect 42720 5256 43076 5284
rect 43070 5244 43076 5256
rect 43128 5244 43134 5296
rect 44174 5284 44180 5296
rect 43456 5256 44180 5284
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23382 5216 23388 5228
rect 22879 5188 23388 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 25866 5176 25872 5228
rect 25924 5176 25930 5228
rect 26234 5176 26240 5228
rect 26292 5176 26298 5228
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5216 33195 5219
rect 33318 5216 33324 5228
rect 33183 5188 33324 5216
rect 33183 5185 33195 5188
rect 33137 5179 33195 5185
rect 33318 5176 33324 5188
rect 33376 5176 33382 5228
rect 33502 5176 33508 5228
rect 33560 5216 33566 5228
rect 33781 5219 33839 5225
rect 33781 5216 33793 5219
rect 33560 5188 33793 5216
rect 33560 5176 33566 5188
rect 33781 5185 33793 5188
rect 33827 5185 33839 5219
rect 33781 5179 33839 5185
rect 34514 5176 34520 5228
rect 34572 5176 34578 5228
rect 34698 5176 34704 5228
rect 34756 5176 34762 5228
rect 34882 5176 34888 5228
rect 34940 5176 34946 5228
rect 35912 5216 35940 5244
rect 37001 5219 37059 5225
rect 37001 5216 37013 5219
rect 35912 5188 37013 5216
rect 37001 5185 37013 5188
rect 37047 5185 37059 5219
rect 37001 5179 37059 5185
rect 37369 5219 37427 5225
rect 37369 5185 37381 5219
rect 37415 5216 37427 5219
rect 37458 5216 37464 5228
rect 37415 5188 37464 5216
rect 37415 5185 37427 5188
rect 37369 5179 37427 5185
rect 37458 5176 37464 5188
rect 37516 5176 37522 5228
rect 37636 5219 37694 5225
rect 37636 5185 37648 5219
rect 37682 5216 37694 5219
rect 38194 5216 38200 5228
rect 37682 5188 38200 5216
rect 37682 5185 37694 5188
rect 37636 5179 37694 5185
rect 38194 5176 38200 5188
rect 38252 5176 38258 5228
rect 39114 5176 39120 5228
rect 39172 5216 39178 5228
rect 39172 5188 43024 5216
rect 39172 5176 39178 5188
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 22204 5120 22937 5148
rect 19429 5111 19487 5117
rect 22925 5117 22937 5120
rect 22971 5148 22983 5151
rect 25314 5148 25320 5160
rect 22971 5120 25320 5148
rect 22971 5117 22983 5120
rect 22925 5111 22983 5117
rect 25314 5108 25320 5120
rect 25372 5108 25378 5160
rect 25884 5148 25912 5176
rect 27893 5151 27951 5157
rect 27893 5148 27905 5151
rect 25884 5120 27905 5148
rect 27893 5117 27905 5120
rect 27939 5117 27951 5151
rect 27893 5111 27951 5117
rect 29549 5151 29607 5157
rect 29549 5117 29561 5151
rect 29595 5117 29607 5151
rect 34716 5148 34744 5176
rect 35529 5151 35587 5157
rect 35529 5148 35541 5151
rect 34716 5120 35541 5148
rect 29549 5111 29607 5117
rect 35529 5117 35541 5120
rect 35575 5117 35587 5151
rect 35529 5111 35587 5117
rect 17221 5083 17279 5089
rect 17221 5080 17233 5083
rect 16172 5052 17233 5080
rect 16172 5040 16178 5052
rect 17221 5049 17233 5052
rect 17267 5049 17279 5083
rect 17221 5043 17279 5049
rect 18785 5083 18843 5089
rect 18785 5049 18797 5083
rect 18831 5049 18843 5083
rect 18785 5043 18843 5049
rect 29273 5083 29331 5089
rect 29273 5049 29285 5083
rect 29319 5080 29331 5083
rect 29564 5080 29592 5111
rect 39942 5108 39948 5160
rect 40000 5148 40006 5160
rect 40862 5148 40868 5160
rect 40000 5120 40868 5148
rect 40000 5108 40006 5120
rect 40862 5108 40868 5120
rect 40920 5148 40926 5160
rect 41049 5151 41107 5157
rect 41049 5148 41061 5151
rect 40920 5120 41061 5148
rect 40920 5108 40926 5120
rect 41049 5117 41061 5120
rect 41095 5148 41107 5151
rect 41506 5148 41512 5160
rect 41095 5120 41512 5148
rect 41095 5117 41107 5120
rect 41049 5111 41107 5117
rect 41506 5108 41512 5120
rect 41564 5108 41570 5160
rect 42245 5151 42303 5157
rect 42245 5117 42257 5151
rect 42291 5148 42303 5151
rect 42889 5151 42947 5157
rect 42291 5120 42472 5148
rect 42291 5117 42303 5120
rect 42245 5111 42303 5117
rect 36170 5080 36176 5092
rect 29319 5052 29592 5080
rect 31726 5052 36176 5080
rect 29319 5049 29331 5052
rect 29273 5043 29331 5049
rect 7760 4984 11652 5012
rect 14829 5015 14887 5021
rect 14829 4981 14841 5015
rect 14875 5012 14887 5015
rect 14918 5012 14924 5024
rect 14875 4984 14924 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 14918 4972 14924 4984
rect 14976 5012 14982 5024
rect 17586 5012 17592 5024
rect 14976 4984 17592 5012
rect 14976 4972 14982 4984
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18196 4984 18889 5012
rect 18196 4972 18202 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18877 4975 18935 4981
rect 19886 4972 19892 5024
rect 19944 5012 19950 5024
rect 20990 5012 20996 5024
rect 19944 4984 20996 5012
rect 19944 4972 19950 4984
rect 20990 4972 20996 4984
rect 21048 4972 21054 5024
rect 21361 5015 21419 5021
rect 21361 4981 21373 5015
rect 21407 5012 21419 5015
rect 21726 5012 21732 5024
rect 21407 4984 21732 5012
rect 21407 4981 21419 4984
rect 21361 4975 21419 4981
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 23290 4972 23296 5024
rect 23348 5012 23354 5024
rect 23385 5015 23443 5021
rect 23385 5012 23397 5015
rect 23348 4984 23397 5012
rect 23348 4972 23354 4984
rect 23385 4981 23397 4984
rect 23431 4981 23443 5015
rect 23385 4975 23443 4981
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 24026 5012 24032 5024
rect 23891 4984 24032 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 30193 5015 30251 5021
rect 30193 4981 30205 5015
rect 30239 5012 30251 5015
rect 30282 5012 30288 5024
rect 30239 4984 30288 5012
rect 30239 4981 30251 4984
rect 30193 4975 30251 4981
rect 30282 4972 30288 4984
rect 30340 4972 30346 5024
rect 30650 4972 30656 5024
rect 30708 5012 30714 5024
rect 31726 5012 31754 5052
rect 36170 5040 36176 5052
rect 36228 5040 36234 5092
rect 42444 5089 42472 5120
rect 42889 5117 42901 5151
rect 42935 5117 42947 5151
rect 42996 5148 43024 5188
rect 43073 5151 43131 5157
rect 43073 5148 43085 5151
rect 42996 5120 43085 5148
rect 42889 5111 42947 5117
rect 43073 5117 43085 5120
rect 43119 5148 43131 5151
rect 43456 5148 43484 5256
rect 44174 5244 44180 5256
rect 44232 5244 44238 5296
rect 45312 5287 45370 5293
rect 45312 5253 45324 5287
rect 45358 5284 45370 5287
rect 45572 5284 45600 5312
rect 45358 5256 45600 5284
rect 46017 5287 46075 5293
rect 45358 5253 45370 5256
rect 45312 5247 45370 5253
rect 46017 5253 46029 5287
rect 46063 5284 46075 5287
rect 46584 5284 46612 5324
rect 47026 5312 47032 5324
rect 47084 5312 47090 5364
rect 49694 5312 49700 5364
rect 49752 5352 49758 5364
rect 49973 5355 50031 5361
rect 49973 5352 49985 5355
rect 49752 5324 49985 5352
rect 49752 5312 49758 5324
rect 49973 5321 49985 5324
rect 50019 5321 50031 5355
rect 49973 5315 50031 5321
rect 51169 5355 51227 5361
rect 51169 5321 51181 5355
rect 51215 5352 51227 5355
rect 51350 5352 51356 5364
rect 51215 5324 51356 5352
rect 51215 5321 51227 5324
rect 51169 5315 51227 5321
rect 51350 5312 51356 5324
rect 51408 5312 51414 5364
rect 51537 5355 51595 5361
rect 51537 5321 51549 5355
rect 51583 5352 51595 5355
rect 51626 5352 51632 5364
rect 51583 5324 51632 5352
rect 51583 5321 51595 5324
rect 51537 5315 51595 5321
rect 51626 5312 51632 5324
rect 51684 5312 51690 5364
rect 51905 5355 51963 5361
rect 51905 5321 51917 5355
rect 51951 5352 51963 5355
rect 51951 5324 52684 5352
rect 51951 5321 51963 5324
rect 51905 5315 51963 5321
rect 47305 5287 47363 5293
rect 47305 5284 47317 5287
rect 46063 5256 46612 5284
rect 46860 5256 47317 5284
rect 46063 5253 46075 5256
rect 46017 5247 46075 5253
rect 44085 5219 44143 5225
rect 44085 5185 44097 5219
rect 44131 5216 44143 5219
rect 45557 5219 45615 5225
rect 44131 5188 45508 5216
rect 44131 5185 44143 5188
rect 44085 5179 44143 5185
rect 43119 5120 43484 5148
rect 43533 5151 43591 5157
rect 43119 5117 43131 5120
rect 43073 5111 43131 5117
rect 43533 5117 43545 5151
rect 43579 5117 43591 5151
rect 45480 5148 45508 5188
rect 45557 5185 45569 5219
rect 45603 5216 45615 5219
rect 45922 5216 45928 5228
rect 45603 5188 45928 5216
rect 45603 5185 45615 5188
rect 45557 5179 45615 5185
rect 45922 5176 45928 5188
rect 45980 5176 45986 5228
rect 46474 5176 46480 5228
rect 46532 5216 46538 5228
rect 46860 5225 46888 5256
rect 47305 5253 47317 5256
rect 47351 5284 47363 5287
rect 51994 5284 52000 5296
rect 47351 5256 52000 5284
rect 47351 5253 47363 5256
rect 47305 5247 47363 5253
rect 51994 5244 52000 5256
rect 52052 5284 52058 5296
rect 52362 5284 52368 5296
rect 52052 5256 52368 5284
rect 52052 5244 52058 5256
rect 52362 5244 52368 5256
rect 52420 5244 52426 5296
rect 52656 5284 52684 5324
rect 52730 5312 52736 5364
rect 52788 5312 52794 5364
rect 53101 5355 53159 5361
rect 53101 5321 53113 5355
rect 53147 5352 53159 5355
rect 53374 5352 53380 5364
rect 53147 5324 53380 5352
rect 53147 5321 53159 5324
rect 53101 5315 53159 5321
rect 53374 5312 53380 5324
rect 53432 5312 53438 5364
rect 55401 5355 55459 5361
rect 55401 5321 55413 5355
rect 55447 5352 55459 5355
rect 55490 5352 55496 5364
rect 55447 5324 55496 5352
rect 55447 5321 55459 5324
rect 55401 5315 55459 5321
rect 55490 5312 55496 5324
rect 55548 5312 55554 5364
rect 55582 5312 55588 5364
rect 55640 5352 55646 5364
rect 55769 5355 55827 5361
rect 55769 5352 55781 5355
rect 55640 5324 55781 5352
rect 55640 5312 55646 5324
rect 55769 5321 55781 5324
rect 55815 5321 55827 5355
rect 55769 5315 55827 5321
rect 57698 5312 57704 5364
rect 57756 5312 57762 5364
rect 52656 5256 53880 5284
rect 46845 5219 46903 5225
rect 46845 5216 46857 5219
rect 46532 5188 46857 5216
rect 46532 5176 46538 5188
rect 46845 5185 46857 5188
rect 46891 5185 46903 5219
rect 46845 5179 46903 5185
rect 47029 5219 47087 5225
rect 47029 5185 47041 5219
rect 47075 5216 47087 5219
rect 47581 5219 47639 5225
rect 47581 5216 47593 5219
rect 47075 5188 47593 5216
rect 47075 5185 47087 5188
rect 47029 5179 47087 5185
rect 47581 5185 47593 5188
rect 47627 5185 47639 5219
rect 47581 5179 47639 5185
rect 47688 5188 48268 5216
rect 45646 5148 45652 5160
rect 45480 5120 45652 5148
rect 43533 5111 43591 5117
rect 42429 5083 42487 5089
rect 42429 5049 42441 5083
rect 42475 5049 42487 5083
rect 42429 5043 42487 5049
rect 30708 4984 31754 5012
rect 30708 4972 30714 4984
rect 32398 4972 32404 5024
rect 32456 5012 32462 5024
rect 34054 5012 34060 5024
rect 32456 4984 34060 5012
rect 32456 4972 32462 4984
rect 34054 4972 34060 4984
rect 34112 4972 34118 5024
rect 34790 4972 34796 5024
rect 34848 5012 34854 5024
rect 34885 5015 34943 5021
rect 34885 5012 34897 5015
rect 34848 4984 34897 5012
rect 34848 4972 34854 4984
rect 34885 4981 34897 4984
rect 34931 4981 34943 5015
rect 34885 4975 34943 4981
rect 38746 4972 38752 5024
rect 38804 4972 38810 5024
rect 38838 4972 38844 5024
rect 38896 5012 38902 5024
rect 39025 5015 39083 5021
rect 39025 5012 39037 5015
rect 38896 4984 39037 5012
rect 38896 4972 38902 4984
rect 39025 4981 39037 4984
rect 39071 4981 39083 5015
rect 39025 4975 39083 4981
rect 40678 4972 40684 5024
rect 40736 5012 40742 5024
rect 41417 5015 41475 5021
rect 41417 5012 41429 5015
rect 40736 4984 41429 5012
rect 40736 4972 40742 4984
rect 41417 4981 41429 4984
rect 41463 5012 41475 5015
rect 41506 5012 41512 5024
rect 41463 4984 41512 5012
rect 41463 4981 41475 4984
rect 41417 4975 41475 4981
rect 41506 4972 41512 4984
rect 41564 4972 41570 5024
rect 41598 4972 41604 5024
rect 41656 4972 41662 5024
rect 42242 4972 42248 5024
rect 42300 5012 42306 5024
rect 42904 5012 42932 5111
rect 43548 5080 43576 5111
rect 45646 5108 45652 5120
rect 45704 5148 45710 5160
rect 46109 5151 46167 5157
rect 46109 5148 46121 5151
rect 45704 5120 46121 5148
rect 45704 5108 45710 5120
rect 46109 5117 46121 5120
rect 46155 5117 46167 5151
rect 46109 5111 46167 5117
rect 46290 5108 46296 5160
rect 46348 5148 46354 5160
rect 46753 5151 46811 5157
rect 46753 5148 46765 5151
rect 46348 5120 46765 5148
rect 46348 5108 46354 5120
rect 46753 5117 46765 5120
rect 46799 5148 46811 5151
rect 47688 5148 47716 5188
rect 46799 5120 47716 5148
rect 46799 5117 46811 5120
rect 46753 5111 46811 5117
rect 47854 5108 47860 5160
rect 47912 5148 47918 5160
rect 48133 5151 48191 5157
rect 48133 5148 48145 5151
rect 47912 5120 48145 5148
rect 47912 5108 47918 5120
rect 48133 5117 48145 5120
rect 48179 5117 48191 5151
rect 48240 5148 48268 5188
rect 50430 5176 50436 5228
rect 50488 5216 50494 5228
rect 50525 5219 50583 5225
rect 50525 5216 50537 5219
rect 50488 5188 50537 5216
rect 50488 5176 50494 5188
rect 50525 5185 50537 5188
rect 50571 5185 50583 5219
rect 50525 5179 50583 5185
rect 51258 5176 51264 5228
rect 51316 5216 51322 5228
rect 52181 5219 52239 5225
rect 52181 5216 52193 5219
rect 51316 5188 52193 5216
rect 51316 5176 51322 5188
rect 52181 5185 52193 5188
rect 52227 5185 52239 5219
rect 52181 5179 52239 5185
rect 53193 5219 53251 5225
rect 53193 5185 53205 5219
rect 53239 5216 53251 5219
rect 53558 5216 53564 5228
rect 53239 5188 53564 5216
rect 53239 5185 53251 5188
rect 53193 5179 53251 5185
rect 53558 5176 53564 5188
rect 53616 5176 53622 5228
rect 53852 5225 53880 5256
rect 53837 5219 53895 5225
rect 53837 5185 53849 5219
rect 53883 5216 53895 5219
rect 53926 5216 53932 5228
rect 53883 5188 53932 5216
rect 53883 5185 53895 5188
rect 53837 5179 53895 5185
rect 53926 5176 53932 5188
rect 53984 5216 53990 5228
rect 55122 5216 55128 5228
rect 53984 5188 55128 5216
rect 53984 5176 53990 5188
rect 55122 5176 55128 5188
rect 55180 5176 55186 5228
rect 55398 5216 55404 5228
rect 55232 5188 55404 5216
rect 55232 5157 55260 5188
rect 55398 5176 55404 5188
rect 55456 5216 55462 5228
rect 55456 5188 55996 5216
rect 55456 5176 55462 5188
rect 55968 5157 55996 5188
rect 56318 5176 56324 5228
rect 56376 5176 56382 5228
rect 56410 5176 56416 5228
rect 56468 5216 56474 5228
rect 56577 5219 56635 5225
rect 56577 5216 56589 5219
rect 56468 5188 56589 5216
rect 56468 5176 56474 5188
rect 56577 5185 56589 5188
rect 56623 5185 56635 5219
rect 56577 5179 56635 5185
rect 58434 5176 58440 5228
rect 58492 5176 58498 5228
rect 52457 5151 52515 5157
rect 52457 5148 52469 5151
rect 48240 5120 52469 5148
rect 48133 5111 48191 5117
rect 52457 5117 52469 5120
rect 52503 5148 52515 5151
rect 53285 5151 53343 5157
rect 53285 5148 53297 5151
rect 52503 5120 53297 5148
rect 52503 5117 52515 5120
rect 52457 5111 52515 5117
rect 53285 5117 53297 5120
rect 53331 5148 53343 5151
rect 55217 5151 55275 5157
rect 55217 5148 55229 5151
rect 53331 5120 55229 5148
rect 53331 5117 53343 5120
rect 53285 5111 53343 5117
rect 55217 5117 55229 5120
rect 55263 5117 55275 5151
rect 55217 5111 55275 5117
rect 55861 5151 55919 5157
rect 55861 5117 55873 5151
rect 55907 5117 55919 5151
rect 55861 5111 55919 5117
rect 55953 5151 56011 5157
rect 55953 5117 55965 5151
rect 55999 5117 56011 5151
rect 55953 5111 56011 5117
rect 44177 5083 44235 5089
rect 44177 5080 44189 5083
rect 43548 5052 44189 5080
rect 44177 5049 44189 5052
rect 44223 5049 44235 5083
rect 44177 5043 44235 5049
rect 45572 5052 49372 5080
rect 42300 4984 42932 5012
rect 42300 4972 42306 4984
rect 43070 4972 43076 5024
rect 43128 5012 43134 5024
rect 45572 5012 45600 5052
rect 49344 5024 49372 5052
rect 50246 5040 50252 5092
rect 50304 5080 50310 5092
rect 51997 5083 52055 5089
rect 51997 5080 52009 5083
rect 50304 5052 52009 5080
rect 50304 5040 50310 5052
rect 51997 5049 52009 5052
rect 52043 5049 52055 5083
rect 51997 5043 52055 5049
rect 54205 5083 54263 5089
rect 54205 5049 54217 5083
rect 54251 5080 54263 5083
rect 55876 5080 55904 5111
rect 56318 5080 56324 5092
rect 54251 5052 54984 5080
rect 55876 5052 56324 5080
rect 54251 5049 54263 5052
rect 54205 5043 54263 5049
rect 43128 4984 45600 5012
rect 43128 4972 43134 4984
rect 46842 4972 46848 5024
rect 46900 5012 46906 5024
rect 47029 5015 47087 5021
rect 47029 5012 47041 5015
rect 46900 4984 47041 5012
rect 46900 4972 46906 4984
rect 47029 4981 47041 4984
rect 47075 4981 47087 5015
rect 47029 4975 47087 4981
rect 49326 4972 49332 5024
rect 49384 4972 49390 5024
rect 49694 4972 49700 5024
rect 49752 5012 49758 5024
rect 50433 5015 50491 5021
rect 50433 5012 50445 5015
rect 49752 4984 50445 5012
rect 49752 4972 49758 4984
rect 50433 4981 50445 4984
rect 50479 5012 50491 5015
rect 50982 5012 50988 5024
rect 50479 4984 50988 5012
rect 50479 4981 50491 4984
rect 50433 4975 50491 4981
rect 50982 4972 50988 4984
rect 51040 4972 51046 5024
rect 51350 4972 51356 5024
rect 51408 5012 51414 5024
rect 54220 5012 54248 5043
rect 51408 4984 54248 5012
rect 54573 5015 54631 5021
rect 51408 4972 51414 4984
rect 54573 4981 54585 5015
rect 54619 5012 54631 5015
rect 54662 5012 54668 5024
rect 54619 4984 54668 5012
rect 54619 4981 54631 4984
rect 54573 4975 54631 4981
rect 54662 4972 54668 4984
rect 54720 4972 54726 5024
rect 54846 4972 54852 5024
rect 54904 4972 54910 5024
rect 54956 5012 54984 5052
rect 56318 5040 56324 5052
rect 56376 5040 56382 5092
rect 56962 5012 56968 5024
rect 54956 4984 56968 5012
rect 56962 4972 56968 4984
rect 57020 4972 57026 5024
rect 57882 4972 57888 5024
rect 57940 4972 57946 5024
rect 1104 4922 58880 4944
rect 1104 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 22616 4922
rect 22668 4870 22680 4922
rect 22732 4870 22744 4922
rect 22796 4870 22808 4922
rect 22860 4870 22872 4922
rect 22924 4870 37060 4922
rect 37112 4870 37124 4922
rect 37176 4870 37188 4922
rect 37240 4870 37252 4922
rect 37304 4870 37316 4922
rect 37368 4870 51504 4922
rect 51556 4870 51568 4922
rect 51620 4870 51632 4922
rect 51684 4870 51696 4922
rect 51748 4870 51760 4922
rect 51812 4870 58880 4922
rect 1104 4848 58880 4870
rect 2774 4768 2780 4820
rect 2832 4768 2838 4820
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3292 4780 3801 4808
rect 3292 4768 3298 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 7742 4808 7748 4820
rect 5123 4780 7748 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 9122 4768 9128 4820
rect 9180 4768 9186 4820
rect 9232 4780 11100 4808
rect 2792 4672 2820 4768
rect 4525 4743 4583 4749
rect 4525 4709 4537 4743
rect 4571 4740 4583 4743
rect 4571 4712 5856 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 2792 4644 3341 4672
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 4430 4632 4436 4684
rect 4488 4632 4494 4684
rect 4724 4644 5304 4672
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 3476 4576 4537 4604
rect 3476 4564 3482 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4724 4604 4752 4644
rect 5276 4616 5304 4644
rect 4797 4607 4855 4613
rect 4797 4604 4809 4607
rect 4724 4576 4809 4604
rect 4525 4567 4583 4573
rect 4797 4573 4809 4576
rect 4843 4573 4855 4607
rect 4797 4567 4855 4573
rect 4890 4564 4896 4616
rect 4948 4613 4954 4616
rect 4948 4567 4959 4613
rect 4948 4564 4954 4567
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 5828 4613 5856 4712
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 9232 4740 9260 4780
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 7064 4712 9260 4740
rect 9784 4712 10057 4740
rect 7064 4700 7070 4712
rect 9784 4681 9812 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10962 4740 10968 4752
rect 10045 4703 10103 4709
rect 10704 4712 10968 4740
rect 10704 4681 10732 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11072 4740 11100 4780
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 11609 4811 11667 4817
rect 11609 4777 11621 4811
rect 11655 4808 11667 4811
rect 11698 4808 11704 4820
rect 11655 4780 11704 4808
rect 11655 4777 11667 4780
rect 11609 4771 11667 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 13081 4811 13139 4817
rect 13081 4777 13093 4811
rect 13127 4808 13139 4811
rect 13446 4808 13452 4820
rect 13127 4780 13452 4808
rect 13127 4777 13139 4780
rect 13081 4771 13139 4777
rect 13446 4768 13452 4780
rect 13504 4808 13510 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 13504 4780 15117 4808
rect 13504 4768 13510 4780
rect 15105 4777 15117 4780
rect 15151 4808 15163 4811
rect 15194 4808 15200 4820
rect 15151 4780 15200 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15194 4768 15200 4780
rect 15252 4808 15258 4820
rect 16482 4808 16488 4820
rect 15252 4780 16488 4808
rect 15252 4768 15258 4780
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 17681 4811 17739 4817
rect 16632 4780 16896 4808
rect 16632 4768 16638 4780
rect 16758 4740 16764 4752
rect 11072 4712 16764 4740
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 16868 4740 16896 4780
rect 17681 4777 17693 4811
rect 17727 4808 17739 4811
rect 17954 4808 17960 4820
rect 17727 4780 17960 4808
rect 17727 4777 17739 4780
rect 17681 4771 17739 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 18380 4780 19349 4808
rect 18380 4768 18386 4780
rect 19337 4777 19349 4780
rect 19383 4777 19395 4811
rect 19337 4771 19395 4777
rect 20990 4768 20996 4820
rect 21048 4808 21054 4820
rect 21450 4808 21456 4820
rect 21048 4780 21456 4808
rect 21048 4768 21054 4780
rect 21450 4768 21456 4780
rect 21508 4808 21514 4820
rect 21545 4811 21603 4817
rect 21545 4808 21557 4811
rect 21508 4780 21557 4808
rect 21508 4768 21514 4780
rect 21545 4777 21557 4780
rect 21591 4808 21603 4811
rect 24762 4808 24768 4820
rect 21591 4780 24768 4808
rect 21591 4777 21603 4780
rect 21545 4771 21603 4777
rect 24762 4768 24768 4780
rect 24820 4808 24826 4820
rect 24857 4811 24915 4817
rect 24857 4808 24869 4811
rect 24820 4780 24869 4808
rect 24820 4768 24826 4780
rect 24857 4777 24869 4780
rect 24903 4777 24915 4811
rect 24857 4771 24915 4777
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 25133 4811 25191 4817
rect 25133 4808 25145 4811
rect 25096 4780 25145 4808
rect 25096 4768 25102 4780
rect 25133 4777 25145 4780
rect 25179 4777 25191 4811
rect 25133 4771 25191 4777
rect 25314 4768 25320 4820
rect 25372 4808 25378 4820
rect 28077 4811 28135 4817
rect 28077 4808 28089 4811
rect 25372 4780 28089 4808
rect 25372 4768 25378 4780
rect 28077 4777 28089 4780
rect 28123 4777 28135 4811
rect 28077 4771 28135 4777
rect 28261 4811 28319 4817
rect 28261 4777 28273 4811
rect 28307 4808 28319 4811
rect 28810 4808 28816 4820
rect 28307 4780 28816 4808
rect 28307 4777 28319 4780
rect 28261 4771 28319 4777
rect 16868 4712 27844 4740
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 9769 4675 9827 4681
rect 7331 4644 9168 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6135 4576 6561 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6549 4573 6561 4576
rect 6595 4604 6607 4607
rect 6917 4607 6975 4613
rect 6917 4604 6929 4607
rect 6595 4576 6929 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 6917 4573 6929 4576
rect 6963 4604 6975 4607
rect 7374 4604 7380 4616
rect 6963 4576 7380 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 4709 4539 4767 4545
rect 2148 4508 4660 4536
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2148 4477 2176 4508
rect 2133 4471 2191 4477
rect 2133 4468 2145 4471
rect 2004 4440 2145 4468
rect 2004 4428 2010 4440
rect 2133 4437 2145 4440
rect 2179 4437 2191 4471
rect 2133 4431 2191 4437
rect 2774 4428 2780 4480
rect 2832 4428 2838 4480
rect 4632 4468 4660 4508
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 5718 4536 5724 4548
rect 4755 4508 5724 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 4982 4468 4988 4480
rect 4632 4440 4988 4468
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5537 4471 5595 4477
rect 5537 4468 5549 4471
rect 5316 4440 5549 4468
rect 5316 4428 5322 4440
rect 5537 4437 5549 4440
rect 5583 4468 5595 4471
rect 6104 4468 6132 4567
rect 7374 4564 7380 4576
rect 7432 4604 7438 4616
rect 8110 4604 8116 4616
rect 7432 4576 8116 4604
rect 7432 4564 7438 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 8444 4576 8677 4604
rect 8444 4564 8450 4576
rect 8665 4573 8677 4576
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 9140 4548 9168 4644
rect 9769 4641 9781 4675
rect 9815 4641 9827 4675
rect 9769 4635 9827 4641
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 16574 4672 16580 4684
rect 10689 4635 10747 4641
rect 10796 4644 16580 4672
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10502 4604 10508 4616
rect 10459 4576 10508 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10796 4604 10824 4644
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 18138 4632 18144 4684
rect 18196 4632 18202 4684
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 18414 4672 18420 4684
rect 18371 4644 18420 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 18414 4632 18420 4644
rect 18472 4632 18478 4684
rect 24946 4672 24952 4684
rect 18524 4644 20300 4672
rect 10612 4576 10824 4604
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8021 4539 8079 4545
rect 8021 4536 8033 4539
rect 7699 4508 8033 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8021 4505 8033 4508
rect 8067 4536 8079 4539
rect 8067 4508 8340 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8312 4480 8340 4508
rect 9122 4496 9128 4548
rect 9180 4536 9186 4548
rect 10612 4536 10640 4576
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 13780 4576 14657 4604
rect 13780 4564 13786 4576
rect 14645 4573 14657 4576
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 16022 4564 16028 4616
rect 16080 4564 16086 4616
rect 17586 4564 17592 4616
rect 17644 4604 17650 4616
rect 18524 4613 18552 4644
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 17644 4576 18521 4604
rect 17644 4564 17650 4576
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 18690 4564 18696 4616
rect 18748 4564 18754 4616
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 9180 4508 10640 4536
rect 9180 4496 9186 4508
rect 10962 4496 10968 4548
rect 11020 4536 11026 4548
rect 13998 4536 14004 4548
rect 11020 4508 14004 4536
rect 11020 4496 11026 4508
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 14090 4496 14096 4548
rect 14148 4496 14154 4548
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 17129 4539 17187 4545
rect 17129 4536 17141 4539
rect 14240 4508 17141 4536
rect 14240 4496 14246 4508
rect 17129 4505 17141 4508
rect 17175 4505 17187 4539
rect 17129 4499 17187 4505
rect 18049 4539 18107 4545
rect 18049 4505 18061 4539
rect 18095 4536 18107 4539
rect 18230 4536 18236 4548
rect 18095 4508 18236 4536
rect 18095 4505 18107 4508
rect 18049 4499 18107 4505
rect 18230 4496 18236 4508
rect 18288 4496 18294 4548
rect 18322 4496 18328 4548
rect 18380 4536 18386 4548
rect 18984 4536 19012 4567
rect 19334 4564 19340 4616
rect 19392 4564 19398 4616
rect 19518 4564 19524 4616
rect 19576 4564 19582 4616
rect 20272 4613 20300 4644
rect 20732 4644 21772 4672
rect 20732 4613 20760 4644
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4604 20315 4607
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20303 4576 20637 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 20625 4573 20637 4576
rect 20671 4604 20683 4607
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20671 4576 20729 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20717 4567 20775 4573
rect 20898 4564 20904 4616
rect 20956 4564 20962 4616
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 18380 4508 19012 4536
rect 19352 4536 19380 4564
rect 21744 4548 21772 4644
rect 23860 4644 24952 4672
rect 23860 4613 23888 4644
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 25038 4632 25044 4684
rect 25096 4672 25102 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 25096 4644 26801 4672
rect 25096 4632 25102 4644
rect 26789 4641 26801 4644
rect 26835 4672 26847 4675
rect 27522 4672 27528 4684
rect 26835 4644 27528 4672
rect 26835 4641 26847 4644
rect 26789 4635 26847 4641
rect 27522 4632 27528 4644
rect 27580 4672 27586 4684
rect 27709 4675 27767 4681
rect 27709 4672 27721 4675
rect 27580 4644 27721 4672
rect 27580 4632 27586 4644
rect 27709 4641 27721 4644
rect 27755 4641 27767 4675
rect 27709 4635 27767 4641
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 23845 4607 23903 4613
rect 23845 4604 23857 4607
rect 22051 4576 23857 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 23845 4573 23857 4576
rect 23891 4573 23903 4607
rect 23845 4567 23903 4573
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4604 24455 4607
rect 25222 4604 25228 4616
rect 24443 4576 25228 4604
rect 24443 4573 24455 4576
rect 24397 4567 24455 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 25314 4564 25320 4616
rect 25372 4564 25378 4616
rect 26329 4607 26387 4613
rect 26329 4573 26341 4607
rect 26375 4604 26387 4607
rect 26375 4576 26409 4604
rect 26375 4573 26387 4576
rect 26329 4567 26387 4573
rect 19797 4539 19855 4545
rect 19797 4536 19809 4539
rect 19352 4508 19809 4536
rect 18380 4496 18386 4508
rect 19797 4505 19809 4508
rect 19843 4536 19855 4539
rect 20070 4536 20076 4548
rect 19843 4508 20076 4536
rect 19843 4505 19855 4508
rect 19797 4499 19855 4505
rect 20070 4496 20076 4508
rect 20128 4496 20134 4548
rect 20438 4496 20444 4548
rect 20496 4536 20502 4548
rect 20809 4539 20867 4545
rect 20809 4536 20821 4539
rect 20496 4508 20821 4536
rect 20496 4496 20502 4508
rect 20809 4505 20821 4508
rect 20855 4505 20867 4539
rect 20809 4499 20867 4505
rect 21726 4496 21732 4548
rect 21784 4536 21790 4548
rect 24026 4536 24032 4548
rect 21784 4508 24032 4536
rect 21784 4496 21790 4508
rect 24026 4496 24032 4508
rect 24084 4536 24090 4548
rect 26145 4539 26203 4545
rect 26145 4536 26157 4539
rect 24084 4508 26157 4536
rect 24084 4496 24090 4508
rect 26145 4505 26157 4508
rect 26191 4536 26203 4539
rect 26344 4536 26372 4567
rect 26510 4564 26516 4616
rect 26568 4564 26574 4616
rect 26191 4508 27476 4536
rect 26191 4505 26203 4508
rect 26145 4499 26203 4505
rect 5583 4440 6132 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 7892 4440 8125 4468
rect 7892 4428 7898 4440
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 8294 4428 8300 4480
rect 8352 4428 8358 4480
rect 10502 4428 10508 4480
rect 10560 4428 10566 4480
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4468 12219 4471
rect 12434 4468 12440 4480
rect 12207 4440 12440 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 12434 4428 12440 4440
rect 12492 4468 12498 4480
rect 13541 4471 13599 4477
rect 13541 4468 13553 4471
rect 12492 4440 13553 4468
rect 12492 4428 12498 4440
rect 13541 4437 13553 4440
rect 13587 4468 13599 4471
rect 13909 4471 13967 4477
rect 13909 4468 13921 4471
rect 13587 4440 13921 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13909 4437 13921 4440
rect 13955 4468 13967 4471
rect 14274 4468 14280 4480
rect 13955 4440 14280 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14274 4428 14280 4440
rect 14332 4468 14338 4480
rect 14918 4468 14924 4480
rect 14332 4440 14924 4468
rect 14332 4428 14338 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15473 4471 15531 4477
rect 15473 4468 15485 4471
rect 15160 4440 15485 4468
rect 15160 4428 15166 4440
rect 15473 4437 15485 4440
rect 15519 4437 15531 4471
rect 15473 4431 15531 4437
rect 16114 4428 16120 4480
rect 16172 4468 16178 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16172 4440 16405 4468
rect 16172 4428 16178 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16393 4431 16451 4437
rect 18598 4428 18604 4480
rect 18656 4428 18662 4480
rect 18782 4428 18788 4480
rect 18840 4428 18846 4480
rect 20622 4428 20628 4480
rect 20680 4468 20686 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 20680 4440 21097 4468
rect 20680 4428 20686 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 22373 4471 22431 4477
rect 22373 4468 22385 4471
rect 22336 4440 22385 4468
rect 22336 4428 22342 4440
rect 22373 4437 22385 4440
rect 22419 4437 22431 4471
rect 22373 4431 22431 4437
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 24121 4471 24179 4477
rect 24121 4468 24133 4471
rect 23348 4440 24133 4468
rect 23348 4428 23354 4440
rect 24121 4437 24133 4440
rect 24167 4468 24179 4471
rect 24210 4468 24216 4480
rect 24167 4440 24216 4468
rect 24167 4437 24179 4440
rect 24121 4431 24179 4437
rect 24210 4428 24216 4440
rect 24268 4428 24274 4480
rect 24578 4428 24584 4480
rect 24636 4428 24642 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 27448 4477 27476 4508
rect 26421 4471 26479 4477
rect 26421 4468 26433 4471
rect 26292 4440 26433 4468
rect 26292 4428 26298 4440
rect 26421 4437 26433 4440
rect 26467 4437 26479 4471
rect 26421 4431 26479 4437
rect 27433 4471 27491 4477
rect 27433 4437 27445 4471
rect 27479 4468 27491 4471
rect 27614 4468 27620 4480
rect 27479 4440 27620 4468
rect 27479 4437 27491 4440
rect 27433 4431 27491 4437
rect 27614 4428 27620 4440
rect 27672 4428 27678 4480
rect 27724 4468 27752 4635
rect 27816 4604 27844 4712
rect 28092 4672 28120 4771
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 28902 4768 28908 4820
rect 28960 4808 28966 4820
rect 31386 4808 31392 4820
rect 28960 4780 31392 4808
rect 28960 4768 28966 4780
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 34146 4808 34152 4820
rect 32600 4780 34152 4808
rect 28166 4700 28172 4752
rect 28224 4740 28230 4752
rect 32600 4740 32628 4780
rect 34146 4768 34152 4780
rect 34204 4768 34210 4820
rect 34793 4811 34851 4817
rect 34793 4777 34805 4811
rect 34839 4808 34851 4811
rect 34882 4808 34888 4820
rect 34839 4780 34888 4808
rect 34839 4777 34851 4780
rect 34793 4771 34851 4777
rect 34882 4768 34888 4780
rect 34940 4768 34946 4820
rect 37277 4811 37335 4817
rect 35360 4780 37228 4808
rect 28224 4712 32628 4740
rect 32677 4743 32735 4749
rect 28224 4700 28230 4712
rect 32677 4709 32689 4743
rect 32723 4709 32735 4743
rect 32677 4703 32735 4709
rect 28813 4675 28871 4681
rect 28813 4672 28825 4675
rect 28092 4644 28825 4672
rect 28813 4641 28825 4644
rect 28859 4672 28871 4675
rect 32125 4675 32183 4681
rect 28859 4644 31754 4672
rect 28859 4641 28871 4644
rect 28813 4635 28871 4641
rect 28166 4604 28172 4616
rect 27816 4576 28172 4604
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28629 4607 28687 4613
rect 28629 4573 28641 4607
rect 28675 4604 28687 4607
rect 29546 4604 29552 4616
rect 28675 4576 29552 4604
rect 28675 4573 28687 4576
rect 28629 4567 28687 4573
rect 29546 4564 29552 4576
rect 29604 4564 29610 4616
rect 29730 4564 29736 4616
rect 29788 4564 29794 4616
rect 30374 4564 30380 4616
rect 30432 4564 30438 4616
rect 31726 4604 31754 4644
rect 32125 4641 32137 4675
rect 32171 4672 32183 4675
rect 32398 4672 32404 4684
rect 32171 4644 32404 4672
rect 32171 4641 32183 4644
rect 32125 4635 32183 4641
rect 32398 4632 32404 4644
rect 32456 4632 32462 4684
rect 32692 4672 32720 4703
rect 34517 4675 34575 4681
rect 34517 4672 34529 4675
rect 32692 4644 34529 4672
rect 34517 4641 34529 4644
rect 34563 4641 34575 4675
rect 35360 4672 35388 4780
rect 37200 4740 37228 4780
rect 37277 4777 37289 4811
rect 37323 4808 37335 4811
rect 37550 4808 37556 4820
rect 37323 4780 37556 4808
rect 37323 4777 37335 4780
rect 37277 4771 37335 4777
rect 37550 4768 37556 4780
rect 37608 4768 37614 4820
rect 38473 4811 38531 4817
rect 38473 4777 38485 4811
rect 38519 4808 38531 4811
rect 38654 4808 38660 4820
rect 38519 4780 38660 4808
rect 38519 4777 38531 4780
rect 38473 4771 38531 4777
rect 38654 4768 38660 4780
rect 38712 4768 38718 4820
rect 40037 4811 40095 4817
rect 40037 4777 40049 4811
rect 40083 4808 40095 4811
rect 42610 4808 42616 4820
rect 40083 4780 42616 4808
rect 40083 4777 40095 4780
rect 40037 4771 40095 4777
rect 42610 4768 42616 4780
rect 42668 4768 42674 4820
rect 42702 4768 42708 4820
rect 42760 4808 42766 4820
rect 42760 4780 49280 4808
rect 42760 4768 42766 4780
rect 39114 4740 39120 4752
rect 37200 4712 39120 4740
rect 37844 4681 37872 4712
rect 39114 4700 39120 4712
rect 39172 4700 39178 4752
rect 42245 4743 42303 4749
rect 42245 4709 42257 4743
rect 42291 4740 42303 4743
rect 45738 4740 45744 4752
rect 42291 4712 42380 4740
rect 42291 4709 42303 4712
rect 42245 4703 42303 4709
rect 34517 4635 34575 4641
rect 34716 4644 35388 4672
rect 35437 4675 35495 4681
rect 31849 4607 31907 4613
rect 31849 4604 31861 4607
rect 31726 4576 31861 4604
rect 31849 4573 31861 4576
rect 31895 4604 31907 4607
rect 32769 4607 32827 4613
rect 32769 4604 32781 4607
rect 31895 4576 32781 4604
rect 31895 4573 31907 4576
rect 31849 4567 31907 4573
rect 32769 4573 32781 4576
rect 32815 4573 32827 4607
rect 33870 4604 33876 4616
rect 32769 4567 32827 4573
rect 33060 4576 33876 4604
rect 28721 4539 28779 4545
rect 28721 4505 28733 4539
rect 28767 4536 28779 4539
rect 30282 4536 30288 4548
rect 28767 4508 30288 4536
rect 28767 4505 28779 4508
rect 28721 4499 28779 4505
rect 30282 4496 30288 4508
rect 30340 4496 30346 4548
rect 31386 4496 31392 4548
rect 31444 4536 31450 4548
rect 31481 4539 31539 4545
rect 31481 4536 31493 4539
rect 31444 4508 31493 4536
rect 31444 4496 31450 4508
rect 31481 4505 31493 4508
rect 31527 4536 31539 4539
rect 32309 4539 32367 4545
rect 31527 4508 32168 4536
rect 31527 4505 31539 4508
rect 31481 4499 31539 4505
rect 32140 4480 32168 4508
rect 32309 4505 32321 4539
rect 32355 4536 32367 4539
rect 33060 4536 33088 4576
rect 33870 4564 33876 4576
rect 33928 4564 33934 4616
rect 34054 4564 34060 4616
rect 34112 4604 34118 4616
rect 34716 4604 34744 4644
rect 35437 4641 35449 4675
rect 35483 4672 35495 4675
rect 35529 4675 35587 4681
rect 35529 4672 35541 4675
rect 35483 4644 35541 4672
rect 35483 4641 35495 4644
rect 35437 4635 35495 4641
rect 35529 4641 35541 4644
rect 35575 4641 35587 4675
rect 37829 4675 37887 4681
rect 35529 4635 35587 4641
rect 35636 4644 36124 4672
rect 34112 4576 34744 4604
rect 34112 4564 34118 4576
rect 34974 4564 34980 4616
rect 35032 4564 35038 4616
rect 32355 4508 33088 4536
rect 33597 4539 33655 4545
rect 32355 4505 32367 4508
rect 32309 4499 32367 4505
rect 33597 4505 33609 4539
rect 33643 4536 33655 4539
rect 34072 4536 34100 4564
rect 33643 4508 34100 4536
rect 33643 4505 33655 4508
rect 33597 4499 33655 4505
rect 34146 4496 34152 4548
rect 34204 4496 34210 4548
rect 34992 4536 35020 4564
rect 35529 4539 35587 4545
rect 35529 4536 35541 4539
rect 34992 4508 35541 4536
rect 35529 4505 35541 4508
rect 35575 4505 35587 4539
rect 35529 4499 35587 4505
rect 28350 4468 28356 4480
rect 27724 4440 28356 4468
rect 28350 4428 28356 4440
rect 28408 4468 28414 4480
rect 29178 4468 29184 4480
rect 28408 4440 29184 4468
rect 28408 4428 28414 4440
rect 29178 4428 29184 4440
rect 29236 4428 29242 4480
rect 29365 4471 29423 4477
rect 29365 4437 29377 4471
rect 29411 4468 29423 4471
rect 29638 4468 29644 4480
rect 29411 4440 29644 4468
rect 29411 4437 29423 4440
rect 29365 4431 29423 4437
rect 29638 4428 29644 4440
rect 29696 4468 29702 4480
rect 31110 4468 31116 4480
rect 29696 4440 31116 4468
rect 29696 4428 29702 4440
rect 31110 4428 31116 4440
rect 31168 4428 31174 4480
rect 32122 4428 32128 4480
rect 32180 4428 32186 4480
rect 32217 4471 32275 4477
rect 32217 4437 32229 4471
rect 32263 4468 32275 4471
rect 33502 4468 33508 4480
rect 32263 4440 33508 4468
rect 32263 4437 32275 4440
rect 32217 4431 32275 4437
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 33870 4428 33876 4480
rect 33928 4428 33934 4480
rect 34164 4468 34192 4496
rect 35636 4468 35664 4644
rect 35894 4564 35900 4616
rect 35952 4613 35958 4616
rect 36096 4613 36124 4644
rect 37829 4641 37841 4675
rect 37875 4641 37887 4675
rect 37829 4635 37887 4641
rect 38746 4632 38752 4684
rect 38804 4632 38810 4684
rect 38838 4632 38844 4684
rect 38896 4672 38902 4684
rect 39390 4672 39396 4684
rect 38896 4644 39396 4672
rect 38896 4632 38902 4644
rect 39390 4632 39396 4644
rect 39448 4672 39454 4684
rect 40313 4675 40371 4681
rect 40313 4672 40325 4675
rect 39448 4644 40325 4672
rect 39448 4632 39454 4644
rect 40313 4641 40325 4644
rect 40359 4672 40371 4675
rect 40681 4675 40739 4681
rect 40681 4672 40693 4675
rect 40359 4644 40693 4672
rect 40359 4641 40371 4644
rect 40313 4635 40371 4641
rect 40681 4641 40693 4644
rect 40727 4641 40739 4675
rect 40681 4635 40739 4641
rect 35952 4604 35960 4613
rect 36081 4607 36139 4613
rect 35952 4576 35997 4604
rect 35952 4567 35960 4576
rect 36081 4573 36093 4607
rect 36127 4604 36139 4607
rect 36817 4607 36875 4613
rect 36817 4604 36829 4607
rect 36127 4576 36829 4604
rect 36127 4573 36139 4576
rect 36081 4567 36139 4573
rect 36817 4573 36829 4576
rect 36863 4573 36875 4607
rect 36817 4567 36875 4573
rect 38105 4607 38163 4613
rect 38105 4573 38117 4607
rect 38151 4604 38163 4607
rect 38286 4604 38292 4616
rect 38151 4576 38292 4604
rect 38151 4573 38163 4576
rect 38105 4567 38163 4573
rect 35952 4564 35958 4567
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 39577 4607 39635 4613
rect 39577 4604 39589 4607
rect 38626 4576 39589 4604
rect 35713 4539 35771 4545
rect 35713 4505 35725 4539
rect 35759 4505 35771 4539
rect 35713 4499 35771 4505
rect 35805 4539 35863 4545
rect 35805 4505 35817 4539
rect 35851 4536 35863 4539
rect 36262 4536 36268 4548
rect 35851 4508 36268 4536
rect 35851 4505 35863 4508
rect 35805 4499 35863 4505
rect 34164 4440 35664 4468
rect 35728 4468 35756 4499
rect 36262 4496 36268 4508
rect 36320 4496 36326 4548
rect 36357 4539 36415 4545
rect 36357 4505 36369 4539
rect 36403 4505 36415 4539
rect 36357 4499 36415 4505
rect 36372 4468 36400 4499
rect 36446 4496 36452 4548
rect 36504 4536 36510 4548
rect 38626 4536 38654 4576
rect 39577 4573 39589 4576
rect 39623 4573 39635 4607
rect 39577 4567 39635 4573
rect 39666 4564 39672 4616
rect 39724 4604 39730 4616
rect 39853 4607 39911 4613
rect 39853 4604 39865 4607
rect 39724 4576 39865 4604
rect 39724 4564 39730 4576
rect 39853 4573 39865 4576
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 40126 4536 40132 4548
rect 36504 4508 38654 4536
rect 39316 4508 40132 4536
rect 36504 4496 36510 4508
rect 37553 4471 37611 4477
rect 37553 4468 37565 4471
rect 35728 4440 37565 4468
rect 37553 4437 37565 4440
rect 37599 4468 37611 4471
rect 37642 4468 37648 4480
rect 37599 4440 37648 4468
rect 37599 4437 37611 4440
rect 37553 4431 37611 4437
rect 37642 4428 37648 4440
rect 37700 4428 37706 4480
rect 39316 4477 39344 4508
rect 40126 4496 40132 4508
rect 40184 4496 40190 4548
rect 40696 4536 40724 4635
rect 40862 4632 40868 4684
rect 40920 4632 40926 4684
rect 42352 4681 42380 4712
rect 44652 4712 45744 4740
rect 44652 4684 44680 4712
rect 45738 4700 45744 4712
rect 45796 4740 45802 4752
rect 46017 4743 46075 4749
rect 46017 4740 46029 4743
rect 45796 4712 46029 4740
rect 45796 4700 45802 4712
rect 46017 4709 46029 4712
rect 46063 4740 46075 4743
rect 46474 4740 46480 4752
rect 46063 4712 46480 4740
rect 46063 4709 46075 4712
rect 46017 4703 46075 4709
rect 46474 4700 46480 4712
rect 46532 4700 46538 4752
rect 42337 4675 42395 4681
rect 42337 4641 42349 4675
rect 42383 4641 42395 4675
rect 44634 4672 44640 4684
rect 42337 4635 42395 4641
rect 42536 4644 44640 4672
rect 41132 4607 41190 4613
rect 41132 4573 41144 4607
rect 41178 4604 41190 4607
rect 41598 4604 41604 4616
rect 41178 4576 41604 4604
rect 41178 4573 41190 4576
rect 41132 4567 41190 4573
rect 41598 4564 41604 4576
rect 41656 4564 41662 4616
rect 42536 4536 42564 4644
rect 43070 4564 43076 4616
rect 43128 4564 43134 4616
rect 43272 4613 43300 4644
rect 44634 4632 44640 4644
rect 44692 4632 44698 4684
rect 45922 4632 45928 4684
rect 45980 4672 45986 4684
rect 49252 4681 49280 4780
rect 49326 4768 49332 4820
rect 49384 4808 49390 4820
rect 51350 4808 51356 4820
rect 49384 4780 51356 4808
rect 49384 4768 49390 4780
rect 51350 4768 51356 4780
rect 51408 4768 51414 4820
rect 51810 4768 51816 4820
rect 51868 4808 51874 4820
rect 53834 4808 53840 4820
rect 51868 4780 53840 4808
rect 51868 4768 51874 4780
rect 53834 4768 53840 4780
rect 53892 4768 53898 4820
rect 54662 4768 54668 4820
rect 54720 4768 54726 4820
rect 56045 4811 56103 4817
rect 56045 4777 56057 4811
rect 56091 4808 56103 4811
rect 56410 4808 56416 4820
rect 56091 4780 56416 4808
rect 56091 4777 56103 4780
rect 56045 4771 56103 4777
rect 56410 4768 56416 4780
rect 56468 4768 56474 4820
rect 57882 4768 57888 4820
rect 57940 4768 57946 4820
rect 50154 4700 50160 4752
rect 50212 4740 50218 4752
rect 50212 4712 52224 4740
rect 50212 4700 50218 4712
rect 46569 4675 46627 4681
rect 46569 4672 46581 4675
rect 45980 4644 46581 4672
rect 45980 4632 45986 4644
rect 46569 4641 46581 4644
rect 46615 4641 46627 4675
rect 46569 4635 46627 4641
rect 49237 4675 49295 4681
rect 49237 4641 49249 4675
rect 49283 4672 49295 4675
rect 49283 4644 51074 4672
rect 49283 4641 49295 4644
rect 49237 4635 49295 4641
rect 43257 4607 43315 4613
rect 43257 4573 43269 4607
rect 43303 4604 43315 4607
rect 43349 4607 43407 4613
rect 43349 4604 43361 4607
rect 43303 4576 43361 4604
rect 43303 4573 43315 4576
rect 43257 4567 43315 4573
rect 43349 4573 43361 4576
rect 43395 4573 43407 4607
rect 43349 4567 43407 4573
rect 43533 4607 43591 4613
rect 43533 4573 43545 4607
rect 43579 4573 43591 4607
rect 43533 4567 43591 4573
rect 40696 4508 42564 4536
rect 42610 4496 42616 4548
rect 42668 4536 42674 4548
rect 43165 4539 43223 4545
rect 43165 4536 43177 4539
rect 42668 4508 43177 4536
rect 42668 4496 42674 4508
rect 43165 4505 43177 4508
rect 43211 4505 43223 4539
rect 43548 4536 43576 4567
rect 43806 4564 43812 4616
rect 43864 4564 43870 4616
rect 44726 4564 44732 4616
rect 44784 4564 44790 4616
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 45020 4576 45201 4604
rect 44085 4539 44143 4545
rect 44085 4536 44097 4539
rect 43548 4508 44097 4536
rect 43165 4499 43223 4505
rect 44085 4505 44097 4508
rect 44131 4505 44143 4539
rect 44085 4499 44143 4505
rect 38013 4471 38071 4477
rect 38013 4437 38025 4471
rect 38059 4468 38071 4471
rect 39301 4471 39359 4477
rect 39301 4468 39313 4471
rect 38059 4440 39313 4468
rect 38059 4437 38071 4440
rect 38013 4431 38071 4437
rect 39301 4437 39313 4440
rect 39347 4437 39359 4471
rect 39301 4431 39359 4437
rect 42242 4428 42248 4480
rect 42300 4468 42306 4480
rect 42981 4471 43039 4477
rect 42981 4468 42993 4471
rect 42300 4440 42993 4468
rect 42300 4428 42306 4440
rect 42981 4437 42993 4440
rect 43027 4437 43039 4471
rect 42981 4431 43039 4437
rect 43441 4471 43499 4477
rect 43441 4437 43453 4471
rect 43487 4468 43499 4471
rect 43530 4468 43536 4480
rect 43487 4440 43536 4468
rect 43487 4437 43499 4440
rect 43441 4431 43499 4437
rect 43530 4428 43536 4440
rect 43588 4428 43594 4480
rect 43622 4428 43628 4480
rect 43680 4428 43686 4480
rect 43714 4428 43720 4480
rect 43772 4468 43778 4480
rect 45020 4468 45048 4576
rect 45189 4573 45201 4576
rect 45235 4604 45247 4607
rect 45278 4604 45284 4616
rect 45235 4576 45284 4604
rect 45235 4573 45247 4576
rect 45189 4567 45247 4573
rect 45278 4564 45284 4576
rect 45336 4604 45342 4616
rect 46198 4604 46204 4616
rect 45336 4576 46204 4604
rect 45336 4564 45342 4576
rect 46198 4564 46204 4576
rect 46256 4604 46262 4616
rect 46842 4613 46848 4616
rect 46293 4607 46351 4613
rect 46293 4604 46305 4607
rect 46256 4576 46305 4604
rect 46256 4564 46262 4576
rect 46293 4573 46305 4576
rect 46339 4573 46351 4607
rect 46836 4604 46848 4613
rect 46803 4576 46848 4604
rect 46293 4567 46351 4573
rect 46836 4567 46848 4576
rect 46842 4564 46848 4567
rect 46900 4564 46906 4616
rect 47762 4564 47768 4616
rect 47820 4604 47826 4616
rect 48225 4607 48283 4613
rect 48225 4604 48237 4607
rect 47820 4576 48237 4604
rect 47820 4564 47826 4576
rect 48225 4573 48237 4576
rect 48271 4604 48283 4607
rect 49513 4607 49571 4613
rect 49513 4604 49525 4607
rect 48271 4576 49525 4604
rect 48271 4573 48283 4576
rect 48225 4567 48283 4573
rect 49513 4573 49525 4576
rect 49559 4604 49571 4607
rect 49697 4607 49755 4613
rect 49697 4604 49709 4607
rect 49559 4576 49709 4604
rect 49559 4573 49571 4576
rect 49513 4567 49571 4573
rect 49697 4573 49709 4576
rect 49743 4573 49755 4607
rect 49697 4567 49755 4573
rect 49878 4564 49884 4616
rect 49936 4564 49942 4616
rect 50154 4564 50160 4616
rect 50212 4564 50218 4616
rect 51046 4604 51074 4644
rect 52196 4613 52224 4712
rect 53650 4700 53656 4752
rect 53708 4740 53714 4752
rect 54680 4740 54708 4768
rect 57900 4740 57928 4768
rect 53708 4712 54708 4740
rect 56060 4712 57928 4740
rect 53708 4700 53714 4712
rect 55048 4644 55904 4672
rect 51905 4607 51963 4613
rect 51905 4604 51917 4607
rect 51046 4576 51917 4604
rect 51905 4573 51917 4576
rect 51951 4573 51963 4607
rect 51905 4567 51963 4573
rect 52181 4607 52239 4613
rect 52181 4573 52193 4607
rect 52227 4604 52239 4607
rect 53006 4604 53012 4616
rect 52227 4576 53012 4604
rect 52227 4573 52239 4576
rect 52181 4567 52239 4573
rect 51810 4536 51816 4548
rect 45112 4508 51816 4536
rect 45112 4480 45140 4508
rect 51810 4496 51816 4508
rect 51868 4496 51874 4548
rect 43772 4440 45048 4468
rect 43772 4428 43778 4440
rect 45094 4428 45100 4480
rect 45152 4428 45158 4480
rect 45462 4428 45468 4480
rect 45520 4468 45526 4480
rect 45557 4471 45615 4477
rect 45557 4468 45569 4471
rect 45520 4440 45569 4468
rect 45520 4428 45526 4440
rect 45557 4437 45569 4440
rect 45603 4468 45615 4471
rect 46658 4468 46664 4480
rect 45603 4440 46664 4468
rect 45603 4437 45615 4440
rect 45557 4431 45615 4437
rect 46658 4428 46664 4440
rect 46716 4428 46722 4480
rect 47118 4428 47124 4480
rect 47176 4468 47182 4480
rect 47854 4468 47860 4480
rect 47176 4440 47860 4468
rect 47176 4428 47182 4440
rect 47854 4428 47860 4440
rect 47912 4428 47918 4480
rect 47946 4428 47952 4480
rect 48004 4428 48010 4480
rect 48682 4428 48688 4480
rect 48740 4468 48746 4480
rect 49694 4468 49700 4480
rect 48740 4440 49700 4468
rect 48740 4428 48746 4440
rect 49694 4428 49700 4440
rect 49752 4428 49758 4480
rect 49789 4471 49847 4477
rect 49789 4437 49801 4471
rect 49835 4468 49847 4471
rect 50062 4468 50068 4480
rect 49835 4440 50068 4468
rect 49835 4437 49847 4440
rect 49789 4431 49847 4437
rect 50062 4428 50068 4440
rect 50120 4428 50126 4480
rect 51920 4468 51948 4567
rect 53006 4564 53012 4576
rect 53064 4564 53070 4616
rect 53742 4564 53748 4616
rect 53800 4564 53806 4616
rect 54846 4564 54852 4616
rect 54904 4604 54910 4616
rect 55048 4613 55076 4644
rect 55876 4613 55904 4644
rect 56060 4613 56088 4712
rect 56318 4632 56324 4684
rect 56376 4632 56382 4684
rect 56686 4632 56692 4684
rect 56744 4672 56750 4684
rect 56873 4675 56931 4681
rect 56873 4672 56885 4675
rect 56744 4644 56885 4672
rect 56744 4632 56750 4644
rect 56873 4641 56885 4644
rect 56919 4641 56931 4675
rect 56873 4635 56931 4641
rect 55033 4607 55091 4613
rect 55033 4604 55045 4607
rect 54904 4576 55045 4604
rect 54904 4564 54910 4576
rect 55033 4573 55045 4576
rect 55079 4573 55091 4607
rect 55033 4567 55091 4573
rect 55769 4607 55827 4613
rect 55769 4573 55781 4607
rect 55815 4573 55827 4607
rect 55769 4567 55827 4573
rect 55861 4607 55919 4613
rect 55861 4573 55873 4607
rect 55907 4573 55919 4607
rect 55861 4567 55919 4573
rect 56045 4607 56103 4613
rect 56045 4573 56057 4607
rect 56091 4573 56103 4607
rect 56045 4567 56103 4573
rect 52448 4539 52506 4545
rect 52448 4505 52460 4539
rect 52494 4536 52506 4539
rect 52638 4536 52644 4548
rect 52494 4508 52644 4536
rect 52494 4505 52506 4508
rect 52448 4499 52506 4505
rect 52638 4496 52644 4508
rect 52696 4496 52702 4548
rect 55784 4536 55812 4567
rect 57146 4564 57152 4616
rect 57204 4564 57210 4616
rect 57790 4536 57796 4548
rect 55784 4508 57796 4536
rect 57790 4496 57796 4508
rect 57848 4496 57854 4548
rect 58345 4539 58403 4545
rect 58345 4505 58357 4539
rect 58391 4536 58403 4539
rect 58618 4536 58624 4548
rect 58391 4508 58624 4536
rect 58391 4505 58403 4508
rect 58345 4499 58403 4505
rect 58618 4496 58624 4508
rect 58676 4496 58682 4548
rect 53190 4468 53196 4480
rect 51920 4440 53196 4468
rect 53190 4428 53196 4440
rect 53248 4428 53254 4480
rect 53561 4471 53619 4477
rect 53561 4437 53573 4471
rect 53607 4468 53619 4471
rect 54110 4468 54116 4480
rect 53607 4440 54116 4468
rect 53607 4437 53619 4440
rect 53561 4431 53619 4437
rect 54110 4428 54116 4440
rect 54168 4428 54174 4480
rect 54294 4428 54300 4480
rect 54352 4428 54358 4480
rect 55214 4428 55220 4480
rect 55272 4468 55278 4480
rect 55585 4471 55643 4477
rect 55585 4468 55597 4471
rect 55272 4440 55597 4468
rect 55272 4428 55278 4440
rect 55585 4437 55597 4440
rect 55631 4437 55643 4471
rect 55585 4431 55643 4437
rect 1104 4378 59040 4400
rect 1104 4326 15394 4378
rect 15446 4326 15458 4378
rect 15510 4326 15522 4378
rect 15574 4326 15586 4378
rect 15638 4326 15650 4378
rect 15702 4326 29838 4378
rect 29890 4326 29902 4378
rect 29954 4326 29966 4378
rect 30018 4326 30030 4378
rect 30082 4326 30094 4378
rect 30146 4326 44282 4378
rect 44334 4326 44346 4378
rect 44398 4326 44410 4378
rect 44462 4326 44474 4378
rect 44526 4326 44538 4378
rect 44590 4326 58726 4378
rect 58778 4326 58790 4378
rect 58842 4326 58854 4378
rect 58906 4326 58918 4378
rect 58970 4326 58982 4378
rect 59034 4326 59040 4378
rect 1104 4304 59040 4326
rect 2608 4236 2912 4264
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2222 4128 2228 4140
rect 2087 4100 2228 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2608 4128 2636 4236
rect 2884 4208 2912 4236
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 6052 4236 6377 4264
rect 6052 4224 6058 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 6365 4227 6423 4233
rect 7484 4236 10640 4264
rect 2676 4199 2734 4205
rect 2676 4165 2688 4199
rect 2722 4196 2734 4199
rect 2774 4196 2780 4208
rect 2722 4168 2780 4196
rect 2722 4165 2734 4168
rect 2676 4159 2734 4165
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 2866 4156 2872 4208
rect 2924 4156 2930 4208
rect 3988 4168 4384 4196
rect 3988 4140 4016 4168
rect 2363 4100 2636 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4356 4137 4384 4168
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 4617 4199 4675 4205
rect 4617 4196 4629 4199
rect 4488 4168 4629 4196
rect 4488 4156 4494 4168
rect 4617 4165 4629 4168
rect 4663 4165 4675 4199
rect 6454 4196 6460 4208
rect 4617 4159 4675 4165
rect 5460 4168 6460 4196
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 3528 4060 3556 4088
rect 4080 4060 4108 4091
rect 3528 4032 4108 4060
rect 2409 4023 2467 4029
rect 1578 3952 1584 4004
rect 1636 3952 1642 4004
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2038 3924 2044 3936
rect 1903 3896 2044 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 2222 3924 2228 3936
rect 2179 3896 2228 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2424 3924 2452 4023
rect 3786 3992 3792 4004
rect 3344 3964 3792 3992
rect 3344 3936 3372 3964
rect 3786 3952 3792 3964
rect 3844 3992 3850 4004
rect 4724 3992 4752 4091
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5350 4128 5356 4140
rect 4856 4100 5356 4128
rect 4856 4088 4862 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5460 4060 5488 4168
rect 6454 4156 6460 4168
rect 6512 4196 6518 4208
rect 7484 4196 7512 4236
rect 7834 4196 7840 4208
rect 6512 4168 7512 4196
rect 7576 4168 7840 4196
rect 6512 4156 6518 4168
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5684 4100 5917 4128
rect 5684 4088 5690 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 6236 4100 7113 4128
rect 6236 4088 6242 4100
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7576 4137 7604 4168
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 8481 4199 8539 4205
rect 8481 4165 8493 4199
rect 8527 4196 8539 4199
rect 9766 4196 9772 4208
rect 8527 4168 9772 4196
rect 8527 4165 8539 4168
rect 8481 4159 8539 4165
rect 9766 4156 9772 4168
rect 9824 4196 9830 4208
rect 10502 4196 10508 4208
rect 9824 4168 10508 4196
rect 9824 4156 9830 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 10612 4196 10640 4236
rect 10962 4224 10968 4276
rect 11020 4224 11026 4276
rect 12434 4224 12440 4276
rect 12492 4224 12498 4276
rect 14642 4264 14648 4276
rect 13188 4236 13676 4264
rect 12452 4196 12480 4224
rect 10612 4168 12480 4196
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 5040 4032 5488 4060
rect 5040 4020 5046 4032
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6328 4032 6929 4060
rect 6328 4020 6334 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 3844 3964 4752 3992
rect 5736 3992 5764 4020
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 5736 3964 7205 3992
rect 3844 3952 3850 3964
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7760 3992 7788 4091
rect 7926 4088 7932 4140
rect 7984 4088 7990 4140
rect 8205 4131 8263 4137
rect 8108 4121 8166 4127
rect 8108 4087 8120 4121
rect 8154 4087 8166 4121
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8108 4081 8166 4087
rect 8128 4004 8156 4081
rect 7760 3964 7880 3992
rect 7193 3955 7251 3961
rect 7852 3936 7880 3964
rect 8110 3952 8116 4004
rect 8168 3952 8174 4004
rect 8220 3992 8248 4091
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8754 4128 8760 4140
rect 8352 4100 8760 4128
rect 8352 4088 8358 4100
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9539 4100 9689 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9784 4100 11652 4128
rect 8386 4020 8392 4072
rect 8444 4020 8450 4072
rect 8570 4020 8576 4072
rect 8628 4020 8634 4072
rect 8662 3992 8668 4004
rect 8220 3964 8668 3992
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 9784 3992 9812 4100
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9916 4032 10241 4060
rect 9916 4020 9922 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11112 4032 11529 4060
rect 11112 4020 11118 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11624 4060 11652 4100
rect 11624 4032 12434 4060
rect 11517 4023 11575 4029
rect 12406 3992 12434 4032
rect 12621 3995 12679 4001
rect 12621 3992 12633 3995
rect 8772 3964 9812 3992
rect 11256 3964 12296 3992
rect 12406 3964 12633 3992
rect 3050 3924 3056 3936
rect 2424 3896 3056 3924
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 7558 3884 7564 3936
rect 7616 3884 7622 3936
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8772 3924 8800 3964
rect 7892 3896 8800 3924
rect 7892 3884 7898 3896
rect 9214 3884 9220 3936
rect 9272 3884 9278 3936
rect 9490 3884 9496 3936
rect 9548 3884 9554 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11256 3933 11284 3964
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10652 3896 11253 3924
rect 10652 3884 10658 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 12158 3884 12164 3936
rect 12216 3884 12222 3936
rect 12268 3924 12296 3964
rect 12621 3961 12633 3964
rect 12667 3961 12679 3995
rect 12621 3955 12679 3961
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12268 3896 12449 3924
rect 12437 3893 12449 3896
rect 12483 3924 12495 3927
rect 13188 3924 13216 4236
rect 13538 4156 13544 4208
rect 13596 4156 13602 4208
rect 13446 4137 13452 4140
rect 13444 4091 13452 4137
rect 13504 4128 13510 4140
rect 13648 4137 13676 4236
rect 13832 4236 14648 4264
rect 13832 4205 13860 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 14734 4224 14740 4276
rect 14792 4264 14798 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14792 4236 15025 4264
rect 14792 4224 14798 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 15120 4236 15516 4264
rect 13817 4199 13875 4205
rect 13817 4165 13829 4199
rect 13863 4165 13875 4199
rect 14274 4196 14280 4208
rect 13817 4159 13875 4165
rect 14016 4168 14280 4196
rect 13633 4131 13691 4137
rect 13504 4100 13544 4128
rect 13446 4088 13452 4091
rect 13504 4088 13510 4100
rect 13633 4097 13645 4131
rect 13679 4128 13691 4131
rect 13915 4131 13973 4137
rect 13679 4100 13860 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 12483 3896 13216 3924
rect 13280 3924 13308 4023
rect 13722 4020 13728 4072
rect 13780 4020 13786 4072
rect 13832 4060 13860 4100
rect 13915 4097 13927 4131
rect 13961 4128 13973 4131
rect 14016 4128 14044 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15120 4196 15148 4236
rect 14844 4168 15148 4196
rect 13961 4100 14044 4128
rect 13961 4097 13973 4100
rect 13915 4091 13973 4097
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14844 4069 14872 4168
rect 15194 4156 15200 4208
rect 15252 4196 15258 4208
rect 15252 4168 15327 4196
rect 15252 4156 15258 4168
rect 14918 4088 14924 4140
rect 14976 4088 14982 4140
rect 15102 4088 15108 4140
rect 15160 4088 15166 4140
rect 15299 4127 15327 4168
rect 15284 4121 15342 4127
rect 15284 4087 15296 4121
rect 15330 4087 15342 4121
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15488 4137 15516 4236
rect 20898 4224 20904 4276
rect 20956 4264 20962 4276
rect 20993 4267 21051 4273
rect 20993 4264 21005 4267
rect 20956 4236 21005 4264
rect 20956 4224 20962 4236
rect 20993 4233 21005 4236
rect 21039 4233 21051 4267
rect 20993 4227 21051 4233
rect 21100 4236 22416 4264
rect 15657 4199 15715 4205
rect 15657 4165 15669 4199
rect 15703 4196 15715 4199
rect 16390 4196 16396 4208
rect 15703 4168 16396 4196
rect 15703 4165 15715 4168
rect 15657 4159 15715 4165
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 16500 4168 17715 4196
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 16114 4128 16120 4140
rect 15519 4100 16120 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 16114 4088 16120 4100
rect 16172 4128 16178 4140
rect 16500 4128 16528 4168
rect 16172 4100 16528 4128
rect 16172 4088 16178 4100
rect 17586 4088 17592 4140
rect 17644 4088 17650 4140
rect 17687 4128 17715 4168
rect 17862 4156 17868 4208
rect 17920 4156 17926 4208
rect 18138 4156 18144 4208
rect 18196 4156 18202 4208
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 21100 4196 21128 4236
rect 21726 4196 21732 4208
rect 18932 4168 21128 4196
rect 21192 4168 21732 4196
rect 18932 4156 18938 4168
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17687 4100 18337 4128
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4097 18475 4131
rect 18417 4091 18475 4097
rect 15284 4081 15342 4087
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 13832 4032 14841 4060
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16022 4060 16028 4072
rect 15611 4032 16028 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16298 4020 16304 4072
rect 16356 4020 16362 4072
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 16448 4032 17233 4060
rect 16448 4020 16454 4032
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17773 4063 17831 4069
rect 17773 4029 17785 4063
rect 17819 4060 17831 4063
rect 18046 4060 18052 4072
rect 17819 4032 18052 4060
rect 17819 4029 17831 4032
rect 17773 4023 17831 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13412 3964 14105 3992
rect 13412 3952 13418 3964
rect 14093 3961 14105 3964
rect 14139 3961 14151 3995
rect 14093 3955 14151 3961
rect 14200 3964 14504 3992
rect 14200 3924 14228 3964
rect 13280 3896 14228 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 14476 3924 14504 3964
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 14792 3964 15761 3992
rect 14792 3952 14798 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 17405 3995 17463 4001
rect 17405 3992 17417 3995
rect 15749 3955 15807 3961
rect 15856 3964 17417 3992
rect 15856 3924 15884 3964
rect 17405 3961 17417 3964
rect 17451 3961 17463 3995
rect 17405 3955 17463 3961
rect 18141 3995 18199 4001
rect 18141 3961 18153 3995
rect 18187 3992 18199 3995
rect 18230 3992 18236 4004
rect 18187 3964 18236 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 14476 3896 15884 3924
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 15988 3896 16681 3924
rect 15988 3884 15994 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 17368 3896 17601 3924
rect 17368 3884 17374 3896
rect 17589 3893 17601 3896
rect 17635 3893 17647 3927
rect 18340 3924 18368 4091
rect 18432 4060 18460 4091
rect 18506 4088 18512 4140
rect 18564 4137 18570 4140
rect 18564 4128 18572 4137
rect 18564 4100 18609 4128
rect 18564 4091 18572 4100
rect 18564 4088 18570 4091
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 19484 4100 19717 4128
rect 19484 4088 19490 4100
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 19886 4088 19892 4140
rect 19944 4088 19950 4140
rect 19978 4088 19984 4140
rect 20036 4088 20042 4140
rect 20070 4088 20076 4140
rect 20128 4137 20134 4140
rect 21192 4137 21220 4168
rect 21468 4137 21496 4168
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 22278 4196 22284 4208
rect 22066 4168 22284 4196
rect 20128 4128 20136 4137
rect 21177 4131 21235 4137
rect 20128 4100 20173 4128
rect 20128 4091 20136 4100
rect 21177 4097 21189 4131
rect 21223 4097 21235 4131
rect 21177 4091 21235 4097
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4097 21511 4131
rect 21453 4091 21511 4097
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4097 21695 4131
rect 21637 4091 21695 4097
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4128 21971 4131
rect 22066 4128 22094 4168
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 22388 4196 22416 4236
rect 23382 4224 23388 4276
rect 23440 4224 23446 4276
rect 27890 4264 27896 4276
rect 24136 4236 27896 4264
rect 24136 4196 24164 4236
rect 27890 4224 27896 4236
rect 27948 4224 27954 4276
rect 27985 4267 28043 4273
rect 27985 4233 27997 4267
rect 28031 4233 28043 4267
rect 27985 4227 28043 4233
rect 22388 4168 24164 4196
rect 24210 4156 24216 4208
rect 24268 4196 24274 4208
rect 24581 4199 24639 4205
rect 24268 4168 24440 4196
rect 24268 4156 24274 4168
rect 22186 4137 22192 4140
rect 21959 4100 22094 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 22180 4091 22192 4137
rect 22244 4128 22250 4140
rect 22244 4100 22280 4128
rect 20128 4088 20134 4091
rect 19058 4060 19064 4072
rect 18432 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 19843 4032 20361 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 21376 4060 21404 4091
rect 21542 4060 21548 4072
rect 21376 4032 21548 4060
rect 20349 4023 20407 4029
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 21652 4060 21680 4091
rect 22186 4088 22192 4091
rect 22244 4088 22250 4100
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 24305 4131 24363 4137
rect 24305 4128 24317 4131
rect 23532 4100 24317 4128
rect 23532 4088 23538 4100
rect 24305 4097 24317 4100
rect 24351 4097 24363 4131
rect 24412 4128 24440 4168
rect 24581 4165 24593 4199
rect 24627 4196 24639 4199
rect 24627 4168 27844 4196
rect 24627 4165 24639 4168
rect 24581 4159 24639 4165
rect 27816 4152 27844 4168
rect 28000 4152 28028 4227
rect 28074 4224 28080 4276
rect 28132 4264 28138 4276
rect 30193 4267 30251 4273
rect 30193 4264 30205 4267
rect 28132 4236 30205 4264
rect 28132 4224 28138 4236
rect 30193 4233 30205 4236
rect 30239 4233 30251 4267
rect 30193 4227 30251 4233
rect 30282 4224 30288 4276
rect 30340 4224 30346 4276
rect 30374 4224 30380 4276
rect 30432 4224 30438 4276
rect 32122 4224 32128 4276
rect 32180 4264 32186 4276
rect 33410 4264 33416 4276
rect 32180 4236 33416 4264
rect 32180 4224 32186 4236
rect 33410 4224 33416 4236
rect 33468 4224 33474 4276
rect 33502 4224 33508 4276
rect 33560 4264 33566 4276
rect 33962 4264 33968 4276
rect 33560 4236 33968 4264
rect 33560 4224 33566 4236
rect 33962 4224 33968 4236
rect 34020 4264 34026 4276
rect 34241 4267 34299 4273
rect 34241 4264 34253 4267
rect 34020 4236 34253 4264
rect 34020 4224 34026 4236
rect 34241 4233 34253 4236
rect 34287 4233 34299 4267
rect 34241 4227 34299 4233
rect 35066 4224 35072 4276
rect 35124 4264 35130 4276
rect 35894 4264 35900 4276
rect 35124 4236 35900 4264
rect 35124 4224 35130 4236
rect 35894 4224 35900 4236
rect 35952 4264 35958 4276
rect 36265 4267 36323 4273
rect 36265 4264 36277 4267
rect 35952 4236 36277 4264
rect 35952 4224 35958 4236
rect 36265 4233 36277 4236
rect 36311 4264 36323 4267
rect 39298 4264 39304 4276
rect 36311 4236 37596 4264
rect 36311 4233 36323 4236
rect 36265 4227 36323 4233
rect 28537 4199 28595 4205
rect 28537 4165 28549 4199
rect 28583 4196 28595 4199
rect 28583 4168 28994 4196
rect 28583 4165 28595 4168
rect 28537 4159 28595 4165
rect 24946 4137 24952 4140
rect 24913 4131 24952 4137
rect 24913 4128 24925 4131
rect 24412 4100 24925 4128
rect 24305 4091 24363 4097
rect 24913 4097 24925 4100
rect 24913 4091 24952 4097
rect 24946 4088 24952 4091
rect 25004 4088 25010 4140
rect 25038 4088 25044 4140
rect 25096 4088 25102 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4097 25191 4131
rect 25133 4091 25191 4097
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 25406 4128 25412 4140
rect 25363 4100 25412 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 21726 4060 21732 4072
rect 21652 4032 21732 4060
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 23308 4032 23949 4060
rect 18690 3952 18696 4004
rect 18748 3992 18754 4004
rect 23308 4001 23336 4032
rect 23937 4029 23949 4032
rect 23983 4029 23995 4063
rect 23937 4023 23995 4029
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 24397 4063 24455 4069
rect 24397 4060 24409 4063
rect 24176 4032 24409 4060
rect 24176 4020 24182 4032
rect 24397 4029 24409 4032
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25148 4060 25176 4091
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 26786 4088 26792 4140
rect 26844 4088 26850 4140
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 27522 4088 27528 4140
rect 27580 4088 27586 4140
rect 27816 4124 28028 4152
rect 28166 4088 28172 4140
rect 28224 4088 28230 4140
rect 28350 4137 28356 4140
rect 28348 4128 28356 4137
rect 28311 4100 28356 4128
rect 28348 4091 28356 4100
rect 28350 4088 28356 4091
rect 28408 4088 28414 4140
rect 28442 4088 28448 4140
rect 28500 4088 28506 4140
rect 24820 4032 25176 4060
rect 25225 4063 25283 4069
rect 24820 4020 24826 4032
rect 23293 3995 23351 4001
rect 18748 3964 21772 3992
rect 18748 3952 18754 3964
rect 19886 3924 19892 3936
rect 18340 3896 19892 3924
rect 17589 3887 17647 3893
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 21358 3884 21364 3936
rect 21416 3884 21422 3936
rect 21634 3884 21640 3936
rect 21692 3884 21698 3936
rect 21744 3924 21772 3964
rect 23293 3961 23305 3995
rect 23339 3961 23351 3995
rect 23293 3955 23351 3961
rect 24121 3927 24179 3933
rect 24121 3924 24133 3927
rect 21744 3896 24133 3924
rect 24121 3893 24133 3896
rect 24167 3893 24179 3927
rect 24121 3887 24179 3893
rect 24394 3884 24400 3936
rect 24452 3884 24458 3936
rect 24964 3924 24992 4032
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25271 4032 25973 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 27246 4060 27252 4072
rect 25961 4023 26019 4029
rect 26436 4032 27252 4060
rect 25038 3952 25044 4004
rect 25096 3992 25102 4004
rect 25409 3995 25467 4001
rect 25409 3992 25421 3995
rect 25096 3964 25421 3992
rect 25096 3952 25102 3964
rect 25409 3961 25421 3964
rect 25455 3961 25467 3995
rect 25409 3955 25467 3961
rect 26436 3933 26464 4032
rect 27246 4020 27252 4032
rect 27304 4060 27310 4072
rect 27433 4063 27491 4069
rect 27433 4060 27445 4063
rect 27304 4032 27445 4060
rect 27304 4020 27310 4032
rect 27433 4029 27445 4032
rect 27479 4029 27491 4063
rect 27540 4060 27568 4088
rect 27801 4063 27859 4069
rect 27801 4060 27813 4063
rect 27540 4032 27813 4060
rect 27433 4023 27491 4029
rect 27801 4029 27813 4032
rect 27847 4029 27859 4063
rect 28552 4060 28580 4159
rect 28718 4088 28724 4140
rect 28776 4088 28782 4140
rect 28966 4128 28994 4168
rect 29178 4156 29184 4208
rect 29236 4196 29242 4208
rect 29236 4168 29592 4196
rect 29236 4156 29242 4168
rect 29564 4128 29592 4168
rect 29638 4156 29644 4208
rect 29696 4196 29702 4208
rect 29917 4199 29975 4205
rect 29917 4196 29929 4199
rect 29696 4168 29929 4196
rect 29696 4156 29702 4168
rect 29917 4165 29929 4168
rect 29963 4165 29975 4199
rect 29917 4159 29975 4165
rect 30101 4199 30159 4205
rect 30101 4165 30113 4199
rect 30147 4196 30159 4199
rect 30300 4196 30328 4224
rect 30147 4168 30328 4196
rect 30392 4196 30420 4224
rect 33260 4199 33318 4205
rect 30392 4168 30788 4196
rect 30147 4165 30159 4168
rect 30101 4159 30159 4165
rect 29825 4131 29883 4137
rect 28966 4100 29500 4128
rect 29564 4121 29771 4128
rect 29564 4100 29709 4121
rect 27801 4023 27859 4029
rect 27908 4032 28580 4060
rect 28629 4063 28687 4069
rect 27154 3952 27160 4004
rect 27212 3952 27218 4004
rect 27448 3992 27476 4023
rect 27908 3992 27936 4032
rect 28629 4029 28641 4063
rect 28675 4060 28687 4063
rect 29365 4063 29423 4069
rect 29365 4060 29377 4063
rect 28675 4032 29377 4060
rect 28675 4029 28687 4032
rect 28629 4023 28687 4029
rect 29365 4029 29377 4032
rect 29411 4029 29423 4063
rect 29365 4023 29423 4029
rect 27448 3964 27936 3992
rect 28074 3952 28080 4004
rect 28132 3992 28138 4004
rect 28132 3964 28580 3992
rect 28132 3952 28138 3964
rect 26421 3927 26479 3933
rect 26421 3924 26433 3927
rect 24964 3896 26433 3924
rect 26421 3893 26433 3896
rect 26467 3893 26479 3927
rect 26421 3887 26479 3893
rect 26602 3884 26608 3936
rect 26660 3884 26666 3936
rect 28552 3924 28580 3964
rect 28810 3952 28816 4004
rect 28868 3952 28874 4004
rect 29472 3992 29500 4100
rect 29697 4087 29709 4100
rect 29743 4090 29771 4121
rect 29825 4097 29837 4131
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 29743 4087 29755 4090
rect 29697 4081 29755 4087
rect 29840 4060 29868 4091
rect 30006 4088 30012 4140
rect 30064 4128 30070 4140
rect 30377 4131 30435 4137
rect 30377 4128 30389 4131
rect 30064 4100 30389 4128
rect 30064 4088 30070 4100
rect 30377 4097 30389 4100
rect 30423 4097 30435 4131
rect 30377 4091 30435 4097
rect 30650 4088 30656 4140
rect 30708 4088 30714 4140
rect 30760 4137 30788 4168
rect 33260 4165 33272 4199
rect 33306 4196 33318 4199
rect 33870 4196 33876 4208
rect 33306 4168 33876 4196
rect 33306 4165 33318 4168
rect 33260 4159 33318 4165
rect 33870 4156 33876 4168
rect 33928 4156 33934 4208
rect 34790 4205 34796 4208
rect 34784 4196 34796 4205
rect 34751 4168 34796 4196
rect 34784 4159 34796 4168
rect 34790 4156 34796 4159
rect 34848 4156 34854 4208
rect 30745 4131 30803 4137
rect 30745 4097 30757 4131
rect 30791 4097 30803 4131
rect 30745 4091 30803 4097
rect 30929 4131 30987 4137
rect 30929 4097 30941 4131
rect 30975 4128 30987 4131
rect 31205 4131 31263 4137
rect 31205 4128 31217 4131
rect 30975 4100 31217 4128
rect 30975 4097 30987 4100
rect 30929 4091 30987 4097
rect 31205 4097 31217 4100
rect 31251 4097 31263 4131
rect 31205 4091 31263 4097
rect 32140 4100 33456 4128
rect 29840 4032 30420 4060
rect 30392 4004 30420 4032
rect 30466 4020 30472 4072
rect 30524 4020 30530 4072
rect 30944 4060 30972 4091
rect 30576 4032 30972 4060
rect 29638 3992 29644 4004
rect 29472 3964 29644 3992
rect 29638 3952 29644 3964
rect 29696 3952 29702 4004
rect 29730 3952 29736 4004
rect 29788 3992 29794 4004
rect 30101 3995 30159 4001
rect 30101 3992 30113 3995
rect 29788 3964 30113 3992
rect 29788 3952 29794 3964
rect 30101 3961 30113 3964
rect 30147 3961 30159 3995
rect 30101 3955 30159 3961
rect 30374 3952 30380 4004
rect 30432 3952 30438 4004
rect 30576 3924 30604 4032
rect 32140 4001 32168 4100
rect 33428 4060 33456 4100
rect 33502 4088 33508 4140
rect 33560 4128 33566 4140
rect 34517 4131 34575 4137
rect 34517 4128 34529 4131
rect 33560 4100 34529 4128
rect 33560 4088 33566 4100
rect 34517 4097 34529 4100
rect 34563 4097 34575 4131
rect 34517 4091 34575 4097
rect 36354 4088 36360 4140
rect 36412 4088 36418 4140
rect 36538 4088 36544 4140
rect 36596 4128 36602 4140
rect 36633 4131 36691 4137
rect 36633 4128 36645 4131
rect 36596 4100 36645 4128
rect 36596 4088 36602 4100
rect 36633 4097 36645 4100
rect 36679 4097 36691 4131
rect 36633 4091 36691 4097
rect 36817 4131 36875 4137
rect 36817 4097 36829 4131
rect 36863 4128 36875 4131
rect 37277 4131 37335 4137
rect 37277 4128 37289 4131
rect 36863 4100 37289 4128
rect 36863 4097 36875 4100
rect 36817 4091 36875 4097
rect 37277 4097 37289 4100
rect 37323 4097 37335 4131
rect 37568 4128 37596 4236
rect 38304 4236 39304 4264
rect 37642 4156 37648 4208
rect 37700 4196 37706 4208
rect 38304 4205 38332 4236
rect 39298 4224 39304 4236
rect 39356 4264 39362 4276
rect 44634 4264 44640 4276
rect 39356 4236 39988 4264
rect 39356 4224 39362 4236
rect 38289 4199 38347 4205
rect 38289 4196 38301 4199
rect 37700 4168 38301 4196
rect 37700 4156 37706 4168
rect 38289 4165 38301 4168
rect 38335 4165 38347 4199
rect 38289 4159 38347 4165
rect 38378 4156 38384 4208
rect 38436 4196 38442 4208
rect 38473 4199 38531 4205
rect 38473 4196 38485 4199
rect 38436 4168 38485 4196
rect 38436 4156 38442 4168
rect 38473 4165 38485 4168
rect 38519 4165 38531 4199
rect 38473 4159 38531 4165
rect 38102 4137 38108 4140
rect 38069 4131 38108 4137
rect 38069 4128 38081 4131
rect 37568 4100 38081 4128
rect 37277 4091 37335 4097
rect 38069 4097 38081 4100
rect 38069 4091 38108 4097
rect 38102 4088 38108 4091
rect 38160 4088 38166 4140
rect 38194 4088 38200 4140
rect 38252 4088 38258 4140
rect 38565 4131 38623 4137
rect 38565 4097 38577 4131
rect 38611 4128 38623 4131
rect 38654 4128 38660 4140
rect 38611 4100 38660 4128
rect 38611 4097 38623 4100
rect 38565 4091 38623 4097
rect 38654 4088 38660 4100
rect 38712 4088 38718 4140
rect 38749 4131 38807 4137
rect 38749 4097 38761 4131
rect 38795 4128 38807 4131
rect 38841 4131 38899 4137
rect 38841 4128 38853 4131
rect 38795 4100 38853 4128
rect 38795 4097 38807 4100
rect 38749 4091 38807 4097
rect 38841 4097 38853 4100
rect 38887 4097 38899 4131
rect 38841 4091 38899 4097
rect 38948 4100 39620 4128
rect 33597 4063 33655 4069
rect 33597 4060 33609 4063
rect 33428 4032 33609 4060
rect 33597 4029 33609 4032
rect 33643 4029 33655 4063
rect 36262 4060 36268 4072
rect 33597 4023 33655 4029
rect 35912 4032 36268 4060
rect 35912 4001 35940 4032
rect 36262 4020 36268 4032
rect 36320 4060 36326 4072
rect 36906 4060 36912 4072
rect 36320 4032 36912 4060
rect 36320 4020 36326 4032
rect 36906 4020 36912 4032
rect 36964 4020 36970 4072
rect 37921 4063 37979 4069
rect 37921 4029 37933 4063
rect 37967 4060 37979 4063
rect 38381 4063 38439 4069
rect 38381 4060 38393 4063
rect 37967 4032 38393 4060
rect 37967 4029 37979 4032
rect 37921 4023 37979 4029
rect 38381 4029 38393 4032
rect 38427 4029 38439 4063
rect 38948 4060 38976 4100
rect 38381 4023 38439 4029
rect 38488 4032 38976 4060
rect 39485 4063 39543 4069
rect 32125 3995 32183 4001
rect 32125 3961 32137 3995
rect 32171 3961 32183 3995
rect 32125 3955 32183 3961
rect 35897 3995 35955 4001
rect 35897 3961 35909 3995
rect 35943 3961 35955 3995
rect 35897 3955 35955 3961
rect 36541 3995 36599 4001
rect 36541 3961 36553 3995
rect 36587 3992 36599 3995
rect 38488 3992 38516 4032
rect 39485 4029 39497 4063
rect 39531 4029 39543 4063
rect 39592 4060 39620 4100
rect 39758 4088 39764 4140
rect 39816 4088 39822 4140
rect 39960 4128 39988 4236
rect 40052 4236 44640 4264
rect 40052 4205 40080 4236
rect 44634 4224 44640 4236
rect 44692 4224 44698 4276
rect 44818 4224 44824 4276
rect 44876 4264 44882 4276
rect 44876 4236 45416 4264
rect 44876 4224 44882 4236
rect 40037 4199 40095 4205
rect 40037 4165 40049 4199
rect 40083 4165 40095 4199
rect 40037 4159 40095 4165
rect 40126 4156 40132 4208
rect 40184 4156 40190 4208
rect 41233 4199 41291 4205
rect 41233 4196 41245 4199
rect 40328 4168 41245 4196
rect 40328 4137 40356 4168
rect 41233 4165 41245 4168
rect 41279 4165 41291 4199
rect 41233 4159 41291 4165
rect 40313 4131 40371 4137
rect 40313 4128 40325 4131
rect 39960 4100 40325 4128
rect 40313 4097 40325 4100
rect 40359 4097 40371 4131
rect 40313 4091 40371 4097
rect 40405 4131 40463 4137
rect 40405 4097 40417 4131
rect 40451 4097 40463 4131
rect 40405 4091 40463 4097
rect 40533 4131 40591 4137
rect 40533 4097 40545 4131
rect 40579 4128 40591 4131
rect 40579 4100 40724 4128
rect 40579 4097 40591 4100
rect 40533 4091 40591 4097
rect 39853 4063 39911 4069
rect 39853 4060 39865 4063
rect 39592 4032 39865 4060
rect 39485 4023 39543 4029
rect 39853 4029 39865 4032
rect 39899 4029 39911 4063
rect 39853 4023 39911 4029
rect 36587 3964 38516 3992
rect 39500 3992 39528 4023
rect 39942 4020 39948 4072
rect 40000 4060 40006 4072
rect 40420 4060 40448 4091
rect 40696 4072 40724 4100
rect 40000 4032 40448 4060
rect 40000 4020 40006 4032
rect 40678 4020 40684 4072
rect 40736 4020 40742 4072
rect 41248 4060 41276 4159
rect 41506 4156 41512 4208
rect 41564 4196 41570 4208
rect 41564 4168 42196 4196
rect 41564 4156 41570 4168
rect 41414 4088 41420 4140
rect 41472 4088 41478 4140
rect 41856 4137 41884 4168
rect 41841 4131 41899 4137
rect 41841 4097 41853 4131
rect 41887 4097 41899 4131
rect 41841 4091 41899 4097
rect 41966 4088 41972 4140
rect 42024 4088 42030 4140
rect 42061 4131 42119 4137
rect 42061 4097 42073 4131
rect 42107 4097 42119 4131
rect 42168 4128 42196 4168
rect 42242 4156 42248 4208
rect 42300 4156 42306 4208
rect 43714 4196 43720 4208
rect 43180 4168 43720 4196
rect 43180 4128 43208 4168
rect 43714 4156 43720 4168
rect 43772 4156 43778 4208
rect 44361 4199 44419 4205
rect 44361 4165 44373 4199
rect 44407 4196 44419 4199
rect 45094 4196 45100 4208
rect 44407 4168 45100 4196
rect 44407 4165 44419 4168
rect 44361 4159 44419 4165
rect 45094 4156 45100 4168
rect 45152 4156 45158 4208
rect 45388 4205 45416 4236
rect 45646 4224 45652 4276
rect 45704 4224 45710 4276
rect 47026 4264 47032 4276
rect 46952 4236 47032 4264
rect 45373 4199 45431 4205
rect 45373 4165 45385 4199
rect 45419 4165 45431 4199
rect 45373 4159 45431 4165
rect 45462 4156 45468 4208
rect 45520 4156 45526 4208
rect 42168 4100 43208 4128
rect 43257 4131 43315 4137
rect 42061 4091 42119 4097
rect 43257 4097 43269 4131
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 44085 4131 44143 4137
rect 44085 4097 44097 4131
rect 44131 4128 44143 4131
rect 44131 4100 44312 4128
rect 45278 4127 45284 4140
rect 44131 4097 44143 4100
rect 44085 4091 44143 4097
rect 42076 4060 42104 4091
rect 41248 4032 42104 4060
rect 40129 3995 40187 4001
rect 40129 3992 40141 3995
rect 39500 3964 40141 3992
rect 36587 3961 36599 3964
rect 36541 3955 36599 3961
rect 40129 3961 40141 3964
rect 40175 3961 40187 3995
rect 41506 3992 41512 4004
rect 40129 3955 40187 3961
rect 40604 3964 41512 3992
rect 28552 3896 30604 3924
rect 30650 3884 30656 3936
rect 30708 3884 30714 3936
rect 30742 3884 30748 3936
rect 30800 3884 30806 3936
rect 31662 3884 31668 3936
rect 31720 3924 31726 3936
rect 32858 3924 32864 3936
rect 31720 3896 32864 3924
rect 31720 3884 31726 3896
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 35618 3884 35624 3936
rect 35676 3924 35682 3936
rect 36446 3924 36452 3936
rect 35676 3896 36452 3924
rect 35676 3884 35682 3896
rect 36446 3884 36452 3896
rect 36504 3884 36510 3936
rect 36814 3884 36820 3936
rect 36872 3884 36878 3936
rect 38746 3884 38752 3936
rect 38804 3884 38810 3936
rect 39574 3884 39580 3936
rect 39632 3884 39638 3936
rect 39945 3927 40003 3933
rect 39945 3893 39957 3927
rect 39991 3924 40003 3927
rect 40604 3924 40632 3964
rect 41506 3952 41512 3964
rect 41564 3952 41570 4004
rect 42076 3992 42104 4032
rect 42153 4063 42211 4069
rect 42153 4029 42165 4063
rect 42199 4060 42211 4063
rect 42429 4063 42487 4069
rect 42429 4060 42441 4063
rect 42199 4032 42441 4060
rect 42199 4029 42211 4032
rect 42153 4023 42211 4029
rect 42429 4029 42441 4032
rect 42475 4029 42487 4063
rect 42429 4023 42487 4029
rect 43070 4020 43076 4072
rect 43128 4020 43134 4072
rect 42978 3992 42984 4004
rect 42076 3964 42984 3992
rect 42978 3952 42984 3964
rect 43036 3952 43042 4004
rect 43272 3992 43300 4091
rect 44177 4063 44235 4069
rect 44177 4029 44189 4063
rect 44223 4029 44235 4063
rect 44284 4060 44312 4100
rect 45276 4088 45284 4127
rect 45336 4088 45342 4140
rect 45664 4137 45692 4224
rect 46290 4156 46296 4208
rect 46348 4196 46354 4208
rect 46348 4168 46612 4196
rect 46348 4156 46354 4168
rect 45649 4131 45707 4137
rect 45649 4097 45661 4131
rect 45695 4097 45707 4131
rect 45649 4091 45707 4097
rect 45738 4088 45744 4140
rect 45796 4088 45802 4140
rect 46584 4137 46612 4168
rect 46658 4156 46664 4208
rect 46716 4156 46722 4208
rect 46952 4205 46980 4236
rect 47026 4224 47032 4236
rect 47084 4224 47090 4276
rect 47228 4236 47440 4264
rect 47228 4205 47256 4236
rect 46937 4199 46995 4205
rect 46937 4165 46949 4199
rect 46983 4165 46995 4199
rect 47121 4199 47179 4205
rect 47121 4196 47133 4199
rect 46937 4159 46995 4165
rect 47025 4168 47133 4196
rect 45925 4131 45983 4137
rect 45925 4097 45937 4131
rect 45971 4128 45983 4131
rect 46017 4131 46075 4137
rect 46017 4128 46029 4131
rect 45971 4100 46029 4128
rect 45971 4097 45983 4100
rect 45925 4091 45983 4097
rect 46017 4097 46029 4100
rect 46063 4097 46075 4131
rect 46017 4091 46075 4097
rect 46569 4131 46627 4137
rect 46569 4097 46581 4131
rect 46615 4097 46627 4131
rect 46676 4128 46704 4156
rect 47025 4128 47053 4168
rect 47121 4165 47133 4168
rect 47167 4165 47179 4199
rect 47121 4159 47179 4165
rect 47213 4199 47271 4205
rect 47213 4165 47225 4199
rect 47259 4165 47271 4199
rect 47412 4196 47440 4236
rect 47762 4224 47768 4276
rect 47820 4264 47826 4276
rect 48593 4267 48651 4273
rect 47820 4236 48084 4264
rect 47820 4224 47826 4236
rect 47412 4168 47992 4196
rect 47213 4159 47271 4165
rect 46676 4100 47053 4128
rect 47325 4137 47383 4143
rect 47964 4140 47992 4168
rect 47325 4103 47337 4137
rect 47371 4134 47383 4137
rect 47371 4128 47440 4134
rect 47371 4106 47532 4128
rect 47371 4103 47383 4106
rect 47325 4097 47383 4103
rect 47412 4100 47532 4106
rect 46569 4091 46627 4097
rect 45276 4087 45288 4088
rect 45322 4087 45334 4088
rect 45276 4081 45334 4087
rect 47504 4072 47532 4100
rect 47946 4088 47952 4140
rect 48004 4088 48010 4140
rect 48056 4137 48084 4236
rect 48593 4233 48605 4267
rect 48639 4264 48651 4267
rect 48682 4264 48688 4276
rect 48639 4236 48688 4264
rect 48639 4233 48651 4236
rect 48593 4227 48651 4233
rect 48682 4224 48688 4236
rect 48740 4224 48746 4276
rect 49878 4224 49884 4276
rect 49936 4264 49942 4276
rect 50157 4267 50215 4273
rect 50157 4264 50169 4267
rect 49936 4236 50169 4264
rect 49936 4224 49942 4236
rect 50157 4233 50169 4236
rect 50203 4233 50215 4267
rect 50157 4227 50215 4233
rect 51000 4236 51120 4264
rect 51000 4208 51028 4236
rect 50982 4156 50988 4208
rect 51040 4156 51046 4208
rect 51092 4205 51120 4236
rect 53558 4224 53564 4276
rect 53616 4224 53622 4276
rect 53926 4264 53932 4276
rect 53668 4236 53932 4264
rect 51077 4199 51135 4205
rect 51077 4165 51089 4199
rect 51123 4165 51135 4199
rect 52917 4199 52975 4205
rect 52917 4196 52929 4199
rect 51077 4159 51135 4165
rect 52196 4168 52929 4196
rect 48041 4131 48099 4137
rect 48041 4097 48053 4131
rect 48087 4097 48099 4131
rect 48041 4091 48099 4097
rect 48225 4131 48283 4137
rect 48225 4097 48237 4131
rect 48271 4128 48283 4131
rect 49234 4128 49240 4140
rect 48271 4100 49240 4128
rect 48271 4097 48283 4100
rect 48225 4091 48283 4097
rect 49234 4088 49240 4100
rect 49292 4088 49298 4140
rect 49418 4088 49424 4140
rect 49476 4088 49482 4140
rect 49881 4131 49939 4137
rect 49881 4097 49893 4131
rect 49927 4128 49939 4131
rect 50430 4128 50436 4140
rect 49927 4100 50436 4128
rect 49927 4097 49939 4100
rect 49881 4091 49939 4097
rect 50430 4088 50436 4100
rect 50488 4088 50494 4140
rect 50706 4088 50712 4140
rect 50764 4128 50770 4140
rect 50893 4131 50951 4137
rect 50893 4128 50905 4131
rect 50764 4100 50905 4128
rect 50764 4088 50770 4100
rect 50893 4097 50905 4100
rect 50939 4097 50951 4131
rect 50893 4091 50951 4097
rect 51166 4088 51172 4140
rect 51224 4088 51230 4140
rect 51297 4131 51355 4137
rect 51297 4128 51309 4131
rect 51281 4097 51309 4128
rect 51343 4128 51355 4131
rect 51994 4128 52000 4140
rect 51343 4100 52000 4128
rect 51343 4097 51355 4100
rect 51281 4091 51355 4097
rect 44453 4063 44511 4069
rect 44453 4060 44465 4063
rect 44284 4032 44465 4060
rect 44177 4023 44235 4029
rect 44453 4029 44465 4032
rect 44499 4029 44511 4063
rect 44453 4023 44511 4029
rect 44082 3992 44088 4004
rect 43272 3964 44088 3992
rect 44082 3952 44088 3964
rect 44140 3952 44146 4004
rect 44192 3992 44220 4023
rect 44726 4020 44732 4072
rect 44784 4020 44790 4072
rect 45002 4020 45008 4072
rect 45060 4020 45066 4072
rect 47118 4020 47124 4072
rect 47176 4060 47182 4072
rect 47213 4063 47271 4069
rect 47213 4060 47225 4063
rect 47176 4032 47225 4060
rect 47176 4020 47182 4032
rect 47213 4029 47225 4032
rect 47259 4029 47271 4063
rect 47213 4023 47271 4029
rect 47486 4020 47492 4072
rect 47544 4020 47550 4072
rect 48958 4020 48964 4072
rect 49016 4060 49022 4072
rect 49605 4063 49663 4069
rect 49016 4032 49556 4060
rect 49016 4020 49022 4032
rect 44744 3992 44772 4020
rect 45649 3995 45707 4001
rect 45649 3992 45661 3995
rect 44192 3964 44404 3992
rect 44744 3964 45661 3992
rect 39991 3896 40632 3924
rect 39991 3893 40003 3896
rect 39945 3887 40003 3893
rect 40678 3884 40684 3936
rect 40736 3924 40742 3936
rect 40865 3927 40923 3933
rect 40865 3924 40877 3927
rect 40736 3896 40877 3924
rect 40736 3884 40742 3896
rect 40865 3893 40877 3896
rect 40911 3893 40923 3927
rect 40865 3887 40923 3893
rect 41601 3927 41659 3933
rect 41601 3893 41613 3927
rect 41647 3924 41659 3927
rect 41782 3924 41788 3936
rect 41647 3896 41788 3924
rect 41647 3893 41659 3896
rect 41601 3887 41659 3893
rect 41782 3884 41788 3896
rect 41840 3884 41846 3936
rect 43438 3884 43444 3936
rect 43496 3884 43502 3936
rect 43898 3884 43904 3936
rect 43956 3884 43962 3936
rect 44174 3884 44180 3936
rect 44232 3884 44238 3936
rect 44376 3924 44404 3964
rect 45649 3961 45661 3964
rect 45695 3961 45707 3995
rect 49237 3995 49295 4001
rect 49237 3992 49249 3995
rect 45649 3955 45707 3961
rect 45756 3964 49249 3992
rect 45756 3924 45784 3964
rect 49237 3961 49249 3964
rect 49283 3961 49295 3995
rect 49528 3992 49556 4032
rect 49605 4029 49617 4063
rect 49651 4060 49663 4063
rect 49786 4060 49792 4072
rect 49651 4032 49792 4060
rect 49651 4029 49663 4032
rect 49605 4023 49663 4029
rect 49786 4020 49792 4032
rect 49844 4020 49850 4072
rect 50801 4063 50859 4069
rect 50801 4029 50813 4063
rect 50847 4060 50859 4063
rect 50985 4063 51043 4069
rect 50985 4060 50997 4063
rect 50847 4032 50997 4060
rect 50847 4029 50859 4032
rect 50801 4023 50859 4029
rect 50985 4029 50997 4032
rect 51031 4029 51043 4063
rect 50985 4023 51043 4029
rect 51281 3992 51309 4091
rect 51994 4088 52000 4100
rect 52052 4128 52058 4140
rect 52196 4128 52224 4168
rect 52917 4165 52929 4168
rect 52963 4196 52975 4199
rect 53668 4196 53696 4236
rect 53926 4224 53932 4236
rect 53984 4224 53990 4276
rect 56318 4224 56324 4276
rect 56376 4224 56382 4276
rect 56594 4224 56600 4276
rect 56652 4264 56658 4276
rect 57146 4264 57152 4276
rect 56652 4236 56737 4264
rect 56652 4224 56658 4236
rect 52963 4168 53696 4196
rect 52963 4165 52975 4168
rect 52917 4159 52975 4165
rect 52052 4100 52224 4128
rect 52273 4131 52331 4137
rect 52052 4088 52058 4100
rect 52273 4097 52285 4131
rect 52319 4128 52331 4131
rect 52365 4131 52423 4137
rect 52365 4128 52377 4131
rect 52319 4100 52377 4128
rect 52319 4097 52331 4100
rect 52273 4091 52331 4097
rect 52365 4097 52377 4100
rect 52411 4097 52423 4131
rect 52365 4091 52423 4097
rect 52454 4088 52460 4140
rect 52512 4128 52518 4140
rect 52549 4131 52607 4137
rect 52549 4128 52561 4131
rect 52512 4100 52561 4128
rect 52512 4088 52518 4100
rect 52549 4097 52561 4100
rect 52595 4097 52607 4131
rect 52549 4091 52607 4097
rect 51629 4063 51687 4069
rect 51629 4029 51641 4063
rect 51675 4029 51687 4063
rect 52564 4060 52592 4091
rect 52822 4088 52828 4140
rect 52880 4128 52886 4140
rect 53193 4131 53251 4137
rect 53193 4128 53205 4131
rect 52880 4100 53205 4128
rect 52880 4088 52886 4100
rect 53193 4097 53205 4100
rect 53239 4097 53251 4131
rect 53193 4091 53251 4097
rect 53374 4088 53380 4140
rect 53432 4088 53438 4140
rect 54110 4088 54116 4140
rect 54168 4088 54174 4140
rect 54294 4088 54300 4140
rect 54352 4088 54358 4140
rect 54481 4131 54539 4137
rect 54481 4097 54493 4131
rect 54527 4097 54539 4131
rect 54481 4091 54539 4097
rect 54496 4060 54524 4091
rect 54570 4088 54576 4140
rect 54628 4128 54634 4140
rect 56336 4137 56364 4224
rect 56709 4159 56737 4236
rect 57072 4236 57152 4264
rect 57072 4205 57100 4236
rect 57146 4224 57152 4236
rect 57204 4224 57210 4276
rect 57057 4199 57115 4205
rect 57057 4165 57069 4199
rect 57103 4165 57115 4199
rect 57238 4196 57244 4208
rect 57057 4159 57115 4165
rect 57164 4168 57244 4196
rect 56709 4153 56767 4159
rect 54757 4131 54815 4137
rect 54757 4128 54769 4131
rect 54628 4100 54769 4128
rect 54628 4088 54634 4100
rect 54757 4097 54769 4100
rect 54803 4097 54815 4131
rect 54757 4091 54815 4097
rect 55217 4131 55275 4137
rect 55217 4097 55229 4131
rect 55263 4097 55275 4131
rect 55217 4091 55275 4097
rect 55401 4131 55459 4137
rect 55401 4097 55413 4131
rect 55447 4128 55459 4131
rect 55585 4131 55643 4137
rect 55585 4128 55597 4131
rect 55447 4100 55597 4128
rect 55447 4097 55459 4100
rect 55401 4091 55459 4097
rect 55585 4097 55597 4100
rect 55631 4097 55643 4131
rect 55585 4091 55643 4097
rect 56321 4131 56379 4137
rect 56321 4097 56333 4131
rect 56367 4097 56379 4131
rect 56321 4091 56379 4097
rect 56505 4131 56563 4137
rect 56505 4097 56517 4131
rect 56551 4097 56563 4131
rect 56505 4091 56563 4097
rect 56597 4131 56655 4137
rect 56597 4097 56609 4131
rect 56643 4097 56655 4131
rect 56709 4119 56721 4153
rect 56755 4119 56767 4153
rect 56962 4137 56968 4140
rect 56709 4113 56767 4119
rect 56597 4091 56655 4097
rect 56960 4091 56968 4137
rect 54846 4060 54852 4072
rect 52564 4032 54852 4060
rect 51629 4023 51687 4029
rect 49528 3964 51309 3992
rect 49237 3955 49295 3961
rect 51350 3952 51356 4004
rect 51408 3992 51414 4004
rect 51644 3992 51672 4023
rect 54846 4020 54852 4032
rect 54904 4060 54910 4072
rect 55033 4063 55091 4069
rect 55033 4060 55045 4063
rect 54904 4032 55045 4060
rect 54904 4020 54910 4032
rect 55033 4029 55045 4032
rect 55079 4060 55091 4063
rect 55232 4060 55260 4091
rect 55079 4032 55260 4060
rect 56229 4063 56287 4069
rect 55079 4029 55091 4032
rect 55033 4023 55091 4029
rect 56229 4029 56241 4063
rect 56275 4060 56287 4063
rect 56413 4063 56471 4069
rect 56413 4060 56425 4063
rect 56275 4032 56425 4060
rect 56275 4029 56287 4032
rect 56229 4023 56287 4029
rect 56413 4029 56425 4032
rect 56459 4029 56471 4063
rect 56413 4023 56471 4029
rect 51408 3964 51672 3992
rect 56520 3992 56548 4091
rect 56612 4060 56640 4091
rect 56962 4088 56968 4091
rect 57020 4088 57026 4140
rect 57164 4137 57192 4168
rect 57238 4156 57244 4168
rect 57296 4156 57302 4208
rect 57330 4156 57336 4208
rect 57388 4156 57394 4208
rect 57149 4131 57207 4137
rect 57149 4097 57161 4131
rect 57195 4097 57207 4131
rect 57149 4091 57207 4097
rect 56870 4060 56876 4072
rect 56612 4032 56876 4060
rect 56870 4020 56876 4032
rect 56928 4020 56934 4072
rect 57164 3992 57192 4091
rect 57422 4088 57428 4140
rect 57480 4088 57486 4140
rect 57241 4063 57299 4069
rect 57241 4029 57253 4063
rect 57287 4060 57299 4063
rect 57885 4063 57943 4069
rect 57885 4060 57897 4063
rect 57287 4032 57897 4060
rect 57287 4029 57299 4032
rect 57241 4023 57299 4029
rect 57885 4029 57897 4032
rect 57931 4029 57943 4063
rect 57885 4023 57943 4029
rect 56520 3964 57192 3992
rect 51408 3952 51414 3964
rect 44376 3896 45784 3924
rect 45830 3884 45836 3936
rect 45888 3924 45894 3936
rect 45925 3927 45983 3933
rect 45925 3924 45937 3927
rect 45888 3896 45937 3924
rect 45888 3884 45894 3896
rect 45925 3893 45937 3896
rect 45971 3893 45983 3927
rect 45925 3887 45983 3893
rect 46474 3884 46480 3936
rect 46532 3924 46538 3936
rect 47762 3924 47768 3936
rect 46532 3896 47768 3924
rect 46532 3884 46538 3896
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 48038 3884 48044 3936
rect 48096 3924 48102 3936
rect 48225 3927 48283 3933
rect 48225 3924 48237 3927
rect 48096 3896 48237 3924
rect 48096 3884 48102 3896
rect 48225 3893 48237 3896
rect 48271 3893 48283 3927
rect 48225 3887 48283 3893
rect 49605 3927 49663 3933
rect 49605 3893 49617 3927
rect 49651 3924 49663 3927
rect 50246 3924 50252 3936
rect 49651 3896 50252 3924
rect 49651 3893 49663 3896
rect 49605 3887 49663 3893
rect 50246 3884 50252 3896
rect 50304 3884 50310 3936
rect 52362 3884 52368 3936
rect 52420 3884 52426 3936
rect 54294 3884 54300 3936
rect 54352 3884 54358 3936
rect 54570 3884 54576 3936
rect 54628 3884 54634 3936
rect 55398 3884 55404 3936
rect 55456 3884 55462 3936
rect 57606 3884 57612 3936
rect 57664 3884 57670 3936
rect 58529 3927 58587 3933
rect 58529 3893 58541 3927
rect 58575 3924 58587 3927
rect 58575 3896 58940 3924
rect 58575 3893 58587 3896
rect 58529 3887 58587 3893
rect 1104 3834 58880 3856
rect 1104 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 22616 3834
rect 22668 3782 22680 3834
rect 22732 3782 22744 3834
rect 22796 3782 22808 3834
rect 22860 3782 22872 3834
rect 22924 3782 37060 3834
rect 37112 3782 37124 3834
rect 37176 3782 37188 3834
rect 37240 3782 37252 3834
rect 37304 3782 37316 3834
rect 37368 3782 51504 3834
rect 51556 3782 51568 3834
rect 51620 3782 51632 3834
rect 51684 3782 51696 3834
rect 51748 3782 51760 3834
rect 51812 3782 58880 3834
rect 1104 3760 58880 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3016 3692 3157 3720
rect 3016 3680 3022 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 6178 3680 6184 3732
rect 6236 3680 6242 3732
rect 6270 3680 6276 3732
rect 6328 3680 6334 3732
rect 6638 3680 6644 3732
rect 6696 3680 6702 3732
rect 10505 3723 10563 3729
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 11054 3720 11060 3732
rect 10551 3692 11060 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 13446 3720 13452 3732
rect 11164 3692 13452 3720
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 11164 3652 11192 3692
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13596 3692 13921 3720
rect 13596 3680 13602 3692
rect 13909 3689 13921 3692
rect 13955 3689 13967 3723
rect 13909 3683 13967 3689
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 16482 3720 16488 3732
rect 14424 3692 16488 3720
rect 14424 3680 14430 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 17586 3680 17592 3732
rect 17644 3680 17650 3732
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18690 3720 18696 3732
rect 18104 3692 18696 3720
rect 18104 3680 18110 3692
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 19058 3680 19064 3732
rect 19116 3680 19122 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20864 3692 20913 3720
rect 20864 3680 20870 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 22465 3723 22523 3729
rect 22465 3689 22477 3723
rect 22511 3689 22523 3723
rect 22465 3683 22523 3689
rect 22741 3723 22799 3729
rect 22741 3689 22753 3723
rect 22787 3720 22799 3723
rect 24118 3720 24124 3732
rect 22787 3692 24124 3720
rect 22787 3689 22799 3692
rect 22741 3683 22799 3689
rect 10008 3624 11192 3652
rect 14185 3655 14243 3661
rect 10008 3612 10014 3624
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3050 3584 3056 3596
rect 3007 3556 3056 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3050 3544 3056 3556
rect 3108 3584 3114 3596
rect 4062 3584 4068 3596
rect 3108 3556 4068 3584
rect 3108 3544 3114 3556
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 4120 3556 4844 3584
rect 4120 3544 4126 3556
rect 3326 3476 3332 3528
rect 3384 3476 3390 3528
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 3605 3519 3663 3525
rect 3605 3516 3617 3519
rect 3568 3488 3617 3516
rect 3568 3476 3574 3488
rect 3605 3485 3617 3488
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3752 3488 4353 3516
rect 3752 3476 3758 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4816 3525 4844 3556
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6420 3556 6500 3584
rect 6420 3544 6426 3556
rect 6472 3525 6500 3556
rect 7852 3556 8984 3584
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 6457 3519 6515 3525
rect 4847 3488 6408 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 2716 3451 2774 3457
rect 1820 3420 2268 3448
rect 1820 3408 1826 3420
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 2130 3380 2136 3392
rect 1627 3352 2136 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 2240 3380 2268 3420
rect 2716 3417 2728 3451
rect 2762 3448 2774 3451
rect 3789 3451 3847 3457
rect 3789 3448 3801 3451
rect 2762 3420 3801 3448
rect 2762 3417 2774 3420
rect 2716 3411 2774 3417
rect 3789 3417 3801 3420
rect 3835 3417 3847 3451
rect 3789 3411 3847 3417
rect 3970 3408 3976 3460
rect 4028 3408 4034 3460
rect 5068 3451 5126 3457
rect 5068 3417 5080 3451
rect 5114 3448 5126 3451
rect 5350 3448 5356 3460
rect 5114 3420 5356 3448
rect 5114 3417 5126 3420
rect 5068 3411 5126 3417
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 6380 3448 6408 3488
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7852 3516 7880 3556
rect 6871 3488 7880 3516
rect 8297 3519 8355 3525
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 8846 3516 8852 3528
rect 8343 3488 8852 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 6840 3448 6868 3479
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 8956 3525 8984 3556
rect 10893 3535 10921 3624
rect 14185 3621 14197 3655
rect 14231 3652 14243 3655
rect 14826 3652 14832 3664
rect 14231 3624 14832 3652
rect 14231 3621 14243 3624
rect 14185 3615 14243 3621
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 15013 3655 15071 3661
rect 15013 3621 15025 3655
rect 15059 3652 15071 3655
rect 15286 3652 15292 3664
rect 15059 3624 15292 3652
rect 15059 3621 15071 3624
rect 15013 3615 15071 3621
rect 15286 3612 15292 3624
rect 15344 3612 15350 3664
rect 22480 3596 22508 3683
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25498 3720 25504 3732
rect 25188 3692 25504 3720
rect 25188 3680 25194 3692
rect 25498 3680 25504 3692
rect 25556 3720 25562 3732
rect 25869 3723 25927 3729
rect 25869 3720 25881 3723
rect 25556 3692 25881 3720
rect 25556 3680 25562 3692
rect 25869 3689 25881 3692
rect 25915 3689 25927 3723
rect 28810 3720 28816 3732
rect 25869 3683 25927 3689
rect 27816 3692 28816 3720
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14553 3587 14611 3593
rect 14332 3556 14504 3584
rect 14332 3544 14338 3556
rect 10878 3529 10936 3535
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 10042 3516 10048 3528
rect 8987 3488 10048 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10878 3495 10890 3529
rect 10924 3495 10936 3529
rect 10878 3489 10936 3495
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12526 3516 12532 3528
rect 12483 3488 12532 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12526 3476 12532 3488
rect 12584 3516 12590 3528
rect 12584 3488 14320 3516
rect 12584 3476 12590 3488
rect 6380 3420 6868 3448
rect 7092 3451 7150 3457
rect 7092 3417 7104 3451
rect 7138 3448 7150 3451
rect 7558 3448 7564 3460
rect 7138 3420 7564 3448
rect 7138 3417 7150 3420
rect 7092 3411 7150 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 8573 3451 8631 3457
rect 8573 3417 8585 3451
rect 8619 3448 8631 3451
rect 8754 3448 8760 3460
rect 8619 3420 8760 3448
rect 8619 3417 8631 3420
rect 8573 3411 8631 3417
rect 8754 3408 8760 3420
rect 8812 3448 8818 3460
rect 9208 3451 9266 3457
rect 8812 3420 9168 3448
rect 8812 3408 8818 3420
rect 3513 3383 3571 3389
rect 3513 3380 3525 3383
rect 2240 3352 3525 3380
rect 3513 3349 3525 3352
rect 3559 3380 3571 3383
rect 3988 3380 4016 3408
rect 3559 3352 4016 3380
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 4706 3340 4712 3392
rect 4764 3340 4770 3392
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8662 3380 8668 3392
rect 8251 3352 8668 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9140 3380 9168 3420
rect 9208 3417 9220 3451
rect 9254 3448 9266 3451
rect 9490 3448 9496 3460
rect 9254 3420 9496 3448
rect 9254 3417 9266 3420
rect 9208 3411 9266 3417
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 10502 3408 10508 3460
rect 10560 3408 10566 3460
rect 10594 3408 10600 3460
rect 10652 3448 10658 3460
rect 10689 3451 10747 3457
rect 10689 3448 10701 3451
rect 10652 3420 10701 3448
rect 10652 3408 10658 3420
rect 10689 3417 10701 3420
rect 10735 3417 10747 3451
rect 10689 3411 10747 3417
rect 10781 3451 10839 3457
rect 10781 3417 10793 3451
rect 10827 3417 10839 3451
rect 10781 3411 10839 3417
rect 12170 3451 12228 3457
rect 12170 3417 12182 3451
rect 12216 3417 12228 3451
rect 12170 3411 12228 3417
rect 12796 3451 12854 3457
rect 12796 3417 12808 3451
rect 12842 3448 12854 3451
rect 13354 3448 13360 3460
rect 12842 3420 13360 3448
rect 12842 3417 12854 3420
rect 12796 3411 12854 3417
rect 9398 3380 9404 3392
rect 9140 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 10284 3352 10333 3380
rect 10284 3340 10290 3352
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 10796 3380 10824 3411
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10796 3352 11069 3380
rect 10321 3343 10379 3349
rect 11057 3349 11069 3352
rect 11103 3380 11115 3383
rect 12066 3380 12072 3392
rect 11103 3352 12072 3380
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12176 3380 12204 3411
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 14292 3448 14320 3488
rect 14366 3476 14372 3528
rect 14424 3476 14430 3528
rect 14476 3525 14504 3556
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 14599 3556 15424 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 14467 3519 14525 3525
rect 14467 3485 14479 3519
rect 14513 3485 14525 3519
rect 14467 3479 14525 3485
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3516 14703 3519
rect 14734 3516 14740 3528
rect 14691 3488 14740 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15396 3516 15424 3556
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 17460 3556 17693 3584
rect 17460 3544 17466 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 21085 3587 21143 3593
rect 21085 3584 21097 3587
rect 17681 3547 17739 3553
rect 20640 3556 21097 3584
rect 15545 3519 15603 3525
rect 15545 3516 15557 3519
rect 15396 3488 15557 3516
rect 15289 3479 15347 3485
rect 15545 3485 15557 3488
rect 15591 3485 15603 3519
rect 15545 3479 15603 3485
rect 14550 3448 14556 3460
rect 14292 3420 14556 3448
rect 14550 3408 14556 3420
rect 14608 3448 14614 3460
rect 15304 3448 15332 3479
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 17696 3516 17724 3547
rect 20640 3525 20668 3556
rect 21085 3553 21097 3556
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 20358 3519 20416 3525
rect 17696 3488 20300 3516
rect 14608 3420 15332 3448
rect 17948 3451 18006 3457
rect 14608 3408 14614 3420
rect 17948 3417 17960 3451
rect 17994 3448 18006 3451
rect 18598 3448 18604 3460
rect 17994 3420 18604 3448
rect 17994 3417 18006 3420
rect 17948 3411 18006 3417
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 12250 3380 12256 3392
rect 12176 3352 12256 3380
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 15194 3340 15200 3392
rect 15252 3380 15258 3392
rect 15930 3380 15936 3392
rect 15252 3352 15936 3380
rect 15252 3340 15258 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 17586 3380 17592 3392
rect 16724 3352 17592 3380
rect 16724 3340 16730 3352
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 19245 3383 19303 3389
rect 19245 3349 19257 3383
rect 19291 3380 19303 3383
rect 19978 3380 19984 3392
rect 19291 3352 19984 3380
rect 19291 3349 19303 3352
rect 19245 3343 19303 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20272 3380 20300 3488
rect 20358 3485 20370 3519
rect 20404 3485 20416 3519
rect 20358 3479 20416 3485
rect 20625 3519 20683 3525
rect 20625 3485 20637 3519
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 20364 3448 20392 3479
rect 20438 3448 20444 3460
rect 20364 3420 20444 3448
rect 20438 3408 20444 3420
rect 20496 3408 20502 3460
rect 20640 3380 20668 3479
rect 20714 3476 20720 3528
rect 20772 3476 20778 3528
rect 21100 3516 21128 3547
rect 22462 3544 22468 3596
rect 22520 3544 22526 3596
rect 22278 3516 22284 3528
rect 21100 3488 22284 3516
rect 22278 3476 22284 3488
rect 22336 3516 22342 3528
rect 22557 3519 22615 3525
rect 22336 3488 22508 3516
rect 22336 3476 22342 3488
rect 21358 3457 21364 3460
rect 21352 3448 21364 3457
rect 21319 3420 21364 3448
rect 21352 3411 21364 3420
rect 21358 3408 21364 3411
rect 21416 3408 21422 3460
rect 21634 3408 21640 3460
rect 21692 3448 21698 3460
rect 22480 3448 22508 3488
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 22738 3516 22744 3528
rect 22603 3488 22744 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 24489 3519 24547 3525
rect 24489 3516 24501 3519
rect 22879 3488 24501 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 24489 3485 24501 3488
rect 24535 3516 24547 3519
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 24535 3488 25973 3516
rect 24535 3485 24547 3488
rect 24489 3479 24547 3485
rect 25961 3485 25973 3488
rect 26007 3516 26019 3519
rect 27617 3519 27675 3525
rect 26007 3488 26372 3516
rect 26007 3485 26019 3488
rect 25961 3479 26019 3485
rect 22848 3448 22876 3479
rect 23078 3451 23136 3457
rect 23078 3448 23090 3451
rect 21692 3420 22094 3448
rect 22480 3420 22876 3448
rect 22940 3420 23090 3448
rect 21692 3408 21698 3420
rect 20272 3352 20668 3380
rect 22066 3380 22094 3420
rect 22940 3380 22968 3420
rect 23078 3417 23090 3420
rect 23124 3417 23136 3451
rect 23078 3411 23136 3417
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 26234 3457 26240 3460
rect 24734 3451 24792 3457
rect 24734 3448 24746 3451
rect 24176 3420 24746 3448
rect 24176 3408 24182 3420
rect 24734 3417 24746 3420
rect 24780 3417 24792 3451
rect 26228 3448 26240 3457
rect 26195 3420 26240 3448
rect 24734 3411 24792 3417
rect 26228 3411 26240 3420
rect 26234 3408 26240 3411
rect 26292 3408 26298 3460
rect 26344 3448 26372 3488
rect 27617 3485 27629 3519
rect 27663 3516 27675 3519
rect 27706 3516 27712 3528
rect 27663 3488 27712 3516
rect 27663 3485 27675 3488
rect 27617 3479 27675 3485
rect 27706 3476 27712 3488
rect 27764 3476 27770 3528
rect 27816 3525 27844 3692
rect 28810 3680 28816 3692
rect 28868 3680 28874 3732
rect 30742 3680 30748 3732
rect 30800 3680 30806 3732
rect 30929 3723 30987 3729
rect 30929 3720 30941 3723
rect 30852 3692 30941 3720
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3485 27859 3519
rect 27801 3479 27859 3485
rect 27893 3519 27951 3525
rect 27893 3485 27905 3519
rect 27939 3516 27951 3519
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 27939 3488 29561 3516
rect 27939 3485 27951 3488
rect 27893 3479 27951 3485
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 29816 3519 29874 3525
rect 29816 3485 29828 3519
rect 29862 3516 29874 3519
rect 30760 3516 30788 3680
rect 29862 3488 30788 3516
rect 29862 3485 29874 3488
rect 29816 3479 29874 3485
rect 27908 3448 27936 3479
rect 30852 3460 30880 3692
rect 30929 3689 30941 3692
rect 30975 3689 30987 3723
rect 31662 3720 31668 3732
rect 30929 3683 30987 3689
rect 31220 3692 31668 3720
rect 31220 3525 31248 3692
rect 31662 3680 31668 3692
rect 31720 3680 31726 3732
rect 33502 3720 33508 3732
rect 33152 3692 33508 3720
rect 31478 3544 31484 3596
rect 31536 3544 31542 3596
rect 33152 3593 33180 3692
rect 33502 3680 33508 3692
rect 33560 3720 33566 3732
rect 37645 3723 37703 3729
rect 33560 3692 36308 3720
rect 33560 3680 33566 3692
rect 34517 3655 34575 3661
rect 34517 3621 34529 3655
rect 34563 3621 34575 3655
rect 34517 3615 34575 3621
rect 33137 3587 33195 3593
rect 33137 3553 33149 3587
rect 33183 3553 33195 3587
rect 33137 3547 33195 3553
rect 31205 3519 31263 3525
rect 31205 3485 31217 3519
rect 31251 3485 31263 3519
rect 31205 3479 31263 3485
rect 31386 3476 31392 3528
rect 31444 3476 31450 3528
rect 34532 3516 34560 3615
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 34664 3624 36216 3652
rect 34664 3612 34670 3624
rect 34793 3587 34851 3593
rect 34793 3553 34805 3587
rect 34839 3584 34851 3587
rect 35437 3587 35495 3593
rect 35437 3584 35449 3587
rect 34839 3556 35449 3584
rect 34839 3553 34851 3556
rect 34793 3547 34851 3553
rect 35437 3553 35449 3556
rect 35483 3553 35495 3587
rect 35437 3547 35495 3553
rect 35802 3516 35808 3528
rect 35860 3525 35866 3528
rect 36188 3525 36216 3624
rect 36280 3593 36308 3692
rect 37645 3689 37657 3723
rect 37691 3720 37703 3723
rect 38194 3720 38200 3732
rect 37691 3692 38200 3720
rect 37691 3689 37703 3692
rect 37645 3683 37703 3689
rect 38194 3680 38200 3692
rect 38252 3680 38258 3732
rect 38562 3680 38568 3732
rect 38620 3720 38626 3732
rect 39758 3720 39764 3732
rect 38620 3692 39764 3720
rect 38620 3680 38626 3692
rect 39758 3680 39764 3692
rect 39816 3680 39822 3732
rect 40034 3720 40040 3732
rect 39868 3692 40040 3720
rect 39301 3655 39359 3661
rect 39301 3621 39313 3655
rect 39347 3652 39359 3655
rect 39868 3652 39896 3692
rect 40034 3680 40040 3692
rect 40092 3680 40098 3732
rect 43349 3723 43407 3729
rect 43349 3689 43361 3723
rect 43395 3720 43407 3723
rect 43395 3692 44404 3720
rect 43395 3689 43407 3692
rect 43349 3683 43407 3689
rect 39347 3624 39896 3652
rect 44376 3652 44404 3692
rect 44818 3680 44824 3732
rect 44876 3680 44882 3732
rect 45922 3720 45928 3732
rect 45296 3692 45928 3720
rect 45005 3655 45063 3661
rect 45005 3652 45017 3655
rect 44376 3624 45017 3652
rect 39347 3621 39359 3624
rect 39301 3615 39359 3621
rect 45005 3621 45017 3624
rect 45051 3621 45063 3655
rect 45005 3615 45063 3621
rect 36265 3587 36323 3593
rect 36265 3553 36277 3587
rect 36311 3553 36323 3587
rect 36265 3547 36323 3553
rect 39592 3556 39896 3584
rect 34532 3488 35572 3516
rect 35768 3488 35808 3516
rect 28138 3451 28196 3457
rect 28138 3448 28150 3451
rect 26344 3420 27936 3448
rect 28000 3420 28150 3448
rect 22066 3352 22968 3380
rect 24210 3340 24216 3392
rect 24268 3340 24274 3392
rect 27338 3340 27344 3392
rect 27396 3340 27402 3392
rect 27709 3383 27767 3389
rect 27709 3349 27721 3383
rect 27755 3380 27767 3383
rect 28000 3380 28028 3420
rect 28138 3417 28150 3420
rect 28184 3417 28196 3451
rect 28138 3411 28196 3417
rect 28442 3408 28448 3460
rect 28500 3408 28506 3460
rect 30374 3408 30380 3460
rect 30432 3448 30438 3460
rect 30834 3448 30840 3460
rect 30432 3420 30840 3448
rect 30432 3408 30438 3420
rect 30834 3408 30840 3420
rect 30892 3408 30898 3460
rect 31297 3451 31355 3457
rect 31297 3417 31309 3451
rect 31343 3448 31355 3451
rect 31726 3451 31784 3457
rect 31726 3448 31738 3451
rect 31343 3420 31738 3448
rect 31343 3417 31355 3420
rect 31297 3411 31355 3417
rect 31726 3417 31738 3420
rect 31772 3417 31784 3451
rect 31726 3411 31784 3417
rect 33404 3451 33462 3457
rect 33404 3417 33416 3451
rect 33450 3448 33462 3451
rect 34882 3448 34888 3460
rect 33450 3420 34888 3448
rect 33450 3417 33462 3420
rect 33404 3411 33462 3417
rect 34882 3408 34888 3420
rect 34940 3408 34946 3460
rect 35158 3408 35164 3460
rect 35216 3448 35222 3460
rect 35437 3451 35495 3457
rect 35437 3448 35449 3451
rect 35216 3420 35449 3448
rect 35216 3408 35222 3420
rect 35437 3417 35449 3420
rect 35483 3417 35495 3451
rect 35437 3411 35495 3417
rect 27755 3352 28028 3380
rect 28460 3380 28488 3408
rect 29270 3380 29276 3392
rect 28460 3352 29276 3380
rect 27755 3349 27767 3352
rect 27709 3343 27767 3349
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 32861 3383 32919 3389
rect 32861 3349 32873 3383
rect 32907 3380 32919 3383
rect 33686 3380 33692 3392
rect 32907 3352 33692 3380
rect 32907 3349 32919 3352
rect 32861 3343 32919 3349
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 35342 3340 35348 3392
rect 35400 3340 35406 3392
rect 35544 3380 35572 3488
rect 35802 3476 35808 3488
rect 35860 3479 35868 3525
rect 36173 3519 36231 3525
rect 36173 3485 36185 3519
rect 36219 3485 36231 3519
rect 36280 3516 36308 3547
rect 37458 3516 37464 3528
rect 36280 3488 37464 3516
rect 36173 3479 36231 3485
rect 35860 3476 35866 3479
rect 37458 3476 37464 3488
rect 37516 3516 37522 3528
rect 37921 3519 37979 3525
rect 37921 3516 37933 3519
rect 37516 3488 37933 3516
rect 37516 3476 37522 3488
rect 37921 3485 37933 3488
rect 37967 3516 37979 3519
rect 39592 3516 39620 3556
rect 39868 3525 39896 3556
rect 40862 3544 40868 3596
rect 40920 3544 40926 3596
rect 45296 3593 45324 3692
rect 45922 3680 45928 3692
rect 45980 3720 45986 3732
rect 50154 3720 50160 3732
rect 45980 3692 50160 3720
rect 45980 3680 45986 3692
rect 46934 3612 46940 3664
rect 46992 3612 46998 3664
rect 47780 3593 47808 3692
rect 50154 3680 50160 3692
rect 50212 3680 50218 3732
rect 53834 3680 53840 3732
rect 53892 3720 53898 3732
rect 54573 3723 54631 3729
rect 54573 3720 54585 3723
rect 53892 3692 54585 3720
rect 53892 3680 53898 3692
rect 54573 3689 54585 3692
rect 54619 3689 54631 3723
rect 54573 3683 54631 3689
rect 55033 3723 55091 3729
rect 55033 3689 55045 3723
rect 55079 3720 55091 3723
rect 56594 3720 56600 3732
rect 55079 3692 56600 3720
rect 55079 3689 55091 3692
rect 55033 3683 55091 3689
rect 56594 3680 56600 3692
rect 56652 3680 56658 3732
rect 56873 3723 56931 3729
rect 56873 3689 56885 3723
rect 56919 3720 56931 3723
rect 57146 3720 57152 3732
rect 56919 3692 57152 3720
rect 56919 3689 56931 3692
rect 56873 3683 56931 3689
rect 57146 3680 57152 3692
rect 57204 3680 57210 3732
rect 58250 3680 58256 3732
rect 58308 3720 58314 3732
rect 58529 3723 58587 3729
rect 58529 3720 58541 3723
rect 58308 3692 58541 3720
rect 58308 3680 58314 3692
rect 58529 3689 58541 3692
rect 58575 3689 58587 3723
rect 58529 3683 58587 3689
rect 49234 3612 49240 3664
rect 49292 3612 49298 3664
rect 50172 3593 50200 3680
rect 43441 3587 43499 3593
rect 43441 3584 43453 3587
rect 42720 3556 43453 3584
rect 37967 3488 39620 3516
rect 39669 3519 39727 3525
rect 37967 3485 37979 3488
rect 37921 3479 37979 3485
rect 39669 3485 39681 3519
rect 39715 3485 39727 3519
rect 39669 3479 39727 3485
rect 39853 3519 39911 3525
rect 39853 3485 39865 3519
rect 39899 3516 39911 3519
rect 40880 3516 40908 3544
rect 42720 3525 42748 3556
rect 43441 3553 43453 3556
rect 43487 3553 43499 3587
rect 43441 3547 43499 3553
rect 45281 3587 45339 3593
rect 45281 3553 45293 3587
rect 45327 3553 45339 3587
rect 45281 3547 45339 3553
rect 47765 3587 47823 3593
rect 47765 3553 47777 3587
rect 47811 3553 47823 3587
rect 47765 3547 47823 3553
rect 50157 3587 50215 3593
rect 50157 3553 50169 3587
rect 50203 3553 50215 3587
rect 50157 3547 50215 3553
rect 54481 3587 54539 3593
rect 54481 3553 54493 3587
rect 54527 3584 54539 3587
rect 54527 3556 55352 3584
rect 54527 3553 54539 3556
rect 54481 3547 54539 3553
rect 42705 3519 42763 3525
rect 42705 3516 42717 3519
rect 39899 3488 42717 3516
rect 39899 3485 39911 3488
rect 39853 3479 39911 3485
rect 42705 3485 42717 3488
rect 42751 3485 42763 3519
rect 42705 3479 42763 3485
rect 43073 3519 43131 3525
rect 43073 3485 43085 3519
rect 43119 3485 43131 3519
rect 43073 3479 43131 3485
rect 35618 3408 35624 3460
rect 35676 3408 35682 3460
rect 35713 3451 35771 3457
rect 35713 3417 35725 3451
rect 35759 3417 35771 3451
rect 35713 3411 35771 3417
rect 36532 3451 36590 3457
rect 36532 3417 36544 3451
rect 36578 3448 36590 3451
rect 36814 3448 36820 3460
rect 36578 3420 36820 3448
rect 36578 3417 36590 3420
rect 36532 3411 36590 3417
rect 35728 3380 35756 3411
rect 36814 3408 36820 3420
rect 36872 3408 36878 3460
rect 38188 3451 38246 3457
rect 38188 3417 38200 3451
rect 38234 3448 38246 3451
rect 38746 3448 38752 3460
rect 38234 3420 38752 3448
rect 38234 3417 38246 3420
rect 38188 3411 38246 3417
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 35894 3380 35900 3392
rect 35544 3352 35900 3380
rect 35894 3340 35900 3352
rect 35952 3340 35958 3392
rect 35989 3383 36047 3389
rect 35989 3349 36001 3383
rect 36035 3380 36047 3383
rect 36170 3380 36176 3392
rect 36035 3352 36176 3380
rect 36035 3349 36047 3352
rect 35989 3343 36047 3349
rect 36170 3340 36176 3352
rect 36228 3340 36234 3392
rect 38102 3340 38108 3392
rect 38160 3380 38166 3392
rect 39390 3380 39396 3392
rect 38160 3352 39396 3380
rect 38160 3340 38166 3352
rect 39390 3340 39396 3352
rect 39448 3340 39454 3392
rect 39482 3340 39488 3392
rect 39540 3340 39546 3392
rect 39684 3380 39712 3479
rect 40126 3457 40132 3460
rect 40120 3411 40132 3457
rect 40126 3408 40132 3411
rect 40184 3408 40190 3460
rect 42460 3451 42518 3457
rect 42460 3417 42472 3451
rect 42506 3448 42518 3451
rect 42610 3448 42616 3460
rect 42506 3420 42616 3448
rect 42506 3417 42518 3420
rect 42460 3411 42518 3417
rect 42610 3408 42616 3420
rect 42668 3408 42674 3460
rect 43088 3448 43116 3479
rect 43162 3476 43168 3528
rect 43220 3476 43226 3528
rect 43530 3476 43536 3528
rect 43588 3516 43594 3528
rect 43697 3519 43755 3525
rect 43697 3516 43709 3519
rect 43588 3488 43709 3516
rect 43588 3476 43594 3488
rect 43697 3485 43709 3488
rect 43743 3485 43755 3519
rect 43697 3479 43755 3485
rect 44634 3476 44640 3528
rect 44692 3516 44698 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44692 3488 45201 3516
rect 44692 3476 44698 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45548 3519 45606 3525
rect 45548 3485 45560 3519
rect 45594 3516 45606 3519
rect 45830 3516 45836 3528
rect 45594 3488 45836 3516
rect 45594 3485 45606 3488
rect 45548 3479 45606 3485
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 47118 3476 47124 3528
rect 47176 3476 47182 3528
rect 48038 3525 48044 3528
rect 48032 3516 48044 3525
rect 47999 3488 48044 3516
rect 48032 3479 48044 3488
rect 48038 3476 48044 3479
rect 48096 3476 48102 3528
rect 49050 3476 49056 3528
rect 49108 3516 49114 3528
rect 49789 3519 49847 3525
rect 49789 3516 49801 3519
rect 49108 3488 49801 3516
rect 49108 3476 49114 3488
rect 49789 3485 49801 3488
rect 49835 3485 49847 3519
rect 49789 3479 49847 3485
rect 50062 3476 50068 3528
rect 50120 3516 50126 3528
rect 50413 3519 50471 3525
rect 50413 3516 50425 3519
rect 50120 3488 50425 3516
rect 50120 3476 50126 3488
rect 50413 3485 50425 3488
rect 50459 3485 50471 3519
rect 50413 3479 50471 3485
rect 52362 3476 52368 3528
rect 52420 3516 52426 3528
rect 52742 3519 52800 3525
rect 52742 3516 52754 3519
rect 52420 3488 52754 3516
rect 52420 3476 52426 3488
rect 52742 3485 52754 3488
rect 52788 3485 52800 3519
rect 52742 3479 52800 3485
rect 53006 3476 53012 3528
rect 53064 3516 53070 3528
rect 54214 3519 54272 3525
rect 53064 3488 54064 3516
rect 53064 3476 53070 3488
rect 42720 3420 43116 3448
rect 42720 3392 42748 3420
rect 43346 3408 43352 3460
rect 43404 3408 43410 3460
rect 46198 3408 46204 3460
rect 46256 3448 46262 3460
rect 47397 3451 47455 3457
rect 47397 3448 47409 3451
rect 46256 3420 47409 3448
rect 46256 3408 46262 3420
rect 47397 3417 47409 3420
rect 47443 3448 47455 3451
rect 47486 3448 47492 3460
rect 47443 3420 47492 3448
rect 47443 3417 47455 3420
rect 47397 3411 47455 3417
rect 47486 3408 47492 3420
rect 47544 3448 47550 3460
rect 48958 3448 48964 3460
rect 47544 3420 48964 3448
rect 47544 3408 47550 3420
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 51166 3408 51172 3460
rect 51224 3448 51230 3460
rect 52178 3448 52184 3460
rect 51224 3420 52184 3448
rect 51224 3408 51230 3420
rect 40494 3380 40500 3392
rect 39684 3352 40500 3380
rect 40494 3340 40500 3352
rect 40552 3340 40558 3392
rect 41230 3340 41236 3392
rect 41288 3340 41294 3392
rect 41325 3383 41383 3389
rect 41325 3349 41337 3383
rect 41371 3380 41383 3383
rect 41966 3380 41972 3392
rect 41371 3352 41972 3380
rect 41371 3349 41383 3352
rect 41325 3343 41383 3349
rect 41966 3340 41972 3352
rect 42024 3380 42030 3392
rect 42334 3380 42340 3392
rect 42024 3352 42340 3380
rect 42024 3340 42030 3352
rect 42334 3340 42340 3352
rect 42392 3340 42398 3392
rect 42702 3340 42708 3392
rect 42760 3340 42766 3392
rect 42889 3383 42947 3389
rect 42889 3349 42901 3383
rect 42935 3380 42947 3383
rect 45002 3380 45008 3392
rect 42935 3352 45008 3380
rect 42935 3349 42947 3352
rect 42889 3343 42947 3349
rect 45002 3340 45008 3352
rect 45060 3340 45066 3392
rect 46566 3340 46572 3392
rect 46624 3380 46630 3392
rect 46661 3383 46719 3389
rect 46661 3380 46673 3383
rect 46624 3352 46673 3380
rect 46624 3340 46630 3352
rect 46661 3349 46673 3352
rect 46707 3349 46719 3383
rect 46661 3343 46719 3349
rect 48590 3340 48596 3392
rect 48648 3380 48654 3392
rect 49142 3380 49148 3392
rect 48648 3352 49148 3380
rect 48648 3340 48654 3352
rect 49142 3340 49148 3352
rect 49200 3340 49206 3392
rect 51552 3389 51580 3420
rect 52178 3408 52184 3420
rect 52236 3408 52242 3460
rect 51537 3383 51595 3389
rect 51537 3349 51549 3383
rect 51583 3349 51595 3383
rect 51537 3343 51595 3349
rect 51629 3383 51687 3389
rect 51629 3349 51641 3383
rect 51675 3380 51687 3383
rect 52546 3380 52552 3392
rect 51675 3352 52552 3380
rect 51675 3349 51687 3352
rect 51629 3343 51687 3349
rect 52546 3340 52552 3352
rect 52604 3340 52610 3392
rect 53098 3340 53104 3392
rect 53156 3340 53162 3392
rect 54036 3380 54064 3488
rect 54214 3485 54226 3519
rect 54260 3485 54272 3519
rect 54214 3479 54272 3485
rect 54220 3448 54248 3479
rect 54294 3448 54300 3460
rect 54220 3420 54300 3448
rect 54294 3408 54300 3420
rect 54352 3408 54358 3460
rect 54496 3380 54524 3547
rect 54849 3519 54907 3525
rect 54849 3485 54861 3519
rect 54895 3485 54907 3519
rect 54849 3479 54907 3485
rect 54864 3448 54892 3479
rect 55122 3476 55128 3528
rect 55180 3476 55186 3528
rect 55214 3476 55220 3528
rect 55272 3476 55278 3528
rect 55324 3525 55352 3556
rect 55309 3519 55367 3525
rect 55309 3485 55321 3519
rect 55355 3516 55367 3519
rect 58253 3519 58311 3525
rect 58253 3516 58265 3519
rect 55355 3488 58265 3516
rect 55355 3485 55367 3488
rect 55309 3479 55367 3485
rect 58253 3485 58265 3488
rect 58299 3485 58311 3519
rect 58253 3479 58311 3485
rect 58345 3519 58403 3525
rect 58345 3485 58357 3519
rect 58391 3485 58403 3519
rect 58345 3479 58403 3485
rect 58541 3519 58599 3525
rect 58541 3485 58553 3519
rect 58587 3516 58599 3519
rect 58912 3516 58940 3896
rect 58587 3488 58940 3516
rect 58587 3485 58599 3488
rect 58541 3479 58599 3485
rect 55232 3448 55260 3476
rect 54864 3420 55260 3448
rect 55398 3408 55404 3460
rect 55456 3448 55462 3460
rect 55554 3451 55612 3457
rect 55554 3448 55566 3451
rect 55456 3420 55566 3448
rect 55456 3408 55462 3420
rect 55554 3417 55566 3420
rect 55600 3417 55612 3451
rect 58008 3451 58066 3457
rect 55554 3411 55612 3417
rect 56612 3420 57928 3448
rect 54036 3352 54524 3380
rect 54938 3340 54944 3392
rect 54996 3380 55002 3392
rect 56612 3380 56640 3420
rect 54996 3352 56640 3380
rect 56689 3383 56747 3389
rect 54996 3340 55002 3352
rect 56689 3349 56701 3383
rect 56735 3380 56747 3383
rect 56870 3380 56876 3392
rect 56735 3352 56876 3380
rect 56735 3349 56747 3352
rect 56689 3343 56747 3349
rect 56870 3340 56876 3352
rect 56928 3340 56934 3392
rect 57900 3380 57928 3420
rect 58008 3417 58020 3451
rect 58054 3448 58066 3451
rect 58158 3448 58164 3460
rect 58054 3420 58164 3448
rect 58054 3417 58066 3420
rect 58008 3411 58066 3417
rect 58158 3408 58164 3420
rect 58216 3408 58222 3460
rect 58360 3380 58388 3479
rect 57900 3352 58388 3380
rect 1104 3290 59040 3312
rect 1104 3238 15394 3290
rect 15446 3238 15458 3290
rect 15510 3238 15522 3290
rect 15574 3238 15586 3290
rect 15638 3238 15650 3290
rect 15702 3238 29838 3290
rect 29890 3238 29902 3290
rect 29954 3238 29966 3290
rect 30018 3238 30030 3290
rect 30082 3238 30094 3290
rect 30146 3238 44282 3290
rect 44334 3238 44346 3290
rect 44398 3238 44410 3290
rect 44462 3238 44474 3290
rect 44526 3238 44538 3290
rect 44590 3238 58726 3290
rect 58778 3238 58790 3290
rect 58842 3238 58854 3290
rect 58906 3238 58918 3290
rect 58970 3238 58982 3290
rect 59034 3238 59040 3290
rect 1104 3216 59040 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 1762 3176 1768 3188
rect 1719 3148 1768 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 2222 3176 2228 3188
rect 2179 3148 2228 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 3694 3176 3700 3188
rect 2547 3148 3700 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4522 3176 4528 3188
rect 4019 3148 4528 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4706 3136 4712 3188
rect 4764 3136 4770 3188
rect 7742 3136 7748 3188
rect 7800 3136 7806 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8018 3176 8024 3188
rect 7883 3148 8024 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8110 3136 8116 3188
rect 8168 3136 8174 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8570 3176 8576 3188
rect 8343 3148 8576 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10594 3176 10600 3188
rect 9456 3148 10600 3176
rect 9456 3136 9462 3148
rect 2240 3108 2268 3136
rect 2240 3080 2774 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 1627 3012 2605 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2746 3040 2774 3080
rect 3510 3068 3516 3120
rect 3568 3108 3574 3120
rect 4724 3108 4752 3136
rect 7760 3108 7788 3136
rect 3568 3080 4660 3108
rect 4724 3080 5580 3108
rect 3568 3068 3574 3080
rect 4632 3049 4660 3080
rect 5552 3049 5580 3080
rect 7024 3080 7788 3108
rect 7024 3049 7052 3080
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 2746 3012 4261 3040
rect 2593 3003 2651 3009
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 1854 2932 1860 2984
rect 1912 2932 1918 2984
rect 2038 2932 2044 2984
rect 2096 2932 2102 2984
rect 2222 2932 2228 2984
rect 2280 2932 2286 2984
rect 2342 2975 2400 2981
rect 2342 2972 2354 2975
rect 2332 2941 2354 2972
rect 2388 2941 2400 2975
rect 3237 2975 3295 2981
rect 2332 2935 2400 2941
rect 2608 2944 3188 2972
rect 2056 2904 2084 2932
rect 2332 2904 2360 2935
rect 2608 2904 2636 2944
rect 2056 2876 2636 2904
rect 3160 2836 3188 2944
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 4154 2972 4160 2984
rect 3467 2944 4160 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 3252 2904 3280 2935
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 3694 2904 3700 2916
rect 3252 2876 3700 2904
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 5368 2904 5396 3003
rect 7098 3000 7104 3052
rect 7156 3000 7162 3052
rect 7650 3000 7656 3052
rect 7708 3000 7714 3052
rect 8128 3040 8156 3136
rect 9232 3049 9260 3136
rect 9585 3111 9643 3117
rect 9585 3077 9597 3111
rect 9631 3108 9643 3111
rect 9674 3108 9680 3120
rect 9631 3080 9680 3108
rect 9631 3077 9643 3080
rect 9585 3071 9643 3077
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 9784 3117 9812 3148
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 10928 3148 11621 3176
rect 10928 3136 10934 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 11609 3139 11667 3145
rect 12406 3148 13553 3176
rect 9769 3111 9827 3117
rect 9769 3077 9781 3111
rect 9815 3077 9827 3111
rect 9769 3071 9827 3077
rect 9861 3111 9919 3117
rect 9861 3077 9873 3111
rect 9907 3108 9919 3111
rect 10226 3108 10232 3120
rect 9907 3080 10232 3108
rect 9907 3077 9919 3080
rect 9861 3071 9919 3077
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10781 3111 10839 3117
rect 10781 3077 10793 3111
rect 10827 3108 10839 3111
rect 12406 3108 12434 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13541 3139 13599 3145
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14424 3148 14473 3176
rect 14424 3136 14430 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 14461 3139 14519 3145
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15746 3176 15752 3188
rect 15436 3148 15752 3176
rect 15436 3136 15442 3148
rect 15746 3136 15752 3148
rect 15804 3176 15810 3188
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 15804 3148 15945 3176
rect 15804 3136 15810 3148
rect 15933 3145 15945 3148
rect 15979 3145 15991 3179
rect 16206 3176 16212 3188
rect 15933 3139 15991 3145
rect 16040 3148 16212 3176
rect 10827 3080 12434 3108
rect 10827 3077 10839 3080
rect 10781 3071 10839 3077
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 14182 3108 14188 3120
rect 13136 3080 14188 3108
rect 13136 3068 13142 3080
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 16040 3117 16068 3148
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16298 3136 16304 3188
rect 16356 3136 16362 3188
rect 16482 3136 16488 3188
rect 16540 3176 16546 3188
rect 16540 3148 16896 3176
rect 16540 3136 16546 3148
rect 14798 3111 14856 3117
rect 14798 3108 14810 3111
rect 14700 3080 14810 3108
rect 14700 3068 14706 3080
rect 14798 3077 14810 3080
rect 14844 3077 14856 3111
rect 14798 3071 14856 3077
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3077 16083 3111
rect 16316 3108 16344 3136
rect 16025 3071 16083 3077
rect 16132 3080 16344 3108
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 7760 3012 8401 3040
rect 6362 2932 6368 2984
rect 6420 2932 6426 2984
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7760 2972 7788 3012
rect 8389 3009 8401 3012
rect 8435 3040 8447 3043
rect 9217 3043 9275 3049
rect 8435 3012 8984 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 7423 2944 7788 2972
rect 8021 2975 8079 2981
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 8021 2941 8033 2975
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 4028 2876 5396 2904
rect 6181 2907 6239 2913
rect 4028 2864 4034 2876
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 6730 2904 6736 2916
rect 6227 2876 6736 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 6730 2864 6736 2876
rect 6788 2904 6794 2916
rect 8036 2904 8064 2935
rect 8110 2932 8116 2984
rect 8168 2932 8174 2984
rect 8956 2981 8984 3012
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9950 3040 9956 3052
rect 10008 3049 10014 3052
rect 9217 3003 9275 3009
rect 9646 3012 9956 3040
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 9646 2972 9674 3012
rect 9950 3000 9956 3012
rect 10008 3040 10016 3049
rect 10008 3012 10053 3040
rect 10008 3003 10016 3012
rect 10008 3000 10014 3003
rect 10134 3000 10140 3052
rect 10192 3000 10198 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 10686 3040 10692 3052
rect 10551 3012 10692 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14458 3040 14464 3052
rect 13771 3012 14464 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14550 3000 14556 3052
rect 14608 3000 14614 3052
rect 8987 2944 9674 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 9858 2932 9864 2984
rect 9916 2932 9922 2984
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10284 2944 10885 2972
rect 10284 2932 10290 2944
rect 10873 2941 10885 2944
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 12032 2944 12541 2972
rect 12032 2932 12038 2944
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 16132 2981 16160 3080
rect 16574 3068 16580 3120
rect 16632 3068 16638 3120
rect 16666 3068 16672 3120
rect 16724 3068 16730 3120
rect 16868 3108 16896 3148
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 17957 3179 18015 3185
rect 17957 3176 17969 3179
rect 17092 3148 17969 3176
rect 17092 3136 17098 3148
rect 17957 3145 17969 3148
rect 18003 3145 18015 3179
rect 17957 3139 18015 3145
rect 19153 3179 19211 3185
rect 19153 3145 19165 3179
rect 19199 3176 19211 3179
rect 19518 3176 19524 3188
rect 19199 3148 19524 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 20070 3136 20076 3188
rect 20128 3136 20134 3188
rect 20901 3179 20959 3185
rect 20901 3145 20913 3179
rect 20947 3176 20959 3179
rect 20990 3176 20996 3188
rect 20947 3148 20996 3176
rect 20947 3145 20959 3148
rect 20901 3139 20959 3145
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 21542 3136 21548 3188
rect 21600 3176 21606 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21600 3148 21833 3176
rect 21600 3136 21606 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 23382 3176 23388 3188
rect 21821 3139 21879 3145
rect 22664 3148 23388 3176
rect 20088 3108 20116 3136
rect 22664 3117 22692 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 24029 3179 24087 3185
rect 24029 3145 24041 3179
rect 24075 3176 24087 3179
rect 24118 3176 24124 3188
rect 24075 3148 24124 3176
rect 24075 3145 24087 3148
rect 24029 3139 24087 3145
rect 24118 3136 24124 3148
rect 24176 3136 24182 3188
rect 25038 3136 25044 3188
rect 25096 3136 25102 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 25685 3179 25743 3185
rect 25685 3176 25697 3179
rect 25280 3148 25697 3176
rect 25280 3136 25286 3148
rect 25685 3145 25697 3148
rect 25731 3145 25743 3179
rect 25685 3139 25743 3145
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 26973 3179 27031 3185
rect 26973 3176 26985 3179
rect 26568 3148 26985 3176
rect 26568 3136 26574 3148
rect 26973 3145 26985 3148
rect 27019 3145 27031 3179
rect 26973 3139 27031 3145
rect 29270 3136 29276 3188
rect 29328 3136 29334 3188
rect 30650 3136 30656 3188
rect 30708 3176 30714 3188
rect 31021 3179 31079 3185
rect 31021 3176 31033 3179
rect 30708 3148 31033 3176
rect 30708 3136 30714 3148
rect 31021 3145 31033 3148
rect 31067 3145 31079 3179
rect 31021 3139 31079 3145
rect 31386 3136 31392 3188
rect 31444 3176 31450 3188
rect 32217 3179 32275 3185
rect 32217 3176 32229 3179
rect 31444 3148 32229 3176
rect 31444 3136 31450 3148
rect 32217 3145 32229 3148
rect 32263 3145 32275 3179
rect 32217 3139 32275 3145
rect 32858 3136 32864 3188
rect 32916 3136 32922 3188
rect 33689 3179 33747 3185
rect 33689 3145 33701 3179
rect 33735 3176 33747 3179
rect 34330 3176 34336 3188
rect 33735 3148 34336 3176
rect 33735 3145 33747 3148
rect 33689 3139 33747 3145
rect 34330 3136 34336 3148
rect 34388 3136 34394 3188
rect 34790 3136 34796 3188
rect 34848 3136 34854 3188
rect 34882 3136 34888 3188
rect 34940 3136 34946 3188
rect 35342 3136 35348 3188
rect 35400 3136 35406 3188
rect 35710 3136 35716 3188
rect 35768 3176 35774 3188
rect 36081 3179 36139 3185
rect 36081 3176 36093 3179
rect 35768 3148 36093 3176
rect 35768 3136 35774 3148
rect 36081 3145 36093 3148
rect 36127 3145 36139 3179
rect 36081 3139 36139 3145
rect 36998 3136 37004 3188
rect 37056 3136 37062 3188
rect 38194 3136 38200 3188
rect 38252 3136 38258 3188
rect 38930 3136 38936 3188
rect 38988 3176 38994 3188
rect 39025 3179 39083 3185
rect 39025 3176 39037 3179
rect 38988 3148 39037 3176
rect 38988 3136 38994 3148
rect 39025 3145 39037 3148
rect 39071 3145 39083 3179
rect 39025 3139 39083 3145
rect 39390 3136 39396 3188
rect 39448 3176 39454 3188
rect 40678 3176 40684 3188
rect 39448 3148 40684 3176
rect 39448 3136 39454 3148
rect 40678 3136 40684 3148
rect 40736 3136 40742 3188
rect 41230 3136 41236 3188
rect 41288 3136 41294 3188
rect 41414 3136 41420 3188
rect 41472 3176 41478 3188
rect 42429 3179 42487 3185
rect 42429 3176 42441 3179
rect 41472 3148 42441 3176
rect 41472 3136 41478 3148
rect 42429 3145 42441 3148
rect 42475 3145 42487 3179
rect 42429 3139 42487 3145
rect 43162 3136 43168 3188
rect 43220 3176 43226 3188
rect 43349 3179 43407 3185
rect 43349 3176 43361 3179
rect 43220 3148 43361 3176
rect 43220 3136 43226 3148
rect 43349 3145 43361 3148
rect 43395 3145 43407 3179
rect 43349 3139 43407 3145
rect 46198 3136 46204 3188
rect 46256 3136 46262 3188
rect 46934 3136 46940 3188
rect 46992 3136 46998 3188
rect 47118 3136 47124 3188
rect 47176 3176 47182 3188
rect 47581 3179 47639 3185
rect 47581 3176 47593 3179
rect 47176 3148 47593 3176
rect 47176 3136 47182 3148
rect 47581 3145 47593 3148
rect 47627 3145 47639 3179
rect 48682 3176 48688 3188
rect 47581 3139 47639 3145
rect 48516 3148 48688 3176
rect 21361 3111 21419 3117
rect 16868 3080 18184 3108
rect 20088 3080 21220 3108
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 16398 3043 16456 3049
rect 16398 3009 16410 3043
rect 16444 3040 16456 3043
rect 16592 3040 16620 3068
rect 16444 3012 16620 3040
rect 16444 3009 16456 3012
rect 16398 3003 16456 3009
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 13688 2944 13829 2972
rect 13688 2932 13694 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2941 16175 2975
rect 16316 2972 16344 3003
rect 16684 2972 16712 3068
rect 17126 3000 17132 3052
rect 17184 3000 17190 3052
rect 17310 3000 17316 3052
rect 17368 3000 17374 3052
rect 18156 3049 18184 3080
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 16316 2944 16712 2972
rect 17221 2975 17279 2981
rect 16117 2935 16175 2941
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 6788 2876 8064 2904
rect 6788 2864 6794 2876
rect 10318 2864 10324 2916
rect 10376 2864 10382 2916
rect 11256 2876 12434 2904
rect 3510 2836 3516 2848
rect 3160 2808 3516 2836
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 5169 2839 5227 2845
rect 5169 2805 5181 2839
rect 5215 2836 5227 2839
rect 7098 2836 7104 2848
rect 5215 2808 7104 2836
rect 5215 2805 5227 2808
rect 5169 2799 5227 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 11256 2845 11284 2876
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7892 2808 8217 2836
rect 7892 2796 7898 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2836 10747 2839
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 10735 2808 10793 2836
rect 10735 2805 10747 2808
rect 10689 2799 10747 2805
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 10781 2799 10839 2805
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2805 11299 2839
rect 12406 2836 12434 2876
rect 16022 2864 16028 2916
rect 16080 2904 16086 2916
rect 17236 2904 17264 2935
rect 16080 2876 17264 2904
rect 16080 2864 16086 2876
rect 17328 2836 17356 3000
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 17911 2944 18245 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 18432 2904 18460 3003
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 19116 3012 19257 3040
rect 19116 3000 19122 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 21082 3000 21088 3052
rect 21140 3000 21146 3052
rect 21192 3040 21220 3080
rect 21361 3077 21373 3111
rect 21407 3108 21419 3111
rect 22649 3111 22707 3117
rect 21407 3080 21864 3108
rect 21407 3077 21419 3080
rect 21361 3071 21419 3077
rect 21836 3052 21864 3080
rect 22649 3077 22661 3111
rect 22695 3077 22707 3111
rect 22649 3071 22707 3077
rect 22738 3068 22744 3120
rect 22796 3108 22802 3120
rect 22833 3111 22891 3117
rect 22833 3108 22845 3111
rect 22796 3080 22845 3108
rect 22796 3068 22802 3080
rect 22833 3077 22845 3080
rect 22879 3077 22891 3111
rect 22833 3071 22891 3077
rect 22925 3111 22983 3117
rect 22925 3077 22937 3111
rect 22971 3108 22983 3111
rect 22971 3080 24256 3108
rect 22971 3077 22983 3080
rect 22925 3071 22983 3077
rect 24228 3052 24256 3080
rect 24302 3068 24308 3120
rect 24360 3108 24366 3120
rect 24670 3108 24676 3120
rect 24360 3080 24676 3108
rect 24360 3068 24366 3080
rect 24670 3068 24676 3080
rect 24728 3068 24734 3120
rect 21248 3043 21306 3049
rect 21248 3040 21260 3043
rect 21192 3012 21260 3040
rect 21248 3009 21260 3012
rect 21294 3040 21306 3043
rect 21294 3012 21404 3040
rect 21294 3009 21306 3012
rect 21248 3003 21306 3009
rect 18598 2932 18604 2984
rect 18656 2932 18662 2984
rect 19150 2932 19156 2984
rect 19208 2972 19214 2984
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 19208 2944 19717 2972
rect 19208 2932 19214 2944
rect 19705 2941 19717 2944
rect 19751 2941 19763 2975
rect 21376 2972 21404 3012
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 21634 3000 21640 3052
rect 21692 3000 21698 3052
rect 21818 3000 21824 3052
rect 21876 3000 21882 3052
rect 23022 3043 23080 3049
rect 23022 3040 23034 3043
rect 21928 3012 23034 3040
rect 21928 2972 21956 3012
rect 23022 3009 23034 3012
rect 23068 3040 23080 3043
rect 23290 3040 23296 3052
rect 23068 3012 23296 3040
rect 23068 3009 23080 3012
rect 23022 3003 23080 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23937 3043 23995 3049
rect 23937 3009 23949 3043
rect 23983 3040 23995 3043
rect 24026 3040 24032 3052
rect 23983 3012 24032 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 24026 3000 24032 3012
rect 24084 3000 24090 3052
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 21376 2944 21956 2972
rect 22066 2944 22385 2972
rect 19705 2935 19763 2941
rect 20622 2904 20628 2916
rect 18432 2876 20628 2904
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 21637 2907 21695 2913
rect 21637 2873 21649 2907
rect 21683 2904 21695 2907
rect 22066 2904 22094 2944
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 22741 2975 22799 2981
rect 22741 2941 22753 2975
rect 22787 2972 22799 2975
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 22787 2944 23765 2972
rect 22787 2941 22799 2944
rect 22741 2935 22799 2941
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 24136 2972 24164 3003
rect 24210 3000 24216 3052
rect 24268 3000 24274 3052
rect 25056 3040 25084 3136
rect 29288 3049 29316 3136
rect 32876 3108 32904 3136
rect 33137 3111 33195 3117
rect 33137 3108 33149 3111
rect 32876 3080 33149 3108
rect 24320 3012 25084 3040
rect 26697 3043 26755 3049
rect 24320 2972 24348 3012
rect 26697 3009 26709 3043
rect 26743 3040 26755 3043
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 26743 3012 27721 3040
rect 26743 3009 26755 3012
rect 26697 3003 26755 3009
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 30926 3000 30932 3052
rect 30984 3000 30990 3052
rect 31202 3000 31208 3052
rect 31260 3000 31266 3052
rect 32876 3040 32904 3080
rect 33137 3077 33149 3080
rect 33183 3077 33195 3111
rect 33137 3071 33195 3077
rect 33410 3049 33416 3052
rect 33403 3043 33416 3049
rect 33403 3040 33415 3043
rect 32784 3012 32904 3040
rect 33371 3012 33415 3040
rect 24136 2944 24348 2972
rect 23753 2935 23811 2941
rect 24670 2932 24676 2984
rect 24728 2932 24734 2984
rect 26237 2975 26295 2981
rect 26237 2941 26249 2975
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 21683 2876 22094 2904
rect 21683 2873 21695 2876
rect 21637 2867 21695 2873
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 26252 2904 26280 2935
rect 27614 2932 27620 2984
rect 27672 2932 27678 2984
rect 28261 2975 28319 2981
rect 28261 2941 28273 2975
rect 28307 2941 28319 2975
rect 28261 2935 28319 2941
rect 23624 2876 26280 2904
rect 26513 2907 26571 2913
rect 23624 2864 23630 2876
rect 26513 2873 26525 2907
rect 26559 2904 26571 2907
rect 26694 2904 26700 2916
rect 26559 2876 26700 2904
rect 26559 2873 26571 2876
rect 26513 2867 26571 2873
rect 26694 2864 26700 2876
rect 26752 2864 26758 2916
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 28276 2904 28304 2935
rect 28534 2932 28540 2984
rect 28592 2932 28598 2984
rect 29362 2932 29368 2984
rect 29420 2972 29426 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 29420 2944 29653 2972
rect 29420 2932 29426 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 30558 2932 30564 2984
rect 30616 2972 30622 2984
rect 31389 2975 31447 2981
rect 30616 2944 30788 2972
rect 30616 2932 30622 2944
rect 30760 2913 30788 2944
rect 31389 2941 31401 2975
rect 31435 2972 31447 2975
rect 31846 2972 31852 2984
rect 31435 2944 31852 2972
rect 31435 2941 31447 2944
rect 31389 2935 31447 2941
rect 31846 2932 31852 2944
rect 31904 2932 31910 2984
rect 26936 2876 28304 2904
rect 30745 2907 30803 2913
rect 26936 2864 26942 2876
rect 30745 2873 30757 2907
rect 30791 2873 30803 2907
rect 30745 2867 30803 2873
rect 12406 2808 17356 2836
rect 18417 2839 18475 2845
rect 11241 2799 11299 2805
rect 18417 2805 18429 2839
rect 18463 2836 18475 2839
rect 18782 2836 18788 2848
rect 18463 2808 18788 2836
rect 18463 2805 18475 2808
rect 18417 2799 18475 2805
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 21726 2796 21732 2848
rect 21784 2836 21790 2848
rect 23201 2839 23259 2845
rect 23201 2836 23213 2839
rect 21784 2808 23213 2836
rect 21784 2796 21790 2808
rect 23201 2805 23213 2808
rect 23247 2805 23259 2839
rect 23201 2799 23259 2805
rect 29086 2796 29092 2848
rect 29144 2796 29150 2848
rect 31938 2796 31944 2848
rect 31996 2796 32002 2848
rect 32784 2836 32812 3012
rect 33403 3009 33415 3012
rect 33403 3003 33416 3009
rect 33410 3000 33416 3003
rect 33468 3000 33474 3052
rect 33505 3043 33563 3049
rect 33505 3009 33517 3043
rect 33551 3040 33563 3043
rect 33873 3043 33931 3049
rect 33873 3040 33885 3043
rect 33551 3012 33885 3040
rect 33551 3009 33563 3012
rect 33505 3003 33563 3009
rect 33873 3009 33885 3012
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 34609 3043 34667 3049
rect 34609 3009 34621 3043
rect 34655 3040 34667 3043
rect 34808 3040 34836 3136
rect 34655 3012 34836 3040
rect 34900 3040 34928 3136
rect 35360 3108 35388 3136
rect 35360 3080 36400 3108
rect 36372 3049 36400 3080
rect 35897 3043 35955 3049
rect 34900 3012 35388 3040
rect 34655 3009 34667 3012
rect 34609 3003 34667 3009
rect 32861 2975 32919 2981
rect 32861 2941 32873 2975
rect 32907 2972 32919 2975
rect 33134 2972 33140 2984
rect 32907 2944 33140 2972
rect 32907 2941 32919 2944
rect 32861 2935 32919 2941
rect 33134 2932 33140 2944
rect 33192 2932 33198 2984
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 34425 2975 34483 2981
rect 34425 2972 34437 2975
rect 33652 2944 34437 2972
rect 33652 2932 33658 2944
rect 34425 2941 34437 2944
rect 34471 2941 34483 2975
rect 34425 2935 34483 2941
rect 34885 2975 34943 2981
rect 34885 2941 34897 2975
rect 34931 2972 34943 2975
rect 35066 2972 35072 2984
rect 34931 2944 35072 2972
rect 34931 2941 34943 2944
rect 34885 2935 34943 2941
rect 35066 2932 35072 2944
rect 35124 2932 35130 2984
rect 35250 2932 35256 2984
rect 35308 2932 35314 2984
rect 35360 2972 35388 3012
rect 35897 3009 35909 3043
rect 35943 3040 35955 3043
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 35943 3012 36277 3040
rect 35943 3009 35955 3012
rect 35897 3003 35955 3009
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 36357 3043 36415 3049
rect 36357 3009 36369 3043
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 36538 3000 36544 3052
rect 36596 3000 36602 3052
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 37553 3043 37611 3049
rect 37553 3009 37565 3043
rect 37599 3040 37611 3043
rect 38212 3040 38240 3136
rect 39298 3068 39304 3120
rect 39356 3068 39362 3120
rect 37599 3012 38240 3040
rect 37599 3009 37611 3012
rect 37553 3003 37611 3009
rect 39206 3000 39212 3052
rect 39264 3000 39270 3052
rect 36449 2975 36507 2981
rect 36449 2972 36461 2975
rect 35360 2944 36461 2972
rect 36449 2941 36461 2944
rect 36495 2941 36507 2975
rect 36449 2935 36507 2941
rect 32950 2864 32956 2916
rect 33008 2904 33014 2916
rect 36170 2904 36176 2916
rect 33008 2876 36176 2904
rect 33008 2864 33014 2876
rect 36170 2864 36176 2876
rect 36228 2864 36234 2916
rect 34698 2836 34704 2848
rect 32784 2808 34704 2836
rect 34698 2796 34704 2808
rect 34756 2836 34762 2848
rect 36556 2836 36584 3000
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37700 2944 37933 2972
rect 37700 2932 37706 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 39316 2972 39344 3068
rect 39408 3040 39436 3136
rect 39577 3111 39635 3117
rect 39577 3077 39589 3111
rect 39623 3108 39635 3111
rect 39623 3080 41000 3108
rect 39623 3077 39635 3080
rect 39577 3071 39635 3077
rect 39464 3043 39522 3049
rect 39464 3040 39476 3043
rect 39408 3012 39476 3040
rect 39464 3009 39476 3012
rect 39510 3009 39522 3043
rect 39464 3003 39522 3009
rect 39669 3043 39727 3049
rect 39669 3009 39681 3043
rect 39715 3009 39727 3043
rect 39669 3003 39727 3009
rect 39853 3043 39911 3049
rect 39853 3009 39865 3043
rect 39899 3040 39911 3043
rect 40218 3040 40224 3052
rect 39899 3012 40224 3040
rect 39899 3009 39911 3012
rect 39853 3003 39911 3009
rect 39684 2972 39712 3003
rect 40218 3000 40224 3012
rect 40276 3000 40282 3052
rect 40972 3049 41000 3080
rect 40957 3043 41015 3049
rect 40957 3009 40969 3043
rect 41003 3040 41015 3043
rect 41248 3040 41276 3136
rect 41003 3012 41276 3040
rect 41003 3009 41015 3012
rect 40957 3003 41015 3009
rect 43622 3000 43628 3052
rect 43680 3040 43686 3052
rect 43901 3043 43959 3049
rect 43901 3040 43913 3043
rect 43680 3012 43913 3040
rect 43680 3000 43686 3012
rect 43901 3009 43913 3012
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 44818 3000 44824 3052
rect 44876 3040 44882 3052
rect 45281 3043 45339 3049
rect 45281 3040 45293 3043
rect 44876 3012 45293 3040
rect 44876 3000 44882 3012
rect 45281 3009 45293 3012
rect 45327 3009 45339 3043
rect 46216 3040 46244 3136
rect 46569 3111 46627 3117
rect 46569 3077 46581 3111
rect 46615 3108 46627 3111
rect 46658 3108 46664 3120
rect 46615 3080 46664 3108
rect 46615 3077 46627 3080
rect 46569 3071 46627 3077
rect 46658 3068 46664 3080
rect 46716 3068 46722 3120
rect 46750 3068 46756 3120
rect 46808 3068 46814 3120
rect 46842 3068 46848 3120
rect 46900 3108 46906 3120
rect 46900 3080 47256 3108
rect 46900 3068 46906 3080
rect 47228 3049 47256 3080
rect 48314 3068 48320 3120
rect 48372 3068 48378 3120
rect 48516 3117 48544 3148
rect 48682 3136 48688 3148
rect 48740 3136 48746 3188
rect 48958 3176 48964 3188
rect 48792 3148 48964 3176
rect 48501 3111 48559 3117
rect 48501 3077 48513 3111
rect 48547 3077 48559 3111
rect 48501 3071 48559 3077
rect 46349 3043 46407 3049
rect 46349 3040 46361 3043
rect 46216 3012 46361 3040
rect 45281 3003 45339 3009
rect 46349 3009 46361 3012
rect 46395 3009 46407 3043
rect 46349 3003 46407 3009
rect 46477 3043 46535 3049
rect 46477 3009 46489 3043
rect 46523 3040 46535 3043
rect 47121 3043 47179 3049
rect 47121 3040 47133 3043
rect 46523 3012 46612 3040
rect 46523 3009 46535 3012
rect 46477 3003 46535 3009
rect 46584 2984 46612 3012
rect 46676 3012 47133 3040
rect 39316 2944 39712 2972
rect 39761 2975 39819 2981
rect 37921 2935 37979 2941
rect 39761 2941 39773 2975
rect 39807 2972 39819 2975
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 39807 2944 40509 2972
rect 39807 2941 39819 2944
rect 39761 2935 39819 2941
rect 40497 2941 40509 2944
rect 40543 2941 40555 2975
rect 40497 2935 40555 2941
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41233 2975 41291 2981
rect 41233 2972 41245 2975
rect 40736 2944 41245 2972
rect 40736 2932 40742 2944
rect 41233 2941 41245 2944
rect 41279 2941 41291 2975
rect 41233 2935 41291 2941
rect 41782 2932 41788 2984
rect 41840 2972 41846 2984
rect 42981 2975 43039 2981
rect 42981 2972 42993 2975
rect 41840 2944 42993 2972
rect 41840 2932 41846 2944
rect 42981 2941 42993 2944
rect 43027 2941 43039 2975
rect 42981 2935 43039 2941
rect 43990 2932 43996 2984
rect 44048 2972 44054 2984
rect 44269 2975 44327 2981
rect 44269 2972 44281 2975
rect 44048 2944 44281 2972
rect 44048 2932 44054 2944
rect 44269 2941 44281 2944
rect 44315 2941 44327 2975
rect 44269 2935 44327 2941
rect 45094 2932 45100 2984
rect 45152 2972 45158 2984
rect 45557 2975 45615 2981
rect 45557 2972 45569 2975
rect 45152 2944 45569 2972
rect 45152 2932 45158 2944
rect 45557 2941 45569 2944
rect 45603 2941 45615 2975
rect 45557 2935 45615 2941
rect 46566 2932 46572 2984
rect 46624 2932 46630 2984
rect 46201 2907 46259 2913
rect 46201 2873 46213 2907
rect 46247 2904 46259 2907
rect 46676 2904 46704 3012
rect 47121 3009 47133 3012
rect 47167 3009 47179 3043
rect 47121 3003 47179 3009
rect 47213 3043 47271 3049
rect 47213 3009 47225 3043
rect 47259 3009 47271 3043
rect 48516 3040 48544 3071
rect 48590 3068 48596 3120
rect 48648 3068 48654 3120
rect 47213 3003 47271 3009
rect 47320 3012 48544 3040
rect 48705 3065 48763 3071
rect 48705 3031 48717 3065
rect 48751 3062 48763 3065
rect 48792 3062 48820 3148
rect 48958 3136 48964 3148
rect 49016 3136 49022 3188
rect 51902 3136 51908 3188
rect 51960 3176 51966 3188
rect 52273 3179 52331 3185
rect 52273 3176 52285 3179
rect 51960 3148 52285 3176
rect 51960 3136 51966 3148
rect 52273 3145 52285 3148
rect 52319 3145 52331 3179
rect 52273 3139 52331 3145
rect 53116 3148 54055 3176
rect 53116 3120 53144 3148
rect 51074 3068 51080 3120
rect 51132 3108 51138 3120
rect 51445 3111 51503 3117
rect 51445 3108 51457 3111
rect 51132 3080 51457 3108
rect 51132 3068 51138 3080
rect 51445 3077 51457 3080
rect 51491 3077 51503 3111
rect 51445 3071 51503 3077
rect 51721 3111 51779 3117
rect 51721 3077 51733 3111
rect 51767 3108 51779 3111
rect 52546 3108 52552 3120
rect 51767 3080 52552 3108
rect 51767 3077 51779 3080
rect 51721 3071 51779 3077
rect 52546 3068 52552 3080
rect 52604 3068 52610 3120
rect 53098 3068 53104 3120
rect 53156 3068 53162 3120
rect 53469 3111 53527 3117
rect 53469 3077 53481 3111
rect 53515 3108 53527 3111
rect 53558 3108 53564 3120
rect 53515 3080 53564 3108
rect 53515 3077 53527 3080
rect 53469 3071 53527 3077
rect 53558 3068 53564 3080
rect 53616 3068 53622 3120
rect 53650 3068 53656 3120
rect 53708 3068 53714 3120
rect 53760 3117 53788 3148
rect 53745 3111 53803 3117
rect 53745 3077 53757 3111
rect 53791 3077 53803 3111
rect 53745 3071 53803 3077
rect 48751 3034 48820 3062
rect 49050 3040 49056 3052
rect 48751 3031 48763 3034
rect 48705 3025 48763 3031
rect 48884 3012 49056 3040
rect 46750 2932 46756 2984
rect 46808 2972 46814 2984
rect 47320 2972 47348 3012
rect 46808 2944 47348 2972
rect 48133 2975 48191 2981
rect 46808 2932 46814 2944
rect 48133 2941 48145 2975
rect 48179 2941 48191 2975
rect 48133 2935 48191 2941
rect 48593 2975 48651 2981
rect 48593 2941 48605 2975
rect 48639 2972 48651 2975
rect 48884 2972 48912 3012
rect 49050 3000 49056 3012
rect 49108 3000 49114 3052
rect 49142 3000 49148 3052
rect 49200 3000 49206 3052
rect 51350 3000 51356 3052
rect 51408 3000 51414 3052
rect 51629 3043 51687 3049
rect 51629 3009 51641 3043
rect 51675 3009 51687 3043
rect 51629 3003 51687 3009
rect 51849 3043 51907 3049
rect 51849 3009 51861 3043
rect 51895 3040 51907 3043
rect 51994 3040 52000 3052
rect 51895 3012 52000 3040
rect 51895 3009 51907 3012
rect 51849 3003 51907 3009
rect 48639 2944 48912 2972
rect 48639 2941 48651 2944
rect 48593 2935 48651 2941
rect 46247 2876 46704 2904
rect 46247 2873 46259 2876
rect 46201 2867 46259 2873
rect 46934 2864 46940 2916
rect 46992 2904 46998 2916
rect 48148 2904 48176 2935
rect 48958 2932 48964 2984
rect 49016 2972 49022 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 49016 2944 49525 2972
rect 49016 2932 49022 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 50062 2932 50068 2984
rect 50120 2972 50126 2984
rect 50525 2975 50583 2981
rect 50525 2972 50537 2975
rect 50120 2944 50537 2972
rect 50120 2932 50126 2944
rect 50525 2941 50537 2944
rect 50571 2941 50583 2975
rect 51368 2972 51396 3000
rect 51445 2975 51503 2981
rect 51445 2972 51457 2975
rect 51368 2944 51457 2972
rect 50525 2935 50583 2941
rect 51445 2941 51457 2944
rect 51491 2941 51503 2975
rect 51445 2935 51503 2941
rect 46992 2876 48176 2904
rect 46992 2864 46998 2876
rect 49418 2864 49424 2916
rect 49476 2864 49482 2916
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 51644 2904 51672 3003
rect 51994 3000 52000 3012
rect 52052 3000 52058 3052
rect 52457 3043 52515 3049
rect 52457 3009 52469 3043
rect 52503 3040 52515 3043
rect 52733 3043 52791 3049
rect 52733 3040 52745 3043
rect 52503 3012 52745 3040
rect 52503 3009 52515 3012
rect 52457 3003 52515 3009
rect 52733 3009 52745 3012
rect 52779 3009 52791 3043
rect 52733 3003 52791 3009
rect 51718 2932 51724 2984
rect 51776 2972 51782 2984
rect 53285 2975 53343 2981
rect 53285 2972 53297 2975
rect 51776 2944 53297 2972
rect 51776 2932 51782 2944
rect 53285 2941 53297 2944
rect 53331 2941 53343 2975
rect 53285 2935 53343 2941
rect 53668 2904 53696 3068
rect 53834 3000 53840 3052
rect 53892 3039 53898 3052
rect 54027 3049 54055 3148
rect 58526 3136 58532 3188
rect 58584 3136 58590 3188
rect 54021 3043 54079 3049
rect 53892 3033 53931 3039
rect 53873 2999 53885 3000
rect 53919 2999 53931 3033
rect 54021 3009 54033 3043
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 57698 3000 57704 3052
rect 57756 3000 57762 3052
rect 53873 2993 53931 2999
rect 53742 2932 53748 2984
rect 53800 2932 53806 2984
rect 54202 2932 54208 2984
rect 54260 2972 54266 2984
rect 54481 2975 54539 2981
rect 54481 2972 54493 2975
rect 54260 2944 54493 2972
rect 54260 2932 54266 2944
rect 54481 2941 54493 2944
rect 54527 2941 54539 2975
rect 54481 2935 54539 2941
rect 55030 2932 55036 2984
rect 55088 2972 55094 2984
rect 55493 2975 55551 2981
rect 55493 2972 55505 2975
rect 55088 2944 55505 2972
rect 55088 2932 55094 2944
rect 55493 2941 55505 2944
rect 55539 2941 55551 2975
rect 55493 2935 55551 2941
rect 57238 2932 57244 2984
rect 57296 2932 57302 2984
rect 57977 2975 58035 2981
rect 57977 2941 57989 2975
rect 58023 2972 58035 2975
rect 58342 2972 58348 2984
rect 58023 2944 58348 2972
rect 58023 2941 58035 2944
rect 57977 2935 58035 2941
rect 58342 2932 58348 2944
rect 58400 2932 58406 2984
rect 51040 2876 53696 2904
rect 51040 2864 51046 2876
rect 38654 2836 38660 2848
rect 34756 2808 38660 2836
rect 34756 2796 34762 2808
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 39758 2796 39764 2848
rect 39816 2836 39822 2848
rect 39945 2839 40003 2845
rect 39945 2836 39957 2839
rect 39816 2808 39957 2836
rect 39816 2796 39822 2808
rect 39945 2805 39957 2808
rect 39991 2805 40003 2839
rect 39945 2799 40003 2805
rect 43438 2796 43444 2848
rect 43496 2836 43502 2848
rect 45554 2836 45560 2848
rect 43496 2808 45560 2836
rect 43496 2796 43502 2808
rect 45554 2796 45560 2808
rect 45612 2796 45618 2848
rect 46290 2796 46296 2848
rect 46348 2836 46354 2848
rect 46753 2839 46811 2845
rect 46753 2836 46765 2839
rect 46348 2808 46765 2836
rect 46348 2796 46354 2808
rect 46753 2805 46765 2808
rect 46799 2805 46811 2839
rect 46753 2799 46811 2805
rect 47397 2839 47455 2845
rect 47397 2805 47409 2839
rect 47443 2836 47455 2839
rect 49436 2836 49464 2864
rect 47443 2808 49464 2836
rect 47443 2805 47455 2808
rect 47397 2799 47455 2805
rect 51166 2796 51172 2848
rect 51224 2796 51230 2848
rect 56137 2839 56195 2845
rect 56137 2805 56149 2839
rect 56183 2836 56195 2839
rect 56962 2836 56968 2848
rect 56183 2808 56968 2836
rect 56183 2805 56195 2808
rect 56137 2799 56195 2805
rect 56962 2796 56968 2808
rect 57020 2796 57026 2848
rect 1104 2746 58880 2768
rect 1104 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 22616 2746
rect 22668 2694 22680 2746
rect 22732 2694 22744 2746
rect 22796 2694 22808 2746
rect 22860 2694 22872 2746
rect 22924 2694 37060 2746
rect 37112 2694 37124 2746
rect 37176 2694 37188 2746
rect 37240 2694 37252 2746
rect 37304 2694 37316 2746
rect 37368 2694 51504 2746
rect 51556 2694 51568 2746
rect 51620 2694 51632 2746
rect 51684 2694 51696 2746
rect 51748 2694 51760 2746
rect 51812 2694 58880 2746
rect 1104 2672 58880 2694
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 4890 2632 4896 2644
rect 4755 2604 4896 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 7285 2635 7343 2641
rect 6595 2604 6914 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2564 4031 2567
rect 6886 2564 6914 2604
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7650 2632 7656 2644
rect 7331 2604 7656 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10134 2632 10140 2644
rect 9815 2604 10140 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10226 2592 10232 2644
rect 10284 2592 10290 2644
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 11848 2604 12173 2632
rect 11848 2592 11854 2604
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12161 2595 12219 2601
rect 12253 2635 12311 2641
rect 12253 2601 12265 2635
rect 12299 2632 12311 2635
rect 12342 2632 12348 2644
rect 12299 2604 12348 2632
rect 12299 2601 12311 2604
rect 12253 2595 12311 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14826 2632 14832 2644
rect 14415 2604 14832 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 16022 2592 16028 2644
rect 16080 2592 16086 2644
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 17497 2635 17555 2641
rect 17497 2632 17509 2635
rect 17184 2604 17509 2632
rect 17184 2592 17190 2604
rect 17497 2601 17509 2604
rect 17543 2601 17555 2635
rect 17497 2595 17555 2601
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 20714 2632 20720 2644
rect 20211 2604 20720 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 21082 2592 21088 2644
rect 21140 2632 21146 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21140 2604 21833 2632
rect 21140 2592 21146 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 21821 2595 21879 2601
rect 24394 2592 24400 2644
rect 24452 2592 24458 2644
rect 25317 2635 25375 2641
rect 25317 2601 25329 2635
rect 25363 2632 25375 2635
rect 25406 2632 25412 2644
rect 25363 2604 25412 2632
rect 25363 2601 25375 2604
rect 25317 2595 25375 2601
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 27433 2635 27491 2641
rect 27433 2601 27445 2635
rect 27479 2632 27491 2635
rect 27614 2632 27620 2644
rect 27479 2604 27620 2632
rect 27479 2601 27491 2604
rect 27433 2595 27491 2601
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 29089 2635 29147 2641
rect 29089 2601 29101 2635
rect 29135 2632 29147 2635
rect 29362 2632 29368 2644
rect 29135 2604 29368 2632
rect 29135 2601 29147 2604
rect 29089 2595 29147 2601
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 29733 2635 29791 2641
rect 29733 2601 29745 2635
rect 29779 2632 29791 2635
rect 30374 2632 30380 2644
rect 29779 2604 30380 2632
rect 29779 2601 29791 2604
rect 29733 2595 29791 2601
rect 30374 2592 30380 2604
rect 30432 2592 30438 2644
rect 30469 2635 30527 2641
rect 30469 2601 30481 2635
rect 30515 2632 30527 2635
rect 30926 2632 30932 2644
rect 30515 2604 30932 2632
rect 30515 2601 30527 2604
rect 30469 2595 30527 2601
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 33134 2592 33140 2644
rect 33192 2632 33198 2644
rect 33965 2635 34023 2641
rect 33965 2632 33977 2635
rect 33192 2604 33977 2632
rect 33192 2592 33198 2604
rect 33965 2601 33977 2604
rect 34011 2601 34023 2635
rect 36078 2632 36084 2644
rect 33965 2595 34023 2601
rect 34164 2604 36084 2632
rect 10244 2564 10272 2592
rect 4019 2536 6316 2564
rect 4019 2533 4031 2536
rect 3973 2527 4031 2533
rect 1854 2456 1860 2508
rect 1912 2456 1918 2508
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2464 2468 2789 2496
rect 2464 2456 2470 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 2004 2400 2053 2428
rect 2004 2388 2010 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2130 2388 2136 2440
rect 2188 2388 2194 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4798 2428 4804 2440
rect 4203 2400 4804 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 3804 2292 3832 2391
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 5258 2320 5264 2372
rect 5316 2320 5322 2372
rect 5994 2292 6000 2304
rect 3804 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 6288 2292 6316 2536
rect 6380 2536 6776 2564
rect 6886 2536 10272 2564
rect 14277 2567 14335 2573
rect 6380 2437 6408 2536
rect 6748 2496 6776 2536
rect 14277 2533 14289 2567
rect 14323 2564 14335 2567
rect 16040 2564 16068 2592
rect 14323 2536 16068 2564
rect 19429 2567 19487 2573
rect 14323 2533 14335 2536
rect 14277 2527 14335 2533
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 23474 2564 23480 2576
rect 19475 2536 23480 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 27522 2524 27528 2576
rect 27580 2524 27586 2576
rect 32309 2567 32367 2573
rect 32309 2533 32321 2567
rect 32355 2564 32367 2567
rect 34164 2564 34192 2604
rect 36078 2592 36084 2604
rect 36136 2592 36142 2644
rect 36814 2592 36820 2644
rect 36872 2632 36878 2644
rect 37093 2635 37151 2641
rect 37093 2632 37105 2635
rect 36872 2604 37105 2632
rect 36872 2592 36878 2604
rect 37093 2601 37105 2604
rect 37139 2601 37151 2635
rect 37093 2595 37151 2601
rect 38562 2592 38568 2644
rect 38620 2592 38626 2644
rect 39206 2592 39212 2644
rect 39264 2632 39270 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 39264 2604 39405 2632
rect 39264 2592 39270 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 39669 2635 39727 2641
rect 39669 2601 39681 2635
rect 39715 2632 39727 2635
rect 40126 2632 40132 2644
rect 39715 2604 40132 2632
rect 39715 2601 39727 2604
rect 39669 2595 39727 2601
rect 40126 2592 40132 2604
rect 40184 2592 40190 2644
rect 40494 2592 40500 2644
rect 40552 2632 40558 2644
rect 41325 2635 41383 2641
rect 41325 2632 41337 2635
rect 40552 2604 41337 2632
rect 40552 2592 40558 2604
rect 41325 2601 41337 2604
rect 41371 2601 41383 2635
rect 41325 2595 41383 2601
rect 41506 2592 41512 2644
rect 41564 2632 41570 2644
rect 42061 2635 42119 2641
rect 42061 2632 42073 2635
rect 41564 2604 42073 2632
rect 41564 2592 41570 2604
rect 42061 2601 42073 2604
rect 42107 2601 42119 2635
rect 42061 2595 42119 2601
rect 43806 2592 43812 2644
rect 43864 2632 43870 2644
rect 43901 2635 43959 2641
rect 43901 2632 43913 2635
rect 43864 2604 43913 2632
rect 43864 2592 43870 2604
rect 43901 2601 43913 2604
rect 43947 2601 43959 2635
rect 43901 2595 43959 2601
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 45005 2635 45063 2641
rect 45005 2632 45017 2635
rect 44232 2604 45017 2632
rect 44232 2592 44238 2604
rect 45005 2601 45017 2604
rect 45051 2601 45063 2635
rect 45005 2595 45063 2601
rect 47210 2592 47216 2644
rect 47268 2592 47274 2644
rect 49786 2592 49792 2644
rect 49844 2592 49850 2644
rect 50154 2592 50160 2644
rect 50212 2592 50218 2644
rect 51166 2592 51172 2644
rect 51224 2592 51230 2644
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 52181 2635 52239 2641
rect 52181 2632 52193 2635
rect 52052 2604 52193 2632
rect 52052 2592 52058 2604
rect 52181 2601 52193 2604
rect 52227 2601 52239 2635
rect 52181 2595 52239 2601
rect 53374 2592 53380 2644
rect 53432 2592 53438 2644
rect 55122 2592 55128 2644
rect 55180 2592 55186 2644
rect 56594 2592 56600 2644
rect 56652 2592 56658 2644
rect 56778 2592 56784 2644
rect 56836 2632 56842 2644
rect 57241 2635 57299 2641
rect 57241 2632 57253 2635
rect 56836 2604 57253 2632
rect 56836 2592 56842 2604
rect 57241 2601 57253 2604
rect 57287 2601 57299 2635
rect 57241 2595 57299 2601
rect 57422 2592 57428 2644
rect 57480 2632 57486 2644
rect 57885 2635 57943 2641
rect 57885 2632 57897 2635
rect 57480 2604 57897 2632
rect 57480 2592 57486 2604
rect 57885 2601 57897 2604
rect 57931 2601 57943 2635
rect 57885 2595 57943 2601
rect 35618 2564 35624 2576
rect 32355 2536 34192 2564
rect 34256 2536 35624 2564
rect 32355 2533 32367 2536
rect 32309 2527 32367 2533
rect 8386 2496 8392 2508
rect 6748 2468 8392 2496
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9824 2468 10333 2496
rect 9824 2456 9830 2468
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 13449 2499 13507 2505
rect 13449 2465 13461 2499
rect 13495 2496 13507 2499
rect 14182 2496 14188 2508
rect 13495 2468 14188 2496
rect 13495 2465 13507 2468
rect 13449 2459 13507 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 15286 2456 15292 2508
rect 15344 2456 15350 2508
rect 15838 2456 15844 2508
rect 15896 2456 15902 2508
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 17920 2468 18061 2496
rect 17920 2456 17926 2468
rect 18049 2465 18061 2468
rect 18095 2465 18107 2499
rect 18049 2459 18107 2465
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20036 2468 20300 2496
rect 20036 2456 20042 2468
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7006 2428 7012 2440
rect 6779 2400 7012 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 8662 2388 8668 2440
rect 8720 2388 8726 2440
rect 9214 2388 9220 2440
rect 9272 2388 9278 2440
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 12216 2400 12265 2428
rect 12216 2388 12222 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 13596 2400 13737 2428
rect 13596 2388 13602 2400
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15304 2428 15332 2456
rect 15243 2400 15332 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 7558 2320 7564 2372
rect 7616 2320 7622 2372
rect 11054 2292 11060 2304
rect 6288 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 14108 2292 14136 2391
rect 15028 2360 15056 2391
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19426 2428 19432 2440
rect 19291 2400 19432 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 20070 2428 20076 2440
rect 19659 2400 20076 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20272 2437 20300 2468
rect 20806 2456 20812 2508
rect 20864 2456 20870 2508
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 22462 2496 22468 2508
rect 21876 2468 22468 2496
rect 21876 2456 21882 2468
rect 22462 2456 22468 2468
rect 22520 2496 22526 2508
rect 22520 2468 22600 2496
rect 22520 2456 22526 2468
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 22186 2388 22192 2440
rect 22244 2428 22250 2440
rect 22572 2437 22600 2468
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22796 2468 23029 2496
rect 22796 2456 22802 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 25866 2456 25872 2508
rect 25924 2456 25930 2508
rect 27540 2496 27568 2524
rect 27080 2468 27568 2496
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22244 2400 22385 2428
rect 22244 2388 22250 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 25222 2428 25228 2440
rect 24811 2400 25228 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 27080 2437 27108 2468
rect 27706 2456 27712 2508
rect 27764 2496 27770 2508
rect 27985 2499 28043 2505
rect 27985 2496 27997 2499
rect 27764 2468 27997 2496
rect 27764 2456 27770 2468
rect 27985 2465 27997 2468
rect 28031 2465 28043 2499
rect 27985 2459 28043 2465
rect 31018 2456 31024 2508
rect 31076 2456 31082 2508
rect 31110 2456 31116 2508
rect 31168 2496 31174 2508
rect 34256 2496 34284 2536
rect 35618 2524 35624 2536
rect 35676 2524 35682 2576
rect 36357 2567 36415 2573
rect 36357 2533 36369 2567
rect 36403 2564 36415 2567
rect 38580 2564 38608 2592
rect 36403 2536 38608 2564
rect 44637 2567 44695 2573
rect 36403 2533 36415 2536
rect 36357 2527 36415 2533
rect 44637 2533 44649 2567
rect 44683 2564 44695 2567
rect 44726 2564 44732 2576
rect 44683 2536 44732 2564
rect 44683 2533 44695 2536
rect 44637 2527 44695 2533
rect 44726 2524 44732 2536
rect 44784 2524 44790 2576
rect 49697 2567 49755 2573
rect 49697 2533 49709 2567
rect 49743 2533 49755 2567
rect 49697 2527 49755 2533
rect 31168 2468 34284 2496
rect 31168 2456 31174 2468
rect 27060 2431 27118 2437
rect 27060 2397 27072 2431
rect 27106 2397 27118 2431
rect 27060 2391 27118 2397
rect 27246 2388 27252 2440
rect 27304 2388 27310 2440
rect 27338 2388 27344 2440
rect 27396 2388 27402 2440
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 27525 2431 27583 2437
rect 27525 2397 27537 2431
rect 27571 2397 27583 2431
rect 27525 2391 27583 2397
rect 15286 2360 15292 2372
rect 15028 2332 15292 2360
rect 15286 2320 15292 2332
rect 15344 2320 15350 2372
rect 27157 2363 27215 2369
rect 27157 2329 27169 2363
rect 27203 2360 27215 2363
rect 27356 2360 27384 2388
rect 27540 2360 27568 2391
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 29273 2431 29331 2437
rect 29273 2428 29285 2431
rect 29144 2400 29285 2428
rect 29144 2388 29150 2400
rect 29273 2397 29285 2400
rect 29319 2397 29331 2431
rect 29273 2391 29331 2397
rect 29546 2388 29552 2440
rect 29604 2388 29610 2440
rect 29917 2431 29975 2437
rect 29917 2397 29929 2431
rect 29963 2428 29975 2431
rect 30190 2428 30196 2440
rect 29963 2400 30196 2428
rect 29963 2397 29975 2400
rect 29917 2391 29975 2397
rect 30190 2388 30196 2400
rect 30248 2388 30254 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30834 2428 30840 2440
rect 30791 2400 30840 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 33686 2388 33692 2440
rect 33744 2428 33750 2440
rect 34149 2431 34207 2437
rect 33744 2400 34100 2428
rect 33744 2388 33750 2400
rect 27203 2332 27568 2360
rect 27203 2329 27215 2332
rect 27157 2323 27215 2329
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 32677 2363 32735 2369
rect 32677 2360 32689 2363
rect 32456 2332 32689 2360
rect 32456 2320 32462 2332
rect 32677 2329 32689 2332
rect 32723 2329 32735 2363
rect 32677 2323 32735 2329
rect 33962 2320 33968 2372
rect 34020 2320 34026 2372
rect 34072 2360 34100 2400
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34256 2428 34284 2468
rect 35066 2456 35072 2508
rect 35124 2456 35130 2508
rect 35802 2456 35808 2508
rect 35860 2496 35866 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 35860 2468 37749 2496
rect 35860 2456 35866 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 38654 2456 38660 2508
rect 38712 2496 38718 2508
rect 38712 2468 38884 2496
rect 38712 2456 38718 2468
rect 34195 2400 34284 2428
rect 34369 2431 34427 2437
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34369 2397 34381 2431
rect 34415 2428 34427 2431
rect 35084 2428 35112 2456
rect 34415 2400 35112 2428
rect 34415 2397 34427 2400
rect 34369 2391 34427 2397
rect 35894 2388 35900 2440
rect 35952 2388 35958 2440
rect 36170 2388 36176 2440
rect 36228 2388 36234 2440
rect 36541 2431 36599 2437
rect 36541 2397 36553 2431
rect 36587 2428 36599 2431
rect 36814 2428 36820 2440
rect 36587 2400 36820 2428
rect 36587 2397 36599 2400
rect 36541 2391 36599 2397
rect 36814 2388 36820 2400
rect 36872 2388 36878 2440
rect 36906 2388 36912 2440
rect 36964 2428 36970 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36964 2400 37289 2428
rect 36964 2388 36970 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 38746 2388 38752 2440
rect 38804 2388 38810 2440
rect 38856 2428 38884 2468
rect 39022 2456 39028 2508
rect 39080 2496 39086 2508
rect 40313 2499 40371 2505
rect 40313 2496 40325 2499
rect 39080 2468 40325 2496
rect 39080 2456 39086 2468
rect 40313 2465 40325 2468
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 42610 2456 42616 2508
rect 42668 2496 42674 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42668 2468 42901 2496
rect 42668 2456 42674 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 45554 2456 45560 2508
rect 45612 2456 45618 2508
rect 47670 2456 47676 2508
rect 47728 2496 47734 2508
rect 48041 2499 48099 2505
rect 48041 2496 48053 2499
rect 47728 2468 48053 2496
rect 47728 2456 47734 2468
rect 48041 2465 48053 2468
rect 48087 2465 48099 2499
rect 49712 2496 49740 2527
rect 51184 2496 51212 2592
rect 53392 2564 53420 2592
rect 55401 2567 55459 2573
rect 55401 2564 55413 2567
rect 53392 2536 55413 2564
rect 55401 2533 55413 2536
rect 55447 2533 55459 2567
rect 56612 2564 56640 2592
rect 57517 2567 57575 2573
rect 57517 2564 57529 2567
rect 56612 2536 57529 2564
rect 55401 2527 55459 2533
rect 57517 2533 57529 2536
rect 57563 2533 57575 2567
rect 57517 2527 57575 2533
rect 49712 2468 50384 2496
rect 51184 2468 52408 2496
rect 48041 2459 48099 2465
rect 39485 2431 39543 2437
rect 39485 2428 39497 2431
rect 38856 2400 39497 2428
rect 39485 2397 39497 2400
rect 39531 2397 39543 2431
rect 39485 2391 39543 2397
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 39942 2388 39948 2440
rect 40000 2388 40006 2440
rect 40126 2388 40132 2440
rect 40184 2428 40190 2440
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 40184 2400 41889 2428
rect 40184 2388 40190 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 42242 2388 42248 2440
rect 42300 2388 42306 2440
rect 42334 2388 42340 2440
rect 42392 2428 42398 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 42392 2400 42441 2428
rect 42392 2388 42398 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 44453 2431 44511 2437
rect 44453 2428 44465 2431
rect 43220 2400 44465 2428
rect 43220 2388 43226 2400
rect 44453 2397 44465 2400
rect 44499 2397 44511 2431
rect 44453 2391 44511 2397
rect 44818 2388 44824 2440
rect 44876 2388 44882 2440
rect 46566 2388 46572 2440
rect 46624 2428 46630 2440
rect 46937 2431 46995 2437
rect 46937 2428 46949 2431
rect 46624 2400 46949 2428
rect 46624 2388 46630 2400
rect 46937 2397 46949 2400
rect 46983 2397 46995 2431
rect 46937 2391 46995 2397
rect 47397 2431 47455 2437
rect 47397 2397 47409 2431
rect 47443 2397 47455 2431
rect 47397 2391 47455 2397
rect 47765 2431 47823 2437
rect 47765 2397 47777 2431
rect 47811 2428 47823 2431
rect 47946 2428 47952 2440
rect 47811 2400 47952 2428
rect 47811 2397 47823 2400
rect 47765 2391 47823 2397
rect 34241 2363 34299 2369
rect 34241 2360 34253 2363
rect 34072 2332 34253 2360
rect 34241 2329 34253 2332
rect 34287 2329 34299 2363
rect 34241 2323 34299 2329
rect 34514 2320 34520 2372
rect 34572 2360 34578 2372
rect 34885 2363 34943 2369
rect 34885 2360 34897 2363
rect 34572 2332 34897 2360
rect 34572 2320 34578 2332
rect 34885 2329 34897 2332
rect 34931 2329 34943 2363
rect 34885 2323 34943 2329
rect 45646 2320 45652 2372
rect 45704 2360 45710 2372
rect 45925 2363 45983 2369
rect 45925 2360 45937 2363
rect 45704 2332 45937 2360
rect 45704 2320 45710 2332
rect 45925 2329 45937 2332
rect 45971 2329 45983 2363
rect 47412 2360 47440 2391
rect 47946 2388 47952 2400
rect 48004 2388 48010 2440
rect 48406 2388 48412 2440
rect 48464 2428 48470 2440
rect 49053 2431 49111 2437
rect 49053 2428 49065 2431
rect 48464 2400 49065 2428
rect 48464 2388 48470 2400
rect 49053 2397 49065 2400
rect 49099 2397 49111 2431
rect 49053 2391 49111 2397
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 50356 2437 50384 2468
rect 49973 2431 50031 2437
rect 49973 2428 49985 2431
rect 49752 2400 49985 2428
rect 49752 2388 49758 2400
rect 49973 2397 49985 2400
rect 50019 2397 50031 2431
rect 49973 2391 50031 2397
rect 50341 2431 50399 2437
rect 50341 2397 50353 2431
rect 50387 2397 50399 2431
rect 50341 2391 50399 2397
rect 52086 2388 52092 2440
rect 52144 2388 52150 2440
rect 52380 2437 52408 2468
rect 52454 2456 52460 2508
rect 52512 2496 52518 2508
rect 53193 2499 53251 2505
rect 53193 2496 53205 2499
rect 52512 2468 53205 2496
rect 52512 2456 52518 2468
rect 53193 2465 53205 2468
rect 53239 2465 53251 2499
rect 53193 2459 53251 2465
rect 54864 2468 55214 2496
rect 52365 2431 52423 2437
rect 52365 2397 52377 2431
rect 52411 2397 52423 2431
rect 52365 2391 52423 2397
rect 52546 2388 52552 2440
rect 52604 2428 52610 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52604 2400 52745 2428
rect 52604 2388 52610 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53374 2388 53380 2440
rect 53432 2428 53438 2440
rect 54864 2437 54892 2468
rect 54205 2431 54263 2437
rect 54205 2428 54217 2431
rect 53432 2400 54217 2428
rect 53432 2388 53438 2400
rect 54205 2397 54217 2400
rect 54251 2397 54263 2431
rect 54205 2391 54263 2397
rect 54849 2431 54907 2437
rect 54849 2397 54861 2431
rect 54895 2397 54907 2431
rect 54849 2391 54907 2397
rect 54941 2431 54999 2437
rect 54941 2397 54953 2431
rect 54987 2397 54999 2431
rect 55186 2428 55214 2468
rect 56778 2456 56784 2508
rect 56836 2496 56842 2508
rect 56836 2468 58480 2496
rect 56836 2456 56842 2468
rect 55585 2431 55643 2437
rect 55585 2428 55597 2431
rect 55186 2400 55597 2428
rect 54941 2391 54999 2397
rect 55585 2397 55597 2400
rect 55631 2397 55643 2431
rect 55585 2391 55643 2397
rect 47854 2360 47860 2372
rect 47412 2332 47860 2360
rect 45925 2323 45983 2329
rect 47854 2320 47860 2332
rect 47912 2320 47918 2372
rect 50798 2320 50804 2372
rect 50856 2360 50862 2372
rect 51077 2363 51135 2369
rect 51077 2360 51089 2363
rect 50856 2332 51089 2360
rect 50856 2320 50862 2332
rect 51077 2329 51089 2332
rect 51123 2329 51135 2363
rect 51077 2323 51135 2329
rect 52914 2320 52920 2372
rect 52972 2360 52978 2372
rect 54956 2360 54984 2391
rect 56870 2388 56876 2440
rect 56928 2388 56934 2440
rect 56962 2388 56968 2440
rect 57020 2428 57026 2440
rect 58452 2437 58480 2468
rect 57425 2431 57483 2437
rect 57425 2428 57437 2431
rect 57020 2400 57437 2428
rect 57020 2388 57026 2400
rect 57425 2397 57437 2400
rect 57471 2397 57483 2431
rect 57425 2391 57483 2397
rect 57701 2431 57759 2437
rect 57701 2397 57713 2431
rect 57747 2397 57759 2431
rect 57701 2391 57759 2397
rect 58437 2431 58495 2437
rect 58437 2397 58449 2431
rect 58483 2397 58495 2431
rect 58437 2391 58495 2397
rect 52972 2332 54984 2360
rect 52972 2320 52978 2332
rect 55674 2320 55680 2372
rect 55732 2360 55738 2372
rect 55861 2363 55919 2369
rect 55861 2360 55873 2363
rect 55732 2332 55873 2360
rect 55732 2320 55738 2332
rect 55861 2329 55873 2332
rect 55907 2329 55919 2363
rect 55861 2323 55919 2329
rect 56318 2320 56324 2372
rect 56376 2360 56382 2372
rect 57716 2360 57744 2391
rect 56376 2332 57744 2360
rect 56376 2320 56382 2332
rect 15194 2292 15200 2304
rect 14108 2264 15200 2292
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 1104 2202 59040 2224
rect 1104 2150 15394 2202
rect 15446 2150 15458 2202
rect 15510 2150 15522 2202
rect 15574 2150 15586 2202
rect 15638 2150 15650 2202
rect 15702 2150 29838 2202
rect 29890 2150 29902 2202
rect 29954 2150 29966 2202
rect 30018 2150 30030 2202
rect 30082 2150 30094 2202
rect 30146 2150 44282 2202
rect 44334 2150 44346 2202
rect 44398 2150 44410 2202
rect 44462 2150 44474 2202
rect 44526 2150 44538 2202
rect 44590 2150 58726 2202
rect 58778 2150 58790 2202
rect 58842 2150 58854 2202
rect 58906 2150 58918 2202
rect 58970 2150 58982 2202
rect 59034 2150 59040 2202
rect 1104 2128 59040 2150
rect 26326 2048 26332 2100
rect 26384 2088 26390 2100
rect 26970 2088 26976 2100
rect 26384 2060 26976 2088
rect 26384 2048 26390 2060
rect 26970 2048 26976 2060
rect 27028 2048 27034 2100
<< via1 >>
rect 8172 27718 8224 27770
rect 8236 27718 8288 27770
rect 8300 27718 8352 27770
rect 8364 27718 8416 27770
rect 8428 27718 8480 27770
rect 22616 27718 22668 27770
rect 22680 27718 22732 27770
rect 22744 27718 22796 27770
rect 22808 27718 22860 27770
rect 22872 27718 22924 27770
rect 37060 27718 37112 27770
rect 37124 27718 37176 27770
rect 37188 27718 37240 27770
rect 37252 27718 37304 27770
rect 37316 27718 37368 27770
rect 51504 27718 51556 27770
rect 51568 27718 51620 27770
rect 51632 27718 51684 27770
rect 51696 27718 51748 27770
rect 51760 27718 51812 27770
rect 51356 27412 51408 27464
rect 51908 27276 51960 27328
rect 15394 27174 15446 27226
rect 15458 27174 15510 27226
rect 15522 27174 15574 27226
rect 15586 27174 15638 27226
rect 15650 27174 15702 27226
rect 29838 27174 29890 27226
rect 29902 27174 29954 27226
rect 29966 27174 30018 27226
rect 30030 27174 30082 27226
rect 30094 27174 30146 27226
rect 44282 27174 44334 27226
rect 44346 27174 44398 27226
rect 44410 27174 44462 27226
rect 44474 27174 44526 27226
rect 44538 27174 44590 27226
rect 58726 27174 58778 27226
rect 58790 27174 58842 27226
rect 58854 27174 58906 27226
rect 58918 27174 58970 27226
rect 58982 27174 59034 27226
rect 30380 27004 30432 27056
rect 17316 26868 17368 26920
rect 28356 26911 28408 26920
rect 28356 26877 28365 26911
rect 28365 26877 28399 26911
rect 28399 26877 28408 26911
rect 28356 26868 28408 26877
rect 28724 26911 28776 26920
rect 28724 26877 28733 26911
rect 28733 26877 28767 26911
rect 28767 26877 28776 26911
rect 28724 26868 28776 26877
rect 30196 26868 30248 26920
rect 30288 26868 30340 26920
rect 45192 26911 45244 26920
rect 45192 26877 45201 26911
rect 45201 26877 45235 26911
rect 45235 26877 45244 26911
rect 45192 26868 45244 26877
rect 46296 26868 46348 26920
rect 46664 26911 46716 26920
rect 46664 26877 46673 26911
rect 46673 26877 46707 26911
rect 46707 26877 46716 26911
rect 46664 26868 46716 26877
rect 48136 26911 48188 26920
rect 48136 26877 48145 26911
rect 48145 26877 48179 26911
rect 48179 26877 48188 26911
rect 48136 26868 48188 26877
rect 49240 26911 49292 26920
rect 49240 26877 49249 26911
rect 49249 26877 49283 26911
rect 49283 26877 49292 26911
rect 49240 26868 49292 26877
rect 50804 26911 50856 26920
rect 50804 26877 50813 26911
rect 50813 26877 50847 26911
rect 50847 26877 50856 26911
rect 50804 26868 50856 26877
rect 51080 26911 51132 26920
rect 51080 26877 51089 26911
rect 51089 26877 51123 26911
rect 51123 26877 51132 26911
rect 51080 26868 51132 26877
rect 52000 26868 52052 26920
rect 54668 26911 54720 26920
rect 54668 26877 54677 26911
rect 54677 26877 54711 26911
rect 54711 26877 54720 26911
rect 54668 26868 54720 26877
rect 45468 26800 45520 26852
rect 48228 26800 48280 26852
rect 18696 26732 18748 26784
rect 18972 26732 19024 26784
rect 27804 26775 27856 26784
rect 27804 26741 27813 26775
rect 27813 26741 27847 26775
rect 27847 26741 27856 26775
rect 27804 26732 27856 26741
rect 30104 26732 30156 26784
rect 31208 26775 31260 26784
rect 31208 26741 31217 26775
rect 31217 26741 31251 26775
rect 31251 26741 31260 26775
rect 31208 26732 31260 26741
rect 45836 26775 45888 26784
rect 45836 26741 45845 26775
rect 45845 26741 45879 26775
rect 45879 26741 45888 26775
rect 45836 26732 45888 26741
rect 47308 26775 47360 26784
rect 47308 26741 47317 26775
rect 47317 26741 47351 26775
rect 47351 26741 47360 26775
rect 47308 26732 47360 26741
rect 47584 26775 47636 26784
rect 47584 26741 47593 26775
rect 47593 26741 47627 26775
rect 47627 26741 47636 26775
rect 47584 26732 47636 26741
rect 48780 26732 48832 26784
rect 50252 26775 50304 26784
rect 50252 26741 50261 26775
rect 50261 26741 50295 26775
rect 50295 26741 50304 26775
rect 50252 26732 50304 26741
rect 50712 26732 50764 26784
rect 52092 26732 52144 26784
rect 53840 26732 53892 26784
rect 8172 26630 8224 26682
rect 8236 26630 8288 26682
rect 8300 26630 8352 26682
rect 8364 26630 8416 26682
rect 8428 26630 8480 26682
rect 22616 26630 22668 26682
rect 22680 26630 22732 26682
rect 22744 26630 22796 26682
rect 22808 26630 22860 26682
rect 22872 26630 22924 26682
rect 37060 26630 37112 26682
rect 37124 26630 37176 26682
rect 37188 26630 37240 26682
rect 37252 26630 37304 26682
rect 37316 26630 37368 26682
rect 51504 26630 51556 26682
rect 51568 26630 51620 26682
rect 51632 26630 51684 26682
rect 51696 26630 51748 26682
rect 51760 26630 51812 26682
rect 17316 26571 17368 26580
rect 17316 26537 17325 26571
rect 17325 26537 17359 26571
rect 17359 26537 17368 26571
rect 17316 26528 17368 26537
rect 48136 26528 48188 26580
rect 51356 26528 51408 26580
rect 48780 26460 48832 26512
rect 54668 26460 54720 26512
rect 15108 26188 15160 26240
rect 15844 26256 15896 26308
rect 17868 26256 17920 26308
rect 19800 26367 19852 26376
rect 19800 26333 19809 26367
rect 19809 26333 19843 26367
rect 19843 26333 19852 26367
rect 19800 26324 19852 26333
rect 22468 26256 22520 26308
rect 16764 26231 16816 26240
rect 16764 26197 16773 26231
rect 16773 26197 16807 26231
rect 16807 26197 16816 26231
rect 16764 26188 16816 26197
rect 17316 26188 17368 26240
rect 27620 26188 27672 26240
rect 29644 26324 29696 26376
rect 30104 26367 30156 26376
rect 30104 26333 30138 26367
rect 30138 26333 30156 26367
rect 30104 26324 30156 26333
rect 46572 26324 46624 26376
rect 47308 26324 47360 26376
rect 48228 26324 48280 26376
rect 49884 26324 49936 26376
rect 28448 26256 28500 26308
rect 44180 26256 44232 26308
rect 29276 26231 29328 26240
rect 29276 26197 29285 26231
rect 29285 26197 29319 26231
rect 29319 26197 29328 26231
rect 29276 26188 29328 26197
rect 30840 26188 30892 26240
rect 31576 26188 31628 26240
rect 45376 26256 45428 26308
rect 48136 26256 48188 26308
rect 50712 26256 50764 26308
rect 54208 26367 54260 26376
rect 54208 26333 54217 26367
rect 54217 26333 54251 26367
rect 54251 26333 54260 26367
rect 54208 26324 54260 26333
rect 54392 26367 54444 26376
rect 54392 26333 54401 26367
rect 54401 26333 54435 26367
rect 54435 26333 54444 26367
rect 54392 26324 54444 26333
rect 45744 26188 45796 26240
rect 46388 26231 46440 26240
rect 46388 26197 46397 26231
rect 46397 26197 46431 26231
rect 46431 26197 46440 26231
rect 46388 26188 46440 26197
rect 46848 26188 46900 26240
rect 48596 26188 48648 26240
rect 51356 26188 51408 26240
rect 52368 26188 52420 26240
rect 54576 26188 54628 26240
rect 15394 26086 15446 26138
rect 15458 26086 15510 26138
rect 15522 26086 15574 26138
rect 15586 26086 15638 26138
rect 15650 26086 15702 26138
rect 29838 26086 29890 26138
rect 29902 26086 29954 26138
rect 29966 26086 30018 26138
rect 30030 26086 30082 26138
rect 30094 26086 30146 26138
rect 44282 26086 44334 26138
rect 44346 26086 44398 26138
rect 44410 26086 44462 26138
rect 44474 26086 44526 26138
rect 44538 26086 44590 26138
rect 58726 26086 58778 26138
rect 58790 26086 58842 26138
rect 58854 26086 58906 26138
rect 58918 26086 58970 26138
rect 58982 26086 59034 26138
rect 16488 25984 16540 26036
rect 19800 25984 19852 26036
rect 28908 25984 28960 26036
rect 29644 25984 29696 26036
rect 29828 25984 29880 26036
rect 45192 25984 45244 26036
rect 45836 25984 45888 26036
rect 46296 25984 46348 26036
rect 46664 25984 46716 26036
rect 46848 26027 46900 26036
rect 46848 25993 46857 26027
rect 46857 25993 46891 26027
rect 46891 25993 46900 26027
rect 46848 25984 46900 25993
rect 47584 25984 47636 26036
rect 49240 25984 49292 26036
rect 51080 25984 51132 26036
rect 52000 26027 52052 26036
rect 52000 25993 52009 26027
rect 52009 25993 52043 26027
rect 52043 25993 52052 26027
rect 52000 25984 52052 25993
rect 27804 25959 27856 25968
rect 15108 25848 15160 25900
rect 27804 25925 27838 25959
rect 27838 25925 27856 25959
rect 27804 25916 27856 25925
rect 45468 25916 45520 25968
rect 27620 25848 27672 25900
rect 29920 25891 29972 25900
rect 29920 25857 29929 25891
rect 29929 25857 29963 25891
rect 29963 25857 29972 25891
rect 29920 25848 29972 25857
rect 30012 25848 30064 25900
rect 46572 25916 46624 25968
rect 7012 25823 7064 25832
rect 7012 25789 7021 25823
rect 7021 25789 7055 25823
rect 7055 25789 7064 25823
rect 7012 25780 7064 25789
rect 7748 25823 7800 25832
rect 7748 25789 7757 25823
rect 7757 25789 7791 25823
rect 7791 25789 7800 25823
rect 7748 25780 7800 25789
rect 8024 25780 8076 25832
rect 10968 25823 11020 25832
rect 10968 25789 10977 25823
rect 10977 25789 11011 25823
rect 11011 25789 11020 25823
rect 10968 25780 11020 25789
rect 13820 25823 13872 25832
rect 13820 25789 13829 25823
rect 13829 25789 13863 25823
rect 13863 25789 13872 25823
rect 13820 25780 13872 25789
rect 14372 25823 14424 25832
rect 14372 25789 14381 25823
rect 14381 25789 14415 25823
rect 14415 25789 14424 25823
rect 14372 25780 14424 25789
rect 17316 25823 17368 25832
rect 17316 25789 17325 25823
rect 17325 25789 17359 25823
rect 17359 25789 17368 25823
rect 17316 25780 17368 25789
rect 17408 25780 17460 25832
rect 17592 25823 17644 25832
rect 17592 25789 17601 25823
rect 17601 25789 17635 25823
rect 17635 25789 17644 25823
rect 17592 25780 17644 25789
rect 12440 25712 12492 25764
rect 6460 25687 6512 25696
rect 6460 25653 6469 25687
rect 6469 25653 6503 25687
rect 6503 25653 6512 25687
rect 6460 25644 6512 25653
rect 7196 25687 7248 25696
rect 7196 25653 7205 25687
rect 7205 25653 7239 25687
rect 7239 25653 7248 25687
rect 7196 25644 7248 25653
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 7932 25644 7984 25653
rect 8852 25687 8904 25696
rect 8852 25653 8861 25687
rect 8861 25653 8895 25687
rect 8895 25653 8904 25687
rect 8852 25644 8904 25653
rect 10416 25687 10468 25696
rect 10416 25653 10425 25687
rect 10425 25653 10459 25687
rect 10459 25653 10468 25687
rect 10416 25644 10468 25653
rect 13176 25712 13228 25764
rect 17868 25755 17920 25764
rect 17868 25721 17877 25755
rect 17877 25721 17911 25755
rect 17911 25721 17920 25755
rect 17868 25712 17920 25721
rect 18696 25780 18748 25832
rect 19248 25780 19300 25832
rect 18972 25712 19024 25764
rect 28724 25780 28776 25832
rect 29552 25780 29604 25832
rect 30840 25780 30892 25832
rect 31300 25823 31352 25832
rect 31300 25789 31309 25823
rect 31309 25789 31343 25823
rect 31343 25789 31352 25823
rect 31300 25780 31352 25789
rect 31576 25712 31628 25764
rect 45652 25848 45704 25900
rect 46848 25848 46900 25900
rect 48136 25848 48188 25900
rect 48596 25848 48648 25900
rect 50252 25916 50304 25968
rect 49884 25848 49936 25900
rect 50896 25848 50948 25900
rect 51908 25848 51960 25900
rect 52276 25848 52328 25900
rect 53840 25916 53892 25968
rect 54484 25984 54536 26036
rect 54392 25916 54444 25968
rect 45744 25823 45796 25832
rect 45744 25789 45753 25823
rect 45753 25789 45787 25823
rect 45787 25789 45796 25823
rect 45744 25780 45796 25789
rect 46664 25780 46716 25832
rect 12900 25644 12952 25696
rect 16580 25644 16632 25696
rect 17500 25644 17552 25696
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 20444 25687 20496 25696
rect 20444 25653 20453 25687
rect 20453 25653 20487 25687
rect 20487 25653 20496 25687
rect 20444 25644 20496 25653
rect 30656 25644 30708 25696
rect 31668 25644 31720 25696
rect 32128 25687 32180 25696
rect 32128 25653 32137 25687
rect 32137 25653 32171 25687
rect 32171 25653 32180 25687
rect 32128 25644 32180 25653
rect 46020 25644 46072 25696
rect 51264 25780 51316 25832
rect 51356 25823 51408 25832
rect 51356 25789 51365 25823
rect 51365 25789 51399 25823
rect 51399 25789 51408 25823
rect 51356 25780 51408 25789
rect 52000 25780 52052 25832
rect 54576 25891 54628 25900
rect 54576 25857 54585 25891
rect 54585 25857 54619 25891
rect 54619 25857 54628 25891
rect 54576 25848 54628 25857
rect 52368 25712 52420 25764
rect 48780 25644 48832 25696
rect 8172 25542 8224 25594
rect 8236 25542 8288 25594
rect 8300 25542 8352 25594
rect 8364 25542 8416 25594
rect 8428 25542 8480 25594
rect 22616 25542 22668 25594
rect 22680 25542 22732 25594
rect 22744 25542 22796 25594
rect 22808 25542 22860 25594
rect 22872 25542 22924 25594
rect 37060 25542 37112 25594
rect 37124 25542 37176 25594
rect 37188 25542 37240 25594
rect 37252 25542 37304 25594
rect 37316 25542 37368 25594
rect 51504 25542 51556 25594
rect 51568 25542 51620 25594
rect 51632 25542 51684 25594
rect 51696 25542 51748 25594
rect 51760 25542 51812 25594
rect 7748 25483 7800 25492
rect 7748 25449 7757 25483
rect 7757 25449 7791 25483
rect 7791 25449 7800 25483
rect 7748 25440 7800 25449
rect 8024 25440 8076 25492
rect 10968 25440 11020 25492
rect 14280 25440 14332 25492
rect 14372 25440 14424 25492
rect 8024 25304 8076 25356
rect 8852 25304 8904 25356
rect 17960 25440 18012 25492
rect 19248 25483 19300 25492
rect 19248 25449 19257 25483
rect 19257 25449 19291 25483
rect 19291 25449 19300 25483
rect 19248 25440 19300 25449
rect 28356 25440 28408 25492
rect 5540 25279 5592 25288
rect 5540 25245 5549 25279
rect 5549 25245 5583 25279
rect 5583 25245 5592 25279
rect 5540 25236 5592 25245
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 6460 25236 6512 25288
rect 9496 25279 9548 25288
rect 9496 25245 9505 25279
rect 9505 25245 9539 25279
rect 9539 25245 9548 25279
rect 9496 25236 9548 25245
rect 11428 25279 11480 25288
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 12440 25236 12492 25288
rect 12900 25236 12952 25288
rect 8576 25168 8628 25220
rect 15752 25347 15804 25356
rect 15752 25313 15761 25347
rect 15761 25313 15795 25347
rect 15795 25313 15804 25347
rect 15752 25304 15804 25313
rect 16488 25347 16540 25356
rect 16120 25236 16172 25288
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 16764 25304 16816 25356
rect 17592 25372 17644 25424
rect 27712 25415 27764 25424
rect 27712 25381 27721 25415
rect 27721 25381 27755 25415
rect 27755 25381 27764 25415
rect 27712 25372 27764 25381
rect 29000 25372 29052 25424
rect 29920 25440 29972 25492
rect 30380 25440 30432 25492
rect 31668 25483 31720 25492
rect 31668 25449 31677 25483
rect 31677 25449 31711 25483
rect 31711 25449 31720 25483
rect 31668 25440 31720 25449
rect 45836 25440 45888 25492
rect 46848 25440 46900 25492
rect 46940 25440 46992 25492
rect 49884 25483 49936 25492
rect 49884 25449 49893 25483
rect 49893 25449 49927 25483
rect 49927 25449 49936 25483
rect 49884 25440 49936 25449
rect 50804 25440 50856 25492
rect 50896 25440 50948 25492
rect 18788 25236 18840 25288
rect 26240 25279 26292 25288
rect 26240 25245 26249 25279
rect 26249 25245 26283 25279
rect 26283 25245 26292 25279
rect 26240 25236 26292 25245
rect 4896 25143 4948 25152
rect 4896 25109 4905 25143
rect 4905 25109 4939 25143
rect 4939 25109 4948 25143
rect 4896 25100 4948 25109
rect 7104 25100 7156 25152
rect 11704 25100 11756 25152
rect 17408 25168 17460 25220
rect 18236 25168 18288 25220
rect 38384 25304 38436 25356
rect 44916 25304 44968 25356
rect 46020 25372 46072 25424
rect 45928 25304 45980 25356
rect 47584 25304 47636 25356
rect 48228 25304 48280 25356
rect 30196 25236 30248 25288
rect 32128 25236 32180 25288
rect 29552 25168 29604 25220
rect 46756 25279 46808 25288
rect 46756 25245 46765 25279
rect 46765 25245 46799 25279
rect 46799 25245 46808 25279
rect 46756 25236 46808 25245
rect 46848 25236 46900 25288
rect 12624 25100 12676 25152
rect 13912 25100 13964 25152
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 16028 25143 16080 25152
rect 16028 25109 16037 25143
rect 16037 25109 16071 25143
rect 16071 25109 16080 25143
rect 16028 25100 16080 25109
rect 25136 25143 25188 25152
rect 25136 25109 25145 25143
rect 25145 25109 25179 25143
rect 25179 25109 25188 25143
rect 25136 25100 25188 25109
rect 25596 25143 25648 25152
rect 25596 25109 25605 25143
rect 25605 25109 25639 25143
rect 25639 25109 25648 25143
rect 25596 25100 25648 25109
rect 27252 25143 27304 25152
rect 27252 25109 27261 25143
rect 27261 25109 27295 25143
rect 27295 25109 27304 25143
rect 27252 25100 27304 25109
rect 29092 25143 29144 25152
rect 29092 25109 29101 25143
rect 29101 25109 29135 25143
rect 29135 25109 29144 25143
rect 29092 25100 29144 25109
rect 45652 25168 45704 25220
rect 45008 25143 45060 25152
rect 45008 25109 45017 25143
rect 45017 25109 45051 25143
rect 45051 25109 45060 25143
rect 45008 25100 45060 25109
rect 48044 25100 48096 25152
rect 52092 25304 52144 25356
rect 52276 25347 52328 25356
rect 52276 25313 52285 25347
rect 52285 25313 52319 25347
rect 52319 25313 52328 25347
rect 52276 25304 52328 25313
rect 52552 25347 52604 25356
rect 52552 25313 52561 25347
rect 52561 25313 52595 25347
rect 52595 25313 52604 25347
rect 52552 25304 52604 25313
rect 52000 25279 52052 25288
rect 52000 25245 52009 25279
rect 52009 25245 52043 25279
rect 52043 25245 52052 25279
rect 52000 25236 52052 25245
rect 54208 25440 54260 25492
rect 54576 25372 54628 25424
rect 53380 25347 53432 25356
rect 53380 25313 53389 25347
rect 53389 25313 53423 25347
rect 53423 25313 53432 25347
rect 53380 25304 53432 25313
rect 54668 25347 54720 25356
rect 54668 25313 54677 25347
rect 54677 25313 54711 25347
rect 54711 25313 54720 25347
rect 54668 25304 54720 25313
rect 48780 25100 48832 25152
rect 50804 25143 50856 25152
rect 50804 25109 50813 25143
rect 50813 25109 50847 25143
rect 50847 25109 50856 25143
rect 50804 25100 50856 25109
rect 53196 25100 53248 25152
rect 15394 24998 15446 25050
rect 15458 24998 15510 25050
rect 15522 24998 15574 25050
rect 15586 24998 15638 25050
rect 15650 24998 15702 25050
rect 29838 24998 29890 25050
rect 29902 24998 29954 25050
rect 29966 24998 30018 25050
rect 30030 24998 30082 25050
rect 30094 24998 30146 25050
rect 44282 24998 44334 25050
rect 44346 24998 44398 25050
rect 44410 24998 44462 25050
rect 44474 24998 44526 25050
rect 44538 24998 44590 25050
rect 58726 24998 58778 25050
rect 58790 24998 58842 25050
rect 58854 24998 58906 25050
rect 58918 24998 58970 25050
rect 58982 24998 59034 25050
rect 4896 24828 4948 24880
rect 7012 24896 7064 24948
rect 7104 24939 7156 24948
rect 7104 24905 7113 24939
rect 7113 24905 7147 24939
rect 7147 24905 7156 24939
rect 7104 24896 7156 24905
rect 7196 24939 7248 24948
rect 7196 24905 7205 24939
rect 7205 24905 7239 24939
rect 7239 24905 7248 24939
rect 7196 24896 7248 24905
rect 9496 24896 9548 24948
rect 11428 24896 11480 24948
rect 5908 24760 5960 24812
rect 7932 24828 7984 24880
rect 10416 24828 10468 24880
rect 13820 24939 13872 24948
rect 13820 24905 13829 24939
rect 13829 24905 13863 24939
rect 13863 24905 13872 24939
rect 13820 24896 13872 24905
rect 14740 24896 14792 24948
rect 17408 24896 17460 24948
rect 18236 24939 18288 24948
rect 18236 24905 18245 24939
rect 18245 24905 18279 24939
rect 18279 24905 18288 24939
rect 18236 24896 18288 24905
rect 29552 24896 29604 24948
rect 30840 24896 30892 24948
rect 3976 24556 4028 24608
rect 6368 24624 6420 24676
rect 8668 24692 8720 24744
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 12532 24735 12584 24744
rect 12532 24701 12541 24735
rect 12541 24701 12575 24735
rect 12575 24701 12584 24735
rect 12532 24692 12584 24701
rect 12624 24692 12676 24744
rect 6184 24599 6236 24608
rect 6184 24565 6193 24599
rect 6193 24565 6227 24599
rect 6227 24565 6236 24599
rect 6184 24556 6236 24565
rect 11244 24556 11296 24608
rect 11888 24599 11940 24608
rect 11888 24565 11897 24599
rect 11897 24565 11931 24599
rect 11931 24565 11940 24599
rect 11888 24556 11940 24565
rect 12348 24556 12400 24608
rect 13176 24624 13228 24676
rect 17868 24828 17920 24880
rect 19800 24828 19852 24880
rect 13544 24735 13596 24744
rect 13544 24701 13553 24735
rect 13553 24701 13587 24735
rect 13587 24701 13596 24735
rect 13544 24692 13596 24701
rect 13636 24692 13688 24744
rect 14280 24760 14332 24812
rect 15752 24760 15804 24812
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 16028 24760 16080 24812
rect 16580 24760 16632 24812
rect 18604 24760 18656 24812
rect 19340 24760 19392 24812
rect 25320 24760 25372 24812
rect 27712 24828 27764 24880
rect 29092 24828 29144 24880
rect 29736 24828 29788 24880
rect 20812 24692 20864 24744
rect 24216 24735 24268 24744
rect 24216 24701 24225 24735
rect 24225 24701 24259 24735
rect 24259 24701 24268 24735
rect 24216 24692 24268 24701
rect 26516 24803 26568 24812
rect 26516 24769 26525 24803
rect 26525 24769 26559 24803
rect 26559 24769 26568 24803
rect 26516 24760 26568 24769
rect 27620 24760 27672 24812
rect 28448 24803 28500 24812
rect 28448 24769 28457 24803
rect 28457 24769 28491 24803
rect 28491 24769 28500 24803
rect 28448 24760 28500 24769
rect 29000 24803 29052 24812
rect 29000 24769 29009 24803
rect 29009 24769 29043 24803
rect 29043 24769 29052 24803
rect 29000 24760 29052 24769
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29276 24760 29328 24769
rect 42708 24760 42760 24812
rect 27988 24692 28040 24744
rect 30840 24735 30892 24744
rect 30840 24701 30849 24735
rect 30849 24701 30883 24735
rect 30883 24701 30892 24735
rect 42892 24803 42944 24812
rect 42892 24769 42901 24803
rect 42901 24769 42935 24803
rect 42935 24769 42944 24803
rect 42892 24760 42944 24769
rect 45928 24939 45980 24948
rect 45928 24905 45937 24939
rect 45937 24905 45971 24939
rect 45971 24905 45980 24939
rect 45928 24896 45980 24905
rect 51172 24896 51224 24948
rect 52000 24896 52052 24948
rect 52552 24896 52604 24948
rect 45008 24760 45060 24812
rect 45376 24760 45428 24812
rect 46388 24760 46440 24812
rect 30840 24692 30892 24701
rect 16212 24624 16264 24676
rect 25228 24624 25280 24676
rect 26240 24556 26292 24608
rect 30288 24556 30340 24608
rect 42248 24599 42300 24608
rect 42248 24565 42257 24599
rect 42257 24565 42291 24599
rect 42291 24565 42300 24599
rect 44640 24735 44692 24744
rect 44640 24701 44649 24735
rect 44649 24701 44683 24735
rect 44683 24701 44692 24735
rect 44640 24692 44692 24701
rect 42708 24624 42760 24676
rect 50620 24760 50672 24812
rect 52552 24803 52604 24812
rect 52552 24769 52561 24803
rect 52561 24769 52595 24803
rect 52595 24769 52604 24803
rect 52552 24760 52604 24769
rect 46664 24624 46716 24676
rect 53380 24896 53432 24948
rect 42248 24556 42300 24565
rect 42800 24556 42852 24608
rect 42984 24556 43036 24608
rect 47492 24556 47544 24608
rect 51264 24599 51316 24608
rect 51264 24565 51273 24599
rect 51273 24565 51307 24599
rect 51307 24565 51316 24599
rect 51264 24556 51316 24565
rect 8172 24454 8224 24506
rect 8236 24454 8288 24506
rect 8300 24454 8352 24506
rect 8364 24454 8416 24506
rect 8428 24454 8480 24506
rect 22616 24454 22668 24506
rect 22680 24454 22732 24506
rect 22744 24454 22796 24506
rect 22808 24454 22860 24506
rect 22872 24454 22924 24506
rect 37060 24454 37112 24506
rect 37124 24454 37176 24506
rect 37188 24454 37240 24506
rect 37252 24454 37304 24506
rect 37316 24454 37368 24506
rect 51504 24454 51556 24506
rect 51568 24454 51620 24506
rect 51632 24454 51684 24506
rect 51696 24454 51748 24506
rect 51760 24454 51812 24506
rect 5540 24352 5592 24404
rect 6184 24352 6236 24404
rect 7196 24352 7248 24404
rect 3976 24259 4028 24268
rect 3976 24225 3985 24259
rect 3985 24225 4019 24259
rect 4019 24225 4028 24259
rect 3976 24216 4028 24225
rect 5908 24259 5960 24268
rect 5908 24225 5917 24259
rect 5917 24225 5951 24259
rect 5951 24225 5960 24259
rect 5908 24216 5960 24225
rect 6092 24259 6144 24268
rect 6092 24225 6101 24259
rect 6101 24225 6135 24259
rect 6135 24225 6144 24259
rect 6092 24216 6144 24225
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 6920 24191 6972 24200
rect 6920 24157 6929 24191
rect 6929 24157 6963 24191
rect 6963 24157 6972 24191
rect 6920 24148 6972 24157
rect 7012 24148 7064 24200
rect 11888 24352 11940 24404
rect 13544 24352 13596 24404
rect 26516 24395 26568 24404
rect 26516 24361 26525 24395
rect 26525 24361 26559 24395
rect 26559 24361 26568 24395
rect 26516 24352 26568 24361
rect 42708 24352 42760 24404
rect 42800 24352 42852 24404
rect 8576 24216 8628 24268
rect 11244 24216 11296 24268
rect 9864 24148 9916 24200
rect 12440 24148 12492 24200
rect 44640 24352 44692 24404
rect 46664 24352 46716 24404
rect 24860 24216 24912 24268
rect 13084 24148 13136 24200
rect 13728 24148 13780 24200
rect 13820 24148 13872 24200
rect 14096 24148 14148 24200
rect 4528 24080 4580 24132
rect 10692 24080 10744 24132
rect 12348 24080 12400 24132
rect 12624 24080 12676 24132
rect 20168 24191 20220 24200
rect 20168 24157 20177 24191
rect 20177 24157 20211 24191
rect 20211 24157 20220 24191
rect 20168 24148 20220 24157
rect 20812 24148 20864 24200
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 22192 24148 22244 24200
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 24952 24148 25004 24200
rect 25136 24148 25188 24200
rect 26056 24148 26108 24200
rect 27068 24191 27120 24200
rect 27068 24157 27077 24191
rect 27077 24157 27111 24191
rect 27111 24157 27120 24191
rect 27068 24148 27120 24157
rect 33508 24191 33560 24200
rect 33508 24157 33517 24191
rect 33517 24157 33551 24191
rect 33551 24157 33560 24191
rect 33508 24148 33560 24157
rect 33692 24191 33744 24200
rect 33692 24157 33701 24191
rect 33701 24157 33735 24191
rect 33735 24157 33744 24191
rect 33692 24148 33744 24157
rect 35992 24191 36044 24200
rect 35992 24157 36001 24191
rect 36001 24157 36035 24191
rect 36035 24157 36044 24191
rect 35992 24148 36044 24157
rect 37556 24191 37608 24200
rect 37556 24157 37565 24191
rect 37565 24157 37599 24191
rect 37599 24157 37608 24191
rect 37556 24148 37608 24157
rect 37740 24191 37792 24200
rect 37740 24157 37749 24191
rect 37749 24157 37783 24191
rect 37783 24157 37792 24191
rect 37740 24148 37792 24157
rect 40408 24191 40460 24200
rect 40408 24157 40417 24191
rect 40417 24157 40451 24191
rect 40451 24157 40460 24191
rect 40408 24148 40460 24157
rect 41144 24191 41196 24200
rect 41144 24157 41153 24191
rect 41153 24157 41187 24191
rect 41187 24157 41196 24191
rect 41144 24148 41196 24157
rect 42340 24191 42392 24200
rect 42340 24157 42349 24191
rect 42349 24157 42383 24191
rect 42383 24157 42392 24191
rect 42340 24148 42392 24157
rect 42524 24148 42576 24200
rect 42984 24148 43036 24200
rect 43996 24191 44048 24200
rect 43996 24157 44005 24191
rect 44005 24157 44039 24191
rect 44039 24157 44048 24191
rect 43996 24148 44048 24157
rect 46480 24191 46532 24200
rect 46480 24157 46489 24191
rect 46489 24157 46523 24191
rect 46523 24157 46532 24191
rect 46480 24148 46532 24157
rect 46756 24191 46808 24200
rect 46756 24157 46765 24191
rect 46765 24157 46799 24191
rect 46799 24157 46808 24191
rect 46756 24148 46808 24157
rect 48136 24191 48188 24200
rect 48136 24157 48145 24191
rect 48145 24157 48179 24191
rect 48179 24157 48188 24191
rect 48136 24148 48188 24157
rect 50988 24191 51040 24200
rect 50988 24157 50997 24191
rect 50997 24157 51031 24191
rect 51031 24157 51040 24191
rect 50988 24148 51040 24157
rect 51908 24191 51960 24200
rect 51908 24157 51917 24191
rect 51917 24157 51951 24191
rect 51951 24157 51960 24191
rect 51908 24148 51960 24157
rect 52644 24191 52696 24200
rect 52644 24157 52653 24191
rect 52653 24157 52687 24191
rect 52687 24157 52696 24191
rect 52644 24148 52696 24157
rect 53288 24191 53340 24200
rect 53288 24157 53297 24191
rect 53297 24157 53331 24191
rect 53331 24157 53340 24191
rect 53288 24148 53340 24157
rect 54392 24191 54444 24200
rect 54392 24157 54401 24191
rect 54401 24157 54435 24191
rect 54435 24157 54444 24191
rect 54392 24148 54444 24157
rect 55312 24191 55364 24200
rect 55312 24157 55321 24191
rect 55321 24157 55355 24191
rect 55355 24157 55364 24191
rect 55312 24148 55364 24157
rect 56876 24148 56928 24200
rect 57244 24148 57296 24200
rect 20260 24080 20312 24132
rect 23296 24080 23348 24132
rect 27528 24080 27580 24132
rect 5356 24055 5408 24064
rect 5356 24021 5365 24055
rect 5365 24021 5399 24055
rect 5399 24021 5408 24055
rect 5356 24012 5408 24021
rect 7564 24012 7616 24064
rect 7656 24012 7708 24064
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 11428 24055 11480 24064
rect 11428 24021 11437 24055
rect 11437 24021 11471 24055
rect 11471 24021 11480 24055
rect 11428 24012 11480 24021
rect 11704 24012 11756 24064
rect 13636 24012 13688 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 21272 24012 21324 24064
rect 21456 24012 21508 24064
rect 22100 24055 22152 24064
rect 22100 24021 22109 24055
rect 22109 24021 22143 24055
rect 22143 24021 22152 24055
rect 22100 24012 22152 24021
rect 23388 24055 23440 24064
rect 23388 24021 23397 24055
rect 23397 24021 23431 24055
rect 23431 24021 23440 24055
rect 23388 24012 23440 24021
rect 25044 24012 25096 24064
rect 26516 24012 26568 24064
rect 27804 24012 27856 24064
rect 32956 24055 33008 24064
rect 32956 24021 32965 24055
rect 32965 24021 32999 24055
rect 32999 24021 33008 24055
rect 32956 24012 33008 24021
rect 34336 24055 34388 24064
rect 34336 24021 34345 24055
rect 34345 24021 34379 24055
rect 34379 24021 34388 24055
rect 34336 24012 34388 24021
rect 35440 24055 35492 24064
rect 35440 24021 35449 24055
rect 35449 24021 35483 24055
rect 35483 24021 35492 24055
rect 35440 24012 35492 24021
rect 36820 24012 36872 24064
rect 38936 24012 38988 24064
rect 39672 24055 39724 24064
rect 39672 24021 39681 24055
rect 39681 24021 39715 24055
rect 39715 24021 39724 24055
rect 39672 24012 39724 24021
rect 39856 24055 39908 24064
rect 39856 24021 39865 24055
rect 39865 24021 39899 24055
rect 39899 24021 39908 24055
rect 39856 24012 39908 24021
rect 40592 24055 40644 24064
rect 40592 24021 40601 24055
rect 40601 24021 40635 24055
rect 40635 24021 40644 24055
rect 40592 24012 40644 24021
rect 41696 24055 41748 24064
rect 41696 24021 41705 24055
rect 41705 24021 41739 24055
rect 41739 24021 41748 24055
rect 41696 24012 41748 24021
rect 44640 24055 44692 24064
rect 44640 24021 44649 24055
rect 44649 24021 44683 24055
rect 44683 24021 44692 24055
rect 44640 24012 44692 24021
rect 45928 24055 45980 24064
rect 45928 24021 45937 24055
rect 45937 24021 45971 24055
rect 45971 24021 45980 24055
rect 45928 24012 45980 24021
rect 47400 24012 47452 24064
rect 48320 24012 48372 24064
rect 50436 24055 50488 24064
rect 50436 24021 50445 24055
rect 50445 24021 50479 24055
rect 50479 24021 50488 24055
rect 50436 24012 50488 24021
rect 51356 24012 51408 24064
rect 52460 24012 52512 24064
rect 52736 24055 52788 24064
rect 52736 24021 52745 24055
rect 52745 24021 52779 24055
rect 52779 24021 52788 24055
rect 52736 24012 52788 24021
rect 53656 24055 53708 24064
rect 53656 24021 53665 24055
rect 53665 24021 53699 24055
rect 53699 24021 53708 24055
rect 53656 24012 53708 24021
rect 53840 24055 53892 24064
rect 53840 24021 53849 24055
rect 53849 24021 53883 24055
rect 53883 24021 53892 24055
rect 53840 24012 53892 24021
rect 54576 24012 54628 24064
rect 55220 24012 55272 24064
rect 56048 24012 56100 24064
rect 56600 24055 56652 24064
rect 56600 24021 56609 24055
rect 56609 24021 56643 24055
rect 56643 24021 56652 24055
rect 56600 24012 56652 24021
rect 57336 24055 57388 24064
rect 57336 24021 57345 24055
rect 57345 24021 57379 24055
rect 57379 24021 57388 24055
rect 57336 24012 57388 24021
rect 15394 23910 15446 23962
rect 15458 23910 15510 23962
rect 15522 23910 15574 23962
rect 15586 23910 15638 23962
rect 15650 23910 15702 23962
rect 29838 23910 29890 23962
rect 29902 23910 29954 23962
rect 29966 23910 30018 23962
rect 30030 23910 30082 23962
rect 30094 23910 30146 23962
rect 44282 23910 44334 23962
rect 44346 23910 44398 23962
rect 44410 23910 44462 23962
rect 44474 23910 44526 23962
rect 44538 23910 44590 23962
rect 58726 23910 58778 23962
rect 58790 23910 58842 23962
rect 58854 23910 58906 23962
rect 58918 23910 58970 23962
rect 58982 23910 59034 23962
rect 5540 23808 5592 23860
rect 5908 23808 5960 23860
rect 5356 23740 5408 23792
rect 5356 23647 5408 23656
rect 5356 23613 5365 23647
rect 5365 23613 5399 23647
rect 5399 23613 5408 23647
rect 5356 23604 5408 23613
rect 7012 23808 7064 23860
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 11428 23808 11480 23860
rect 13544 23808 13596 23860
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 17960 23808 18012 23860
rect 19340 23808 19392 23860
rect 19432 23808 19484 23860
rect 20168 23851 20220 23860
rect 20168 23817 20177 23851
rect 20177 23817 20211 23851
rect 20211 23817 20220 23851
rect 20168 23808 20220 23817
rect 20260 23851 20312 23860
rect 20260 23817 20269 23851
rect 20269 23817 20303 23851
rect 20303 23817 20312 23851
rect 20260 23808 20312 23817
rect 23296 23808 23348 23860
rect 23940 23808 23992 23860
rect 4712 23511 4764 23520
rect 4712 23477 4721 23511
rect 4721 23477 4755 23511
rect 4755 23477 4764 23511
rect 4712 23468 4764 23477
rect 6092 23468 6144 23520
rect 11244 23740 11296 23792
rect 14188 23740 14240 23792
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 13268 23604 13320 23656
rect 18696 23672 18748 23724
rect 21272 23672 21324 23724
rect 22100 23740 22152 23792
rect 25228 23808 25280 23860
rect 27068 23808 27120 23860
rect 27528 23808 27580 23860
rect 31300 23808 31352 23860
rect 31576 23851 31628 23860
rect 31576 23817 31585 23851
rect 31585 23817 31619 23851
rect 31619 23817 31628 23851
rect 31576 23808 31628 23817
rect 24860 23740 24912 23792
rect 15200 23604 15252 23656
rect 16396 23647 16448 23656
rect 16396 23613 16405 23647
rect 16405 23613 16439 23647
rect 16439 23613 16448 23647
rect 16396 23604 16448 23613
rect 17408 23647 17460 23656
rect 17408 23613 17417 23647
rect 17417 23613 17451 23647
rect 17451 23613 17460 23647
rect 17408 23604 17460 23613
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 7012 23468 7064 23520
rect 12624 23468 12676 23520
rect 13728 23468 13780 23520
rect 14832 23511 14884 23520
rect 14832 23477 14841 23511
rect 14841 23477 14875 23511
rect 14875 23477 14884 23511
rect 14832 23468 14884 23477
rect 15844 23511 15896 23520
rect 15844 23477 15853 23511
rect 15853 23477 15887 23511
rect 15887 23477 15896 23511
rect 15844 23468 15896 23477
rect 16212 23468 16264 23520
rect 16856 23511 16908 23520
rect 16856 23477 16865 23511
rect 16865 23477 16899 23511
rect 16899 23477 16908 23511
rect 16856 23468 16908 23477
rect 19892 23536 19944 23588
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 20444 23468 20496 23520
rect 20812 23468 20864 23520
rect 21364 23468 21416 23520
rect 22008 23536 22060 23588
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 25320 23740 25372 23792
rect 25872 23740 25924 23792
rect 29736 23740 29788 23792
rect 30380 23740 30432 23792
rect 33140 23808 33192 23860
rect 33692 23808 33744 23860
rect 34152 23808 34204 23860
rect 37556 23808 37608 23860
rect 38936 23808 38988 23860
rect 39856 23808 39908 23860
rect 41144 23808 41196 23860
rect 45652 23808 45704 23860
rect 46480 23808 46532 23860
rect 48136 23808 48188 23860
rect 50988 23808 51040 23860
rect 53288 23808 53340 23860
rect 54392 23808 54444 23860
rect 32036 23672 32088 23724
rect 32956 23672 33008 23724
rect 25044 23604 25096 23656
rect 27712 23604 27764 23656
rect 29184 23604 29236 23656
rect 35440 23740 35492 23792
rect 35532 23672 35584 23724
rect 23112 23468 23164 23520
rect 24860 23468 24912 23520
rect 27252 23468 27304 23520
rect 28080 23468 28132 23520
rect 30472 23468 30524 23520
rect 30748 23468 30800 23520
rect 31576 23468 31628 23520
rect 34060 23468 34112 23520
rect 37648 23604 37700 23656
rect 38292 23715 38344 23724
rect 38292 23681 38301 23715
rect 38301 23681 38335 23715
rect 38335 23681 38344 23715
rect 38292 23672 38344 23681
rect 38384 23672 38436 23724
rect 38568 23672 38620 23724
rect 42708 23740 42760 23792
rect 42892 23740 42944 23792
rect 40224 23715 40276 23724
rect 40224 23681 40233 23715
rect 40233 23681 40267 23715
rect 40267 23681 40276 23715
rect 40224 23672 40276 23681
rect 40316 23715 40368 23724
rect 40316 23681 40325 23715
rect 40325 23681 40359 23715
rect 40359 23681 40368 23715
rect 40316 23672 40368 23681
rect 34520 23468 34572 23520
rect 35716 23511 35768 23520
rect 35716 23477 35725 23511
rect 35725 23477 35759 23511
rect 35759 23477 35768 23511
rect 35716 23468 35768 23477
rect 35900 23468 35952 23520
rect 39672 23604 39724 23656
rect 41604 23604 41656 23656
rect 44272 23672 44324 23724
rect 44640 23715 44692 23724
rect 44640 23681 44649 23715
rect 44649 23681 44683 23715
rect 44683 23681 44692 23715
rect 44640 23672 44692 23681
rect 49056 23783 49108 23792
rect 49056 23749 49065 23783
rect 49065 23749 49099 23783
rect 49099 23749 49108 23783
rect 49056 23740 49108 23749
rect 55220 23740 55272 23792
rect 56600 23783 56652 23792
rect 45284 23604 45336 23656
rect 46572 23672 46624 23724
rect 50804 23715 50856 23724
rect 50804 23681 50813 23715
rect 50813 23681 50847 23715
rect 50847 23681 50856 23715
rect 50804 23672 50856 23681
rect 52000 23672 52052 23724
rect 46664 23647 46716 23656
rect 46664 23613 46673 23647
rect 46673 23613 46707 23647
rect 46707 23613 46716 23647
rect 46664 23604 46716 23613
rect 47492 23604 47544 23656
rect 48320 23536 48372 23588
rect 48504 23647 48556 23656
rect 48504 23613 48513 23647
rect 48513 23613 48547 23647
rect 48547 23613 48556 23647
rect 48504 23604 48556 23613
rect 50252 23604 50304 23656
rect 51356 23604 51408 23656
rect 52460 23604 52512 23656
rect 53656 23604 53708 23656
rect 54576 23604 54628 23656
rect 55772 23672 55824 23724
rect 56600 23749 56634 23783
rect 56634 23749 56652 23783
rect 56600 23740 56652 23749
rect 56324 23647 56376 23656
rect 56324 23613 56333 23647
rect 56333 23613 56367 23647
rect 56367 23613 56376 23647
rect 56324 23604 56376 23613
rect 57612 23604 57664 23656
rect 41236 23468 41288 23520
rect 41512 23511 41564 23520
rect 41512 23477 41521 23511
rect 41521 23477 41555 23511
rect 41555 23477 41564 23511
rect 41512 23468 41564 23477
rect 42524 23468 42576 23520
rect 44640 23468 44692 23520
rect 45100 23511 45152 23520
rect 45100 23477 45109 23511
rect 45109 23477 45143 23511
rect 45143 23477 45152 23511
rect 45100 23468 45152 23477
rect 45284 23468 45336 23520
rect 48688 23468 48740 23520
rect 50252 23511 50304 23520
rect 50252 23477 50261 23511
rect 50261 23477 50295 23511
rect 50295 23477 50304 23511
rect 50252 23468 50304 23477
rect 53104 23468 53156 23520
rect 55496 23511 55548 23520
rect 55496 23477 55505 23511
rect 55505 23477 55539 23511
rect 55539 23477 55548 23511
rect 55496 23468 55548 23477
rect 58072 23536 58124 23588
rect 57796 23468 57848 23520
rect 57888 23511 57940 23520
rect 57888 23477 57897 23511
rect 57897 23477 57931 23511
rect 57931 23477 57940 23511
rect 57888 23468 57940 23477
rect 8172 23366 8224 23418
rect 8236 23366 8288 23418
rect 8300 23366 8352 23418
rect 8364 23366 8416 23418
rect 8428 23366 8480 23418
rect 22616 23366 22668 23418
rect 22680 23366 22732 23418
rect 22744 23366 22796 23418
rect 22808 23366 22860 23418
rect 22872 23366 22924 23418
rect 37060 23366 37112 23418
rect 37124 23366 37176 23418
rect 37188 23366 37240 23418
rect 37252 23366 37304 23418
rect 37316 23366 37368 23418
rect 51504 23366 51556 23418
rect 51568 23366 51620 23418
rect 51632 23366 51684 23418
rect 51696 23366 51748 23418
rect 51760 23366 51812 23418
rect 4528 23307 4580 23316
rect 4528 23273 4537 23307
rect 4537 23273 4571 23307
rect 4571 23273 4580 23307
rect 4528 23264 4580 23273
rect 5356 23264 5408 23316
rect 12348 23264 12400 23316
rect 16396 23264 16448 23316
rect 19340 23264 19392 23316
rect 4712 23128 4764 23180
rect 11336 23128 11388 23180
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 13728 23060 13780 23112
rect 15108 23060 15160 23112
rect 18788 23128 18840 23180
rect 19892 23171 19944 23180
rect 19892 23137 19901 23171
rect 19901 23137 19935 23171
rect 19935 23137 19944 23171
rect 19892 23128 19944 23137
rect 22100 23264 22152 23316
rect 24216 23307 24268 23316
rect 24216 23273 24225 23307
rect 24225 23273 24259 23307
rect 24259 23273 24268 23307
rect 24216 23264 24268 23273
rect 26792 23264 26844 23316
rect 27712 23264 27764 23316
rect 33508 23264 33560 23316
rect 21180 23171 21232 23180
rect 21180 23137 21189 23171
rect 21189 23137 21223 23171
rect 21223 23137 21232 23171
rect 21180 23128 21232 23137
rect 21272 23128 21324 23180
rect 14832 22992 14884 23044
rect 16856 22992 16908 23044
rect 8576 22924 8628 22976
rect 12992 22967 13044 22976
rect 12992 22933 13001 22967
rect 13001 22933 13035 22967
rect 13035 22933 13044 22967
rect 12992 22924 13044 22933
rect 13268 22924 13320 22976
rect 17592 22924 17644 22976
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 20168 23060 20220 23112
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 21732 23103 21784 23112
rect 21732 23069 21741 23103
rect 21741 23069 21775 23103
rect 21775 23069 21784 23103
rect 21732 23060 21784 23069
rect 22468 23128 22520 23180
rect 24860 23128 24912 23180
rect 26056 23171 26108 23180
rect 26056 23137 26065 23171
rect 26065 23137 26099 23171
rect 26099 23137 26108 23171
rect 26056 23128 26108 23137
rect 26332 23171 26384 23180
rect 26332 23137 26341 23171
rect 26341 23137 26375 23171
rect 26375 23137 26384 23171
rect 26332 23128 26384 23137
rect 23388 23060 23440 23112
rect 25780 23103 25832 23112
rect 25780 23069 25789 23103
rect 25789 23069 25823 23103
rect 25823 23069 25832 23103
rect 25780 23060 25832 23069
rect 25872 23060 25924 23112
rect 27528 23128 27580 23180
rect 28080 23128 28132 23180
rect 21456 22924 21508 22976
rect 22284 22924 22336 22976
rect 24400 22967 24452 22976
rect 24400 22933 24409 22967
rect 24409 22933 24443 22967
rect 24443 22933 24452 22967
rect 24400 22924 24452 22933
rect 25964 22924 26016 22976
rect 27804 23060 27856 23112
rect 29644 23128 29696 23180
rect 30656 23171 30708 23180
rect 30656 23137 30665 23171
rect 30665 23137 30699 23171
rect 30699 23137 30708 23171
rect 30656 23128 30708 23137
rect 31576 23196 31628 23248
rect 31576 23103 31628 23112
rect 31576 23069 31585 23103
rect 31585 23069 31619 23103
rect 31619 23069 31628 23103
rect 31576 23060 31628 23069
rect 30472 22992 30524 23044
rect 27528 22967 27580 22976
rect 27528 22933 27537 22967
rect 27537 22933 27571 22967
rect 27571 22933 27580 22967
rect 27528 22924 27580 22933
rect 27896 22967 27948 22976
rect 27896 22933 27905 22967
rect 27905 22933 27939 22967
rect 27939 22933 27948 22967
rect 27896 22924 27948 22933
rect 29000 22967 29052 22976
rect 29000 22933 29009 22967
rect 29009 22933 29043 22967
rect 29043 22933 29052 22967
rect 29000 22924 29052 22933
rect 29644 22924 29696 22976
rect 30380 22924 30432 22976
rect 30564 22967 30616 22976
rect 30564 22933 30573 22967
rect 30573 22933 30607 22967
rect 30607 22933 30616 22967
rect 30564 22924 30616 22933
rect 31024 22967 31076 22976
rect 31024 22933 31033 22967
rect 31033 22933 31067 22967
rect 31067 22933 31076 22967
rect 31024 22924 31076 22933
rect 34060 23171 34112 23180
rect 34060 23137 34069 23171
rect 34069 23137 34103 23171
rect 34103 23137 34112 23171
rect 36636 23264 36688 23316
rect 37740 23307 37792 23316
rect 37740 23273 37749 23307
rect 37749 23273 37783 23307
rect 37783 23273 37792 23307
rect 37740 23264 37792 23273
rect 38292 23264 38344 23316
rect 40408 23264 40460 23316
rect 39028 23239 39080 23248
rect 39028 23205 39037 23239
rect 39037 23205 39071 23239
rect 39071 23205 39080 23239
rect 39028 23196 39080 23205
rect 34060 23128 34112 23137
rect 38292 23128 38344 23180
rect 38936 23128 38988 23180
rect 40316 23128 40368 23180
rect 40408 23171 40460 23180
rect 40408 23137 40417 23171
rect 40417 23137 40451 23171
rect 40451 23137 40460 23171
rect 40408 23128 40460 23137
rect 32036 23060 32088 23112
rect 34336 23060 34388 23112
rect 34520 23060 34572 23112
rect 36912 23060 36964 23112
rect 38752 23103 38804 23112
rect 38752 23069 38761 23103
rect 38761 23069 38795 23103
rect 38795 23069 38804 23103
rect 38752 23060 38804 23069
rect 41512 23264 41564 23316
rect 42616 23128 42668 23180
rect 44272 23264 44324 23316
rect 45284 23307 45336 23316
rect 45284 23273 45293 23307
rect 45293 23273 45327 23307
rect 45327 23273 45336 23307
rect 45284 23264 45336 23273
rect 46756 23264 46808 23316
rect 48504 23307 48556 23316
rect 48504 23273 48513 23307
rect 48513 23273 48547 23307
rect 48547 23273 48556 23307
rect 48504 23264 48556 23273
rect 51908 23264 51960 23316
rect 52644 23264 52696 23316
rect 55312 23264 55364 23316
rect 55772 23264 55824 23316
rect 43444 23128 43496 23180
rect 56048 23128 56100 23180
rect 57244 23307 57296 23316
rect 57244 23273 57253 23307
rect 57253 23273 57287 23307
rect 57287 23273 57296 23307
rect 57244 23264 57296 23273
rect 56508 23171 56560 23180
rect 56508 23137 56517 23171
rect 56517 23137 56551 23171
rect 56551 23137 56560 23171
rect 56508 23128 56560 23137
rect 32312 22992 32364 23044
rect 34612 22992 34664 23044
rect 33324 22967 33376 22976
rect 33324 22933 33333 22967
rect 33333 22933 33367 22967
rect 33367 22933 33376 22967
rect 33324 22924 33376 22933
rect 34796 22924 34848 22976
rect 36176 22992 36228 23044
rect 36820 22992 36872 23044
rect 40224 23035 40276 23044
rect 40224 23001 40233 23035
rect 40233 23001 40267 23035
rect 40267 23001 40276 23035
rect 40224 22992 40276 23001
rect 43628 23103 43680 23112
rect 43628 23069 43637 23103
rect 43637 23069 43671 23103
rect 43671 23069 43680 23103
rect 43628 23060 43680 23069
rect 43720 23103 43772 23112
rect 43720 23069 43754 23103
rect 43754 23069 43772 23103
rect 43720 23060 43772 23069
rect 45008 23060 45060 23112
rect 45468 23103 45520 23112
rect 45468 23069 45477 23103
rect 45477 23069 45511 23103
rect 45511 23069 45520 23103
rect 45468 23060 45520 23069
rect 47400 23103 47452 23112
rect 47400 23069 47434 23103
rect 47434 23069 47452 23103
rect 47400 23060 47452 23069
rect 51264 23060 51316 23112
rect 41328 22992 41380 23044
rect 41512 23035 41564 23044
rect 41512 23001 41546 23035
rect 41546 23001 41564 23035
rect 41512 22992 41564 23001
rect 35532 22924 35584 22976
rect 36084 22967 36136 22976
rect 36084 22933 36093 22967
rect 36093 22933 36127 22967
rect 36127 22933 36136 22967
rect 36084 22924 36136 22933
rect 40040 22924 40092 22976
rect 40408 22924 40460 22976
rect 40960 22967 41012 22976
rect 40960 22933 40969 22967
rect 40969 22933 41003 22967
rect 41003 22933 41012 22967
rect 40960 22924 41012 22933
rect 42248 22924 42300 22976
rect 43076 22924 43128 22976
rect 43444 22924 43496 22976
rect 45560 22992 45612 23044
rect 45928 22992 45980 23044
rect 46848 22992 46900 23044
rect 50252 22992 50304 23044
rect 50436 23035 50488 23044
rect 50436 23001 50470 23035
rect 50470 23001 50488 23035
rect 50436 22992 50488 23001
rect 52736 23035 52788 23044
rect 52736 23001 52754 23035
rect 52754 23001 52788 23035
rect 52736 22992 52788 23001
rect 55956 23103 56008 23112
rect 55956 23069 55965 23103
rect 55965 23069 55999 23103
rect 55999 23069 56008 23103
rect 55956 23060 56008 23069
rect 56968 23103 57020 23112
rect 56968 23069 56977 23103
rect 56977 23069 57011 23103
rect 57011 23069 57020 23103
rect 56968 23060 57020 23069
rect 53840 22992 53892 23044
rect 57888 23128 57940 23180
rect 44732 22924 44784 22976
rect 50620 22924 50672 22976
rect 51816 22924 51868 22976
rect 53564 22924 53616 22976
rect 56692 22924 56744 22976
rect 57060 22924 57112 22976
rect 57796 22924 57848 22976
rect 15394 22822 15446 22874
rect 15458 22822 15510 22874
rect 15522 22822 15574 22874
rect 15586 22822 15638 22874
rect 15650 22822 15702 22874
rect 29838 22822 29890 22874
rect 29902 22822 29954 22874
rect 29966 22822 30018 22874
rect 30030 22822 30082 22874
rect 30094 22822 30146 22874
rect 44282 22822 44334 22874
rect 44346 22822 44398 22874
rect 44410 22822 44462 22874
rect 44474 22822 44526 22874
rect 44538 22822 44590 22874
rect 58726 22822 58778 22874
rect 58790 22822 58842 22874
rect 58854 22822 58906 22874
rect 58918 22822 58970 22874
rect 58982 22822 59034 22874
rect 7564 22720 7616 22772
rect 13544 22720 13596 22772
rect 13636 22720 13688 22772
rect 15200 22720 15252 22772
rect 15844 22720 15896 22772
rect 16120 22763 16172 22772
rect 16120 22729 16129 22763
rect 16129 22729 16163 22763
rect 16163 22729 16172 22763
rect 16120 22720 16172 22729
rect 17408 22720 17460 22772
rect 17500 22720 17552 22772
rect 20904 22720 20956 22772
rect 22192 22720 22244 22772
rect 24860 22720 24912 22772
rect 7748 22652 7800 22704
rect 12256 22652 12308 22704
rect 7656 22584 7708 22636
rect 19064 22695 19116 22704
rect 19064 22661 19098 22695
rect 19098 22661 19116 22695
rect 19064 22652 19116 22661
rect 20720 22652 20772 22704
rect 21732 22652 21784 22704
rect 22008 22652 22060 22704
rect 16120 22584 16172 22636
rect 17500 22584 17552 22636
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 20168 22584 20220 22636
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 22468 22584 22520 22636
rect 23112 22584 23164 22636
rect 25044 22652 25096 22704
rect 25596 22720 25648 22772
rect 25964 22763 26016 22772
rect 25964 22729 25973 22763
rect 25973 22729 26007 22763
rect 26007 22729 26016 22763
rect 25964 22720 26016 22729
rect 27436 22720 27488 22772
rect 27896 22720 27948 22772
rect 29184 22763 29236 22772
rect 29184 22729 29193 22763
rect 29193 22729 29227 22763
rect 29227 22729 29236 22763
rect 29184 22720 29236 22729
rect 30564 22720 30616 22772
rect 31576 22720 31628 22772
rect 34796 22720 34848 22772
rect 35716 22763 35768 22772
rect 24400 22584 24452 22636
rect 33140 22652 33192 22704
rect 26424 22584 26476 22636
rect 27528 22584 27580 22636
rect 27620 22584 27672 22636
rect 5908 22559 5960 22568
rect 5908 22525 5917 22559
rect 5917 22525 5951 22559
rect 5951 22525 5960 22559
rect 5908 22516 5960 22525
rect 8576 22516 8628 22568
rect 9404 22559 9456 22568
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 10600 22516 10652 22568
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 11888 22559 11940 22568
rect 11888 22525 11897 22559
rect 11897 22525 11931 22559
rect 11931 22525 11940 22559
rect 11888 22516 11940 22525
rect 5448 22448 5500 22500
rect 7564 22448 7616 22500
rect 9128 22448 9180 22500
rect 13544 22448 13596 22500
rect 13912 22516 13964 22568
rect 14740 22516 14792 22568
rect 15568 22516 15620 22568
rect 17132 22491 17184 22500
rect 17132 22457 17141 22491
rect 17141 22457 17175 22491
rect 17175 22457 17184 22491
rect 18604 22559 18656 22568
rect 18604 22525 18613 22559
rect 18613 22525 18647 22559
rect 18647 22525 18656 22559
rect 18604 22516 18656 22525
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 25780 22559 25832 22568
rect 17132 22448 17184 22457
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 6920 22380 6972 22432
rect 8852 22423 8904 22432
rect 8852 22389 8861 22423
rect 8861 22389 8895 22423
rect 8895 22389 8904 22423
rect 8852 22380 8904 22389
rect 10692 22423 10744 22432
rect 10692 22389 10701 22423
rect 10701 22389 10735 22423
rect 10735 22389 10744 22423
rect 10692 22380 10744 22389
rect 12532 22423 12584 22432
rect 12532 22389 12541 22423
rect 12541 22389 12575 22423
rect 12575 22389 12584 22423
rect 12532 22380 12584 22389
rect 17408 22380 17460 22432
rect 22192 22448 22244 22500
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 29736 22516 29788 22568
rect 30104 22559 30156 22568
rect 30104 22525 30122 22559
rect 30122 22525 30156 22559
rect 30104 22516 30156 22525
rect 30564 22516 30616 22568
rect 24952 22380 25004 22432
rect 29092 22448 29144 22500
rect 30656 22448 30708 22500
rect 27988 22380 28040 22432
rect 30932 22559 30984 22568
rect 30932 22525 30941 22559
rect 30941 22525 30975 22559
rect 30975 22525 30984 22559
rect 30932 22516 30984 22525
rect 33416 22584 33468 22636
rect 31392 22448 31444 22500
rect 32128 22516 32180 22568
rect 33048 22559 33100 22568
rect 33048 22525 33057 22559
rect 33057 22525 33091 22559
rect 33091 22525 33100 22559
rect 33048 22516 33100 22525
rect 34336 22627 34388 22636
rect 34336 22593 34345 22627
rect 34345 22593 34379 22627
rect 34379 22593 34388 22627
rect 34336 22584 34388 22593
rect 35716 22729 35725 22763
rect 35725 22729 35759 22763
rect 35759 22729 35768 22763
rect 35716 22720 35768 22729
rect 36176 22763 36228 22772
rect 36176 22729 36185 22763
rect 36185 22729 36219 22763
rect 36219 22729 36228 22763
rect 36176 22720 36228 22729
rect 41604 22720 41656 22772
rect 42340 22720 42392 22772
rect 42892 22763 42944 22772
rect 42892 22729 42901 22763
rect 42901 22729 42935 22763
rect 42935 22729 42944 22763
rect 42892 22720 42944 22729
rect 43996 22720 44048 22772
rect 35808 22652 35860 22704
rect 34060 22559 34112 22568
rect 34060 22525 34069 22559
rect 34069 22525 34103 22559
rect 34103 22525 34112 22559
rect 34060 22516 34112 22525
rect 34152 22516 34204 22568
rect 34612 22559 34664 22568
rect 34612 22525 34621 22559
rect 34621 22525 34655 22559
rect 34655 22525 34664 22559
rect 34612 22516 34664 22525
rect 35256 22559 35308 22568
rect 35256 22525 35265 22559
rect 35265 22525 35299 22559
rect 35299 22525 35308 22559
rect 35256 22516 35308 22525
rect 38016 22584 38068 22636
rect 38660 22584 38712 22636
rect 40592 22584 40644 22636
rect 41420 22652 41472 22704
rect 42524 22652 42576 22704
rect 43720 22652 43772 22704
rect 44180 22652 44232 22704
rect 45100 22652 45152 22704
rect 45560 22652 45612 22704
rect 48780 22720 48832 22772
rect 50620 22720 50672 22772
rect 52000 22720 52052 22772
rect 53104 22763 53156 22772
rect 53104 22729 53113 22763
rect 53113 22729 53147 22763
rect 53147 22729 53156 22763
rect 53104 22720 53156 22729
rect 53196 22763 53248 22772
rect 53196 22729 53205 22763
rect 53205 22729 53239 22763
rect 53239 22729 53248 22763
rect 53196 22720 53248 22729
rect 55772 22763 55824 22772
rect 55772 22729 55781 22763
rect 55781 22729 55815 22763
rect 55815 22729 55824 22763
rect 55772 22720 55824 22729
rect 57612 22763 57664 22772
rect 57612 22729 57621 22763
rect 57621 22729 57655 22763
rect 57655 22729 57664 22763
rect 57612 22720 57664 22729
rect 53564 22652 53616 22704
rect 41696 22584 41748 22636
rect 44640 22627 44692 22636
rect 44640 22593 44649 22627
rect 44649 22593 44683 22627
rect 44683 22593 44692 22627
rect 44640 22584 44692 22593
rect 45468 22584 45520 22636
rect 46204 22627 46256 22636
rect 46204 22593 46238 22627
rect 46238 22593 46256 22627
rect 46204 22584 46256 22593
rect 46940 22584 46992 22636
rect 48320 22584 48372 22636
rect 49056 22584 49108 22636
rect 36728 22559 36780 22568
rect 36728 22525 36737 22559
rect 36737 22525 36771 22559
rect 36771 22525 36780 22559
rect 36728 22516 36780 22525
rect 36912 22516 36964 22568
rect 43168 22516 43220 22568
rect 44916 22516 44968 22568
rect 34796 22448 34848 22500
rect 35992 22448 36044 22500
rect 32404 22423 32456 22432
rect 32404 22389 32413 22423
rect 32413 22389 32447 22423
rect 32447 22389 32456 22423
rect 32404 22380 32456 22389
rect 35532 22380 35584 22432
rect 38660 22423 38712 22432
rect 38660 22389 38669 22423
rect 38669 22389 38703 22423
rect 38703 22389 38712 22423
rect 38660 22380 38712 22389
rect 42248 22423 42300 22432
rect 42248 22389 42257 22423
rect 42257 22389 42291 22423
rect 42291 22389 42300 22423
rect 42248 22380 42300 22389
rect 42616 22380 42668 22432
rect 45008 22423 45060 22432
rect 45008 22389 45017 22423
rect 45017 22389 45051 22423
rect 45051 22389 45060 22423
rect 45008 22380 45060 22389
rect 47308 22423 47360 22432
rect 47308 22389 47317 22423
rect 47317 22389 47351 22423
rect 47351 22389 47360 22423
rect 47308 22380 47360 22389
rect 47584 22423 47636 22432
rect 47584 22389 47593 22423
rect 47593 22389 47627 22423
rect 47627 22389 47636 22423
rect 47584 22380 47636 22389
rect 48228 22380 48280 22432
rect 49240 22559 49292 22568
rect 49240 22525 49249 22559
rect 49249 22525 49283 22559
rect 49283 22525 49292 22559
rect 49240 22516 49292 22525
rect 51172 22516 51224 22568
rect 51632 22627 51684 22636
rect 51632 22593 51641 22627
rect 51641 22593 51675 22627
rect 51675 22593 51684 22627
rect 51632 22584 51684 22593
rect 52460 22584 52512 22636
rect 55496 22584 55548 22636
rect 57336 22652 57388 22704
rect 56324 22584 56376 22636
rect 58072 22584 58124 22636
rect 51448 22516 51500 22568
rect 52368 22559 52420 22568
rect 52368 22525 52377 22559
rect 52377 22525 52411 22559
rect 52411 22525 52420 22559
rect 52368 22516 52420 22525
rect 52644 22516 52696 22568
rect 48780 22491 48832 22500
rect 48780 22457 48789 22491
rect 48789 22457 48823 22491
rect 48823 22457 48832 22491
rect 48780 22448 48832 22457
rect 49608 22448 49660 22500
rect 51816 22448 51868 22500
rect 51172 22380 51224 22432
rect 52736 22423 52788 22432
rect 52736 22389 52745 22423
rect 52745 22389 52779 22423
rect 52779 22389 52788 22423
rect 52736 22380 52788 22389
rect 56968 22380 57020 22432
rect 8172 22278 8224 22330
rect 8236 22278 8288 22330
rect 8300 22278 8352 22330
rect 8364 22278 8416 22330
rect 8428 22278 8480 22330
rect 22616 22278 22668 22330
rect 22680 22278 22732 22330
rect 22744 22278 22796 22330
rect 22808 22278 22860 22330
rect 22872 22278 22924 22330
rect 37060 22278 37112 22330
rect 37124 22278 37176 22330
rect 37188 22278 37240 22330
rect 37252 22278 37304 22330
rect 37316 22278 37368 22330
rect 51504 22278 51556 22330
rect 51568 22278 51620 22330
rect 51632 22278 51684 22330
rect 51696 22278 51748 22330
rect 51760 22278 51812 22330
rect 5448 22176 5500 22228
rect 5908 22176 5960 22228
rect 9404 22176 9456 22228
rect 11336 22176 11388 22228
rect 11888 22176 11940 22228
rect 12256 22176 12308 22228
rect 6920 22108 6972 22160
rect 7748 22108 7800 22160
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 8852 22040 8904 22092
rect 9680 21972 9732 22024
rect 5172 21947 5224 21956
rect 5172 21913 5181 21947
rect 5181 21913 5215 21947
rect 5215 21913 5224 21947
rect 5172 21904 5224 21913
rect 7196 21904 7248 21956
rect 7472 21904 7524 21956
rect 13912 22219 13964 22228
rect 13912 22185 13921 22219
rect 13921 22185 13955 22219
rect 13955 22185 13964 22219
rect 13912 22176 13964 22185
rect 14740 22176 14792 22228
rect 16396 22176 16448 22228
rect 17132 22176 17184 22228
rect 17592 22176 17644 22228
rect 18604 22176 18656 22228
rect 20168 22219 20220 22228
rect 20168 22185 20177 22219
rect 20177 22185 20211 22219
rect 20211 22185 20220 22219
rect 20168 22176 20220 22185
rect 13636 22040 13688 22092
rect 14740 22083 14792 22092
rect 10324 21972 10376 22024
rect 12440 21972 12492 22024
rect 12808 22015 12860 22024
rect 12808 21981 12842 22015
rect 12842 21981 12860 22015
rect 12808 21972 12860 21981
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 15844 22040 15896 22092
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 4804 21879 4856 21888
rect 4804 21845 4813 21879
rect 4813 21845 4847 21879
rect 4847 21845 4856 21879
rect 4804 21836 4856 21845
rect 5540 21836 5592 21888
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 7288 21836 7340 21888
rect 8300 21836 8352 21888
rect 9404 21879 9456 21888
rect 9404 21845 9413 21879
rect 9413 21845 9447 21879
rect 9447 21845 9456 21879
rect 9404 21836 9456 21845
rect 10692 21904 10744 21956
rect 10600 21836 10652 21888
rect 11060 21836 11112 21888
rect 13728 21904 13780 21956
rect 17132 22083 17184 22092
rect 17132 22049 17141 22083
rect 17141 22049 17175 22083
rect 17175 22049 17184 22083
rect 17132 22040 17184 22049
rect 16580 21972 16632 22024
rect 17224 22015 17276 22024
rect 17224 21981 17258 22015
rect 17258 21981 17276 22015
rect 17224 21972 17276 21981
rect 12532 21836 12584 21888
rect 12992 21836 13044 21888
rect 16304 21836 16356 21888
rect 17316 21836 17368 21888
rect 20628 21904 20680 21956
rect 19800 21836 19852 21888
rect 19892 21836 19944 21888
rect 20444 21836 20496 21888
rect 21180 22176 21232 22228
rect 25780 22176 25832 22228
rect 57060 22176 57112 22228
rect 22468 22040 22520 22092
rect 26332 22108 26384 22160
rect 26976 22108 27028 22160
rect 22192 21972 22244 22024
rect 24860 21836 24912 21888
rect 25044 21836 25096 21888
rect 27804 22083 27856 22092
rect 27804 22049 27813 22083
rect 27813 22049 27847 22083
rect 27847 22049 27856 22083
rect 27804 22040 27856 22049
rect 28908 22040 28960 22092
rect 32128 22151 32180 22160
rect 32128 22117 32137 22151
rect 32137 22117 32171 22151
rect 32171 22117 32180 22151
rect 32128 22108 32180 22117
rect 32312 22151 32364 22160
rect 32312 22117 32321 22151
rect 32321 22117 32355 22151
rect 32355 22117 32364 22151
rect 32312 22108 32364 22117
rect 33416 22108 33468 22160
rect 34152 22108 34204 22160
rect 32404 22040 32456 22092
rect 33048 22040 33100 22092
rect 33324 22040 33376 22092
rect 31024 21972 31076 22024
rect 35256 22108 35308 22160
rect 36636 22108 36688 22160
rect 38016 22151 38068 22160
rect 38016 22117 38025 22151
rect 38025 22117 38059 22151
rect 38059 22117 38068 22151
rect 38016 22108 38068 22117
rect 38752 22151 38804 22160
rect 36084 22083 36136 22092
rect 36084 22049 36093 22083
rect 36093 22049 36127 22083
rect 36127 22049 36136 22083
rect 36084 22040 36136 22049
rect 38752 22117 38761 22151
rect 38761 22117 38795 22151
rect 38795 22117 38804 22151
rect 38752 22108 38804 22117
rect 41512 22151 41564 22160
rect 41512 22117 41521 22151
rect 41521 22117 41555 22151
rect 41555 22117 41564 22151
rect 41512 22108 41564 22117
rect 42616 22108 42668 22160
rect 28264 21904 28316 21956
rect 30840 21904 30892 21956
rect 31300 21904 31352 21956
rect 35808 21972 35860 22024
rect 38660 22040 38712 22092
rect 41328 22040 41380 22092
rect 43628 22108 43680 22160
rect 29276 21836 29328 21888
rect 34060 21879 34112 21888
rect 34060 21845 34069 21879
rect 34069 21845 34103 21879
rect 34103 21845 34112 21879
rect 34060 21836 34112 21845
rect 34888 21836 34940 21888
rect 36728 21836 36780 21888
rect 37648 21836 37700 21888
rect 43076 22083 43128 22092
rect 43076 22049 43085 22083
rect 43085 22049 43119 22083
rect 43119 22049 43128 22083
rect 43076 22040 43128 22049
rect 46388 22083 46440 22092
rect 46388 22049 46397 22083
rect 46397 22049 46431 22083
rect 46431 22049 46440 22083
rect 46388 22040 46440 22049
rect 46848 22040 46900 22092
rect 46940 22015 46992 22024
rect 46940 21981 46949 22015
rect 46949 21981 46983 22015
rect 46983 21981 46992 22015
rect 46940 21972 46992 21981
rect 48044 22083 48096 22092
rect 48044 22049 48053 22083
rect 48053 22049 48087 22083
rect 48087 22049 48096 22083
rect 48044 22040 48096 22049
rect 55956 22108 56008 22160
rect 56508 22108 56560 22160
rect 47584 21972 47636 22024
rect 50160 22015 50212 22024
rect 50160 21981 50169 22015
rect 50169 21981 50203 22015
rect 50203 21981 50212 22015
rect 50160 21972 50212 21981
rect 51356 22040 51408 22092
rect 52644 22083 52696 22092
rect 52644 22049 52653 22083
rect 52653 22049 52687 22083
rect 52687 22049 52696 22083
rect 52644 22040 52696 22049
rect 50988 21904 51040 21956
rect 42892 21836 42944 21888
rect 43168 21836 43220 21888
rect 44640 21836 44692 21888
rect 46480 21879 46532 21888
rect 46480 21845 46489 21879
rect 46489 21845 46523 21879
rect 46523 21845 46532 21879
rect 46480 21836 46532 21845
rect 46664 21836 46716 21888
rect 48320 21836 48372 21888
rect 48964 21836 49016 21888
rect 50068 21836 50120 21888
rect 51080 21836 51132 21888
rect 56048 22040 56100 22092
rect 55220 21836 55272 21888
rect 55864 21836 55916 21888
rect 56968 22015 57020 22024
rect 56968 21981 56977 22015
rect 56977 21981 57011 22015
rect 57011 21981 57020 22015
rect 56968 21972 57020 21981
rect 57796 21972 57848 22024
rect 57980 22015 58032 22024
rect 57980 21981 57989 22015
rect 57989 21981 58023 22015
rect 58023 21981 58032 22015
rect 57980 21972 58032 21981
rect 56876 21836 56928 21888
rect 57428 21879 57480 21888
rect 57428 21845 57437 21879
rect 57437 21845 57471 21879
rect 57471 21845 57480 21879
rect 57428 21836 57480 21845
rect 15394 21734 15446 21786
rect 15458 21734 15510 21786
rect 15522 21734 15574 21786
rect 15586 21734 15638 21786
rect 15650 21734 15702 21786
rect 29838 21734 29890 21786
rect 29902 21734 29954 21786
rect 29966 21734 30018 21786
rect 30030 21734 30082 21786
rect 30094 21734 30146 21786
rect 44282 21734 44334 21786
rect 44346 21734 44398 21786
rect 44410 21734 44462 21786
rect 44474 21734 44526 21786
rect 44538 21734 44590 21786
rect 58726 21734 58778 21786
rect 58790 21734 58842 21786
rect 58854 21734 58906 21786
rect 58918 21734 58970 21786
rect 58982 21734 59034 21786
rect 5172 21632 5224 21684
rect 6460 21632 6512 21684
rect 5356 21564 5408 21616
rect 7656 21632 7708 21684
rect 9404 21632 9456 21684
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 24860 21632 24912 21684
rect 25688 21632 25740 21684
rect 30196 21632 30248 21684
rect 30656 21632 30708 21684
rect 31392 21675 31444 21684
rect 31392 21641 31401 21675
rect 31401 21641 31435 21675
rect 31435 21641 31444 21675
rect 31392 21632 31444 21641
rect 33048 21632 33100 21684
rect 35440 21632 35492 21684
rect 35716 21632 35768 21684
rect 43720 21632 43772 21684
rect 46204 21632 46256 21684
rect 46940 21632 46992 21684
rect 48228 21675 48280 21684
rect 48228 21641 48237 21675
rect 48237 21641 48271 21675
rect 48271 21641 48280 21675
rect 48228 21632 48280 21641
rect 50988 21675 51040 21684
rect 50988 21641 50997 21675
rect 50997 21641 51031 21675
rect 51031 21641 51040 21675
rect 50988 21632 51040 21641
rect 51172 21632 51224 21684
rect 55404 21632 55456 21684
rect 55956 21632 56008 21684
rect 56692 21675 56744 21684
rect 56692 21641 56701 21675
rect 56701 21641 56735 21675
rect 56735 21641 56744 21675
rect 56692 21632 56744 21641
rect 57980 21632 58032 21684
rect 7196 21539 7248 21548
rect 7196 21505 7214 21539
rect 7214 21505 7248 21539
rect 7196 21496 7248 21505
rect 7288 21539 7340 21548
rect 7288 21505 7297 21539
rect 7297 21505 7331 21539
rect 7331 21505 7340 21539
rect 7288 21496 7340 21505
rect 13820 21564 13872 21616
rect 29000 21564 29052 21616
rect 51356 21564 51408 21616
rect 52828 21564 52880 21616
rect 55220 21564 55272 21616
rect 8300 21539 8352 21548
rect 8300 21505 8309 21539
rect 8309 21505 8343 21539
rect 8343 21505 8352 21539
rect 8300 21496 8352 21505
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 7012 21471 7064 21480
rect 7012 21437 7021 21471
rect 7021 21437 7055 21471
rect 7055 21437 7064 21471
rect 7012 21428 7064 21437
rect 5908 21292 5960 21344
rect 7288 21292 7340 21344
rect 7932 21428 7984 21480
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 13912 21539 13964 21548
rect 13912 21505 13921 21539
rect 13921 21505 13955 21539
rect 13955 21505 13964 21539
rect 13912 21496 13964 21505
rect 29276 21539 29328 21548
rect 29276 21505 29285 21539
rect 29285 21505 29319 21539
rect 29319 21505 29328 21539
rect 29276 21496 29328 21505
rect 30380 21539 30432 21548
rect 30380 21505 30389 21539
rect 30389 21505 30423 21539
rect 30423 21505 30432 21539
rect 30380 21496 30432 21505
rect 42248 21496 42300 21548
rect 46480 21496 46532 21548
rect 47308 21496 47360 21548
rect 48964 21539 49016 21548
rect 48964 21505 48973 21539
rect 48973 21505 49007 21539
rect 49007 21505 49016 21539
rect 48964 21496 49016 21505
rect 12348 21428 12400 21480
rect 14464 21428 14516 21480
rect 13176 21360 13228 21412
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 19064 21471 19116 21480
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 17040 21360 17092 21412
rect 36728 21428 36780 21480
rect 42524 21428 42576 21480
rect 48596 21428 48648 21480
rect 29644 21360 29696 21412
rect 50252 21471 50304 21480
rect 50252 21437 50261 21471
rect 50261 21437 50295 21471
rect 50295 21437 50304 21471
rect 50252 21428 50304 21437
rect 50804 21428 50856 21480
rect 51264 21428 51316 21480
rect 52736 21496 52788 21548
rect 55772 21496 55824 21548
rect 57612 21428 57664 21480
rect 8024 21292 8076 21344
rect 8484 21292 8536 21344
rect 8760 21292 8812 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 10508 21335 10560 21344
rect 10508 21301 10517 21335
rect 10517 21301 10551 21335
rect 10551 21301 10560 21335
rect 10508 21292 10560 21301
rect 10692 21292 10744 21344
rect 11980 21335 12032 21344
rect 11980 21301 11989 21335
rect 11989 21301 12023 21335
rect 12023 21301 12032 21335
rect 11980 21292 12032 21301
rect 12716 21292 12768 21344
rect 13912 21292 13964 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 15292 21292 15344 21344
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 25964 21292 26016 21344
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 28448 21335 28500 21344
rect 28448 21301 28457 21335
rect 28457 21301 28491 21335
rect 28491 21301 28500 21335
rect 28448 21292 28500 21301
rect 31024 21335 31076 21344
rect 31024 21301 31033 21335
rect 31033 21301 31067 21335
rect 31067 21301 31076 21335
rect 31024 21292 31076 21301
rect 35624 21335 35676 21344
rect 35624 21301 35633 21335
rect 35633 21301 35667 21335
rect 35667 21301 35676 21335
rect 35624 21292 35676 21301
rect 37832 21292 37884 21344
rect 42156 21335 42208 21344
rect 42156 21301 42165 21335
rect 42165 21301 42199 21335
rect 42199 21301 42208 21335
rect 42156 21292 42208 21301
rect 42616 21292 42668 21344
rect 48412 21335 48464 21344
rect 48412 21301 48421 21335
rect 48421 21301 48455 21335
rect 48455 21301 48464 21335
rect 48412 21292 48464 21301
rect 49056 21292 49108 21344
rect 51356 21292 51408 21344
rect 56784 21292 56836 21344
rect 57888 21335 57940 21344
rect 57888 21301 57897 21335
rect 57897 21301 57931 21335
rect 57931 21301 57940 21335
rect 57888 21292 57940 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 22616 21190 22668 21242
rect 22680 21190 22732 21242
rect 22744 21190 22796 21242
rect 22808 21190 22860 21242
rect 22872 21190 22924 21242
rect 37060 21190 37112 21242
rect 37124 21190 37176 21242
rect 37188 21190 37240 21242
rect 37252 21190 37304 21242
rect 37316 21190 37368 21242
rect 51504 21190 51556 21242
rect 51568 21190 51620 21242
rect 51632 21190 51684 21242
rect 51696 21190 51748 21242
rect 51760 21190 51812 21242
rect 4160 21088 4212 21140
rect 7288 21088 7340 21140
rect 7564 21088 7616 21140
rect 10692 21088 10744 21140
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 9680 20952 9732 21004
rect 10324 20952 10376 21004
rect 11980 21020 12032 21072
rect 12348 21088 12400 21140
rect 16120 21088 16172 21140
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 28264 21131 28316 21140
rect 28264 21097 28273 21131
rect 28273 21097 28307 21131
rect 28307 21097 28316 21131
rect 28264 21088 28316 21097
rect 28448 21088 28500 21140
rect 33324 21088 33376 21140
rect 34060 21088 34112 21140
rect 5540 20816 5592 20868
rect 7196 20816 7248 20868
rect 6000 20748 6052 20800
rect 7472 20748 7524 20800
rect 10508 20884 10560 20936
rect 8024 20816 8076 20868
rect 13452 20927 13504 20936
rect 13452 20893 13461 20927
rect 13461 20893 13495 20927
rect 13495 20893 13504 20927
rect 13452 20884 13504 20893
rect 18604 20952 18656 21004
rect 38292 21020 38344 21072
rect 36728 20952 36780 21004
rect 37832 20952 37884 21004
rect 46388 21088 46440 21140
rect 46756 21088 46808 21140
rect 50252 21088 50304 21140
rect 44824 21020 44876 21072
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 19340 20927 19392 20936
rect 19340 20893 19349 20927
rect 19349 20893 19383 20927
rect 19383 20893 19392 20927
rect 19340 20884 19392 20893
rect 23020 20884 23072 20936
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 25228 20927 25280 20936
rect 25228 20893 25237 20927
rect 25237 20893 25271 20927
rect 25271 20893 25280 20927
rect 25228 20884 25280 20893
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 25780 20884 25832 20936
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 27528 20884 27580 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 34152 20927 34204 20936
rect 34152 20893 34161 20927
rect 34161 20893 34195 20927
rect 34195 20893 34204 20927
rect 34152 20884 34204 20893
rect 37556 20927 37608 20936
rect 37556 20893 37565 20927
rect 37565 20893 37599 20927
rect 37599 20893 37608 20927
rect 37556 20884 37608 20893
rect 37740 20927 37792 20936
rect 37740 20893 37749 20927
rect 37749 20893 37783 20927
rect 37783 20893 37792 20927
rect 37740 20884 37792 20893
rect 38936 20927 38988 20936
rect 38936 20893 38945 20927
rect 38945 20893 38979 20927
rect 38979 20893 38988 20927
rect 38936 20884 38988 20893
rect 40500 20884 40552 20936
rect 42340 20884 42392 20936
rect 43168 20884 43220 20936
rect 44180 20884 44232 20936
rect 36728 20816 36780 20868
rect 43904 20816 43956 20868
rect 52092 21088 52144 21140
rect 52368 21088 52420 21140
rect 57612 21131 57664 21140
rect 57612 21097 57621 21131
rect 57621 21097 57655 21131
rect 57655 21097 57664 21131
rect 57612 21088 57664 21097
rect 57888 21088 57940 21140
rect 52184 20927 52236 20936
rect 52184 20893 52193 20927
rect 52193 20893 52227 20927
rect 52227 20893 52236 20927
rect 52184 20884 52236 20893
rect 53564 20884 53616 20936
rect 54300 20927 54352 20936
rect 54300 20893 54309 20927
rect 54309 20893 54343 20927
rect 54343 20893 54352 20927
rect 54300 20884 54352 20893
rect 55680 20884 55732 20936
rect 53840 20816 53892 20868
rect 56784 20816 56836 20868
rect 7932 20748 7984 20800
rect 12808 20791 12860 20800
rect 12808 20757 12817 20791
rect 12817 20757 12851 20791
rect 12851 20757 12860 20791
rect 12808 20748 12860 20757
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 15844 20748 15896 20800
rect 19524 20748 19576 20800
rect 22008 20748 22060 20800
rect 22376 20748 22428 20800
rect 22468 20748 22520 20800
rect 24584 20791 24636 20800
rect 24584 20757 24593 20791
rect 24593 20757 24627 20791
rect 24627 20757 24636 20791
rect 24584 20748 24636 20757
rect 26056 20748 26108 20800
rect 26516 20748 26568 20800
rect 26884 20748 26936 20800
rect 30380 20791 30432 20800
rect 30380 20757 30389 20791
rect 30389 20757 30423 20791
rect 30423 20757 30432 20791
rect 30380 20748 30432 20757
rect 32680 20748 32732 20800
rect 33600 20791 33652 20800
rect 33600 20757 33609 20791
rect 33609 20757 33643 20791
rect 33643 20757 33652 20791
rect 33600 20748 33652 20757
rect 36912 20748 36964 20800
rect 38384 20791 38436 20800
rect 38384 20757 38393 20791
rect 38393 20757 38427 20791
rect 38427 20757 38436 20791
rect 38384 20748 38436 20757
rect 38752 20791 38804 20800
rect 38752 20757 38761 20791
rect 38761 20757 38795 20791
rect 38795 20757 38804 20791
rect 38752 20748 38804 20757
rect 39580 20791 39632 20800
rect 39580 20757 39589 20791
rect 39589 20757 39623 20791
rect 39623 20757 39632 20791
rect 39580 20748 39632 20757
rect 40224 20791 40276 20800
rect 40224 20757 40233 20791
rect 40233 20757 40267 20791
rect 40267 20757 40276 20791
rect 40224 20748 40276 20757
rect 40408 20748 40460 20800
rect 42892 20748 42944 20800
rect 43076 20791 43128 20800
rect 43076 20757 43085 20791
rect 43085 20757 43119 20791
rect 43119 20757 43128 20791
rect 43076 20748 43128 20757
rect 44640 20748 44692 20800
rect 45560 20791 45612 20800
rect 45560 20757 45569 20791
rect 45569 20757 45603 20791
rect 45603 20757 45612 20791
rect 45560 20748 45612 20757
rect 53196 20748 53248 20800
rect 54024 20748 54076 20800
rect 54852 20791 54904 20800
rect 54852 20757 54861 20791
rect 54861 20757 54895 20791
rect 54895 20757 54904 20791
rect 54852 20748 54904 20757
rect 56324 20748 56376 20800
rect 57520 20791 57572 20800
rect 57520 20757 57529 20791
rect 57529 20757 57563 20791
rect 57563 20757 57572 20791
rect 57520 20748 57572 20757
rect 57980 20791 58032 20800
rect 57980 20757 57989 20791
rect 57989 20757 58023 20791
rect 58023 20757 58032 20791
rect 57980 20748 58032 20757
rect 58072 20791 58124 20800
rect 58072 20757 58081 20791
rect 58081 20757 58115 20791
rect 58115 20757 58124 20791
rect 58072 20748 58124 20757
rect 15394 20646 15446 20698
rect 15458 20646 15510 20698
rect 15522 20646 15574 20698
rect 15586 20646 15638 20698
rect 15650 20646 15702 20698
rect 29838 20646 29890 20698
rect 29902 20646 29954 20698
rect 29966 20646 30018 20698
rect 30030 20646 30082 20698
rect 30094 20646 30146 20698
rect 44282 20646 44334 20698
rect 44346 20646 44398 20698
rect 44410 20646 44462 20698
rect 44474 20646 44526 20698
rect 44538 20646 44590 20698
rect 58726 20646 58778 20698
rect 58790 20646 58842 20698
rect 58854 20646 58906 20698
rect 58918 20646 58970 20698
rect 58982 20646 59034 20698
rect 5540 20544 5592 20596
rect 7196 20544 7248 20596
rect 13452 20544 13504 20596
rect 14004 20544 14056 20596
rect 15292 20544 15344 20596
rect 16580 20544 16632 20596
rect 16672 20544 16724 20596
rect 17316 20544 17368 20596
rect 19340 20544 19392 20596
rect 22468 20544 22520 20596
rect 7932 20476 7984 20528
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 9680 20451 9732 20460
rect 9680 20417 9714 20451
rect 9714 20417 9732 20451
rect 9680 20408 9732 20417
rect 10416 20408 10468 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 16396 20476 16448 20528
rect 18052 20476 18104 20528
rect 19616 20519 19668 20528
rect 19616 20485 19634 20519
rect 19634 20485 19668 20519
rect 19616 20476 19668 20485
rect 21180 20476 21232 20528
rect 24860 20544 24912 20596
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 26332 20544 26384 20596
rect 26700 20544 26752 20596
rect 29736 20544 29788 20596
rect 30932 20544 30984 20596
rect 38108 20544 38160 20596
rect 38752 20544 38804 20596
rect 38936 20544 38988 20596
rect 42892 20587 42944 20596
rect 42892 20553 42901 20587
rect 42901 20553 42935 20587
rect 42935 20553 42944 20587
rect 42892 20544 42944 20553
rect 43720 20544 43772 20596
rect 44732 20587 44784 20596
rect 44732 20553 44741 20587
rect 44741 20553 44775 20587
rect 44775 20553 44784 20587
rect 44732 20544 44784 20553
rect 48412 20544 48464 20596
rect 52184 20544 52236 20596
rect 53564 20587 53616 20596
rect 53564 20553 53573 20587
rect 53573 20553 53607 20587
rect 53607 20553 53616 20587
rect 53564 20544 53616 20553
rect 54024 20587 54076 20596
rect 54024 20553 54033 20587
rect 54033 20553 54067 20587
rect 54067 20553 54076 20587
rect 54024 20544 54076 20553
rect 55772 20544 55824 20596
rect 57428 20544 57480 20596
rect 24584 20476 24636 20528
rect 25412 20476 25464 20528
rect 28080 20476 28132 20528
rect 38660 20476 38712 20528
rect 40224 20476 40276 20528
rect 42984 20476 43036 20528
rect 49424 20476 49476 20528
rect 50160 20476 50212 20528
rect 7472 20340 7524 20392
rect 9036 20340 9088 20392
rect 10876 20340 10928 20392
rect 14556 20340 14608 20392
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 11704 20247 11756 20256
rect 11704 20213 11713 20247
rect 11713 20213 11747 20247
rect 11747 20213 11756 20247
rect 11704 20204 11756 20213
rect 13176 20204 13228 20256
rect 20536 20408 20588 20460
rect 21272 20408 21324 20460
rect 26056 20408 26108 20460
rect 26424 20408 26476 20460
rect 33508 20408 33560 20460
rect 33876 20408 33928 20460
rect 37648 20451 37700 20460
rect 37648 20417 37657 20451
rect 37657 20417 37691 20451
rect 37691 20417 37700 20451
rect 37648 20408 37700 20417
rect 38568 20408 38620 20460
rect 40868 20408 40920 20460
rect 18236 20383 18288 20392
rect 18236 20349 18245 20383
rect 18245 20349 18279 20383
rect 18279 20349 18288 20383
rect 18236 20340 18288 20349
rect 19984 20383 20036 20392
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 22008 20340 22060 20392
rect 20444 20272 20496 20324
rect 21456 20272 21508 20324
rect 25228 20340 25280 20392
rect 25964 20383 26016 20392
rect 25964 20349 25973 20383
rect 25973 20349 26007 20383
rect 26007 20349 26016 20383
rect 25964 20340 26016 20349
rect 26608 20340 26660 20392
rect 27252 20340 27304 20392
rect 29000 20340 29052 20392
rect 31116 20383 31168 20392
rect 31116 20349 31125 20383
rect 31125 20349 31159 20383
rect 31159 20349 31168 20383
rect 31116 20340 31168 20349
rect 32588 20383 32640 20392
rect 32588 20349 32597 20383
rect 32597 20349 32631 20383
rect 32631 20349 32640 20383
rect 32588 20340 32640 20349
rect 32680 20383 32732 20392
rect 32680 20349 32689 20383
rect 32689 20349 32723 20383
rect 32723 20349 32732 20383
rect 32680 20340 32732 20349
rect 32956 20383 33008 20392
rect 32956 20349 32965 20383
rect 32965 20349 32999 20383
rect 32999 20349 33008 20383
rect 32956 20340 33008 20349
rect 35808 20383 35860 20392
rect 35808 20349 35817 20383
rect 35817 20349 35851 20383
rect 35851 20349 35860 20383
rect 35808 20340 35860 20349
rect 15292 20204 15344 20256
rect 17592 20204 17644 20256
rect 17868 20204 17920 20256
rect 19708 20204 19760 20256
rect 21548 20204 21600 20256
rect 21824 20204 21876 20256
rect 23204 20247 23256 20256
rect 23204 20213 23213 20247
rect 23213 20213 23247 20247
rect 23247 20213 23256 20247
rect 23204 20204 23256 20213
rect 23940 20204 23992 20256
rect 24860 20204 24912 20256
rect 26148 20204 26200 20256
rect 27344 20204 27396 20256
rect 28448 20247 28500 20256
rect 28448 20213 28457 20247
rect 28457 20213 28491 20247
rect 28491 20213 28500 20247
rect 28448 20204 28500 20213
rect 29460 20247 29512 20256
rect 29460 20213 29469 20247
rect 29469 20213 29503 20247
rect 29503 20213 29512 20247
rect 29460 20204 29512 20213
rect 31392 20204 31444 20256
rect 37464 20383 37516 20392
rect 37464 20349 37473 20383
rect 37473 20349 37507 20383
rect 37507 20349 37516 20383
rect 37464 20340 37516 20349
rect 37832 20340 37884 20392
rect 38108 20340 38160 20392
rect 38844 20340 38896 20392
rect 36912 20272 36964 20324
rect 35716 20204 35768 20256
rect 35992 20247 36044 20256
rect 35992 20213 36001 20247
rect 36001 20213 36035 20247
rect 36035 20213 36044 20247
rect 35992 20204 36044 20213
rect 37832 20204 37884 20256
rect 38016 20247 38068 20256
rect 38016 20213 38025 20247
rect 38025 20213 38059 20247
rect 38059 20213 38068 20247
rect 38016 20204 38068 20213
rect 43812 20408 43864 20460
rect 43260 20383 43312 20392
rect 43260 20349 43269 20383
rect 43269 20349 43303 20383
rect 43303 20349 43312 20383
rect 43260 20340 43312 20349
rect 46756 20408 46808 20460
rect 44456 20340 44508 20392
rect 44640 20340 44692 20392
rect 45284 20383 45336 20392
rect 45284 20349 45293 20383
rect 45293 20349 45327 20383
rect 45327 20349 45336 20383
rect 45284 20340 45336 20349
rect 43628 20272 43680 20324
rect 43996 20272 44048 20324
rect 44824 20272 44876 20324
rect 49148 20383 49200 20392
rect 49148 20349 49157 20383
rect 49157 20349 49191 20383
rect 49191 20349 49200 20383
rect 49148 20340 49200 20349
rect 52736 20408 52788 20460
rect 47492 20272 47544 20324
rect 39120 20204 39172 20256
rect 41052 20247 41104 20256
rect 41052 20213 41061 20247
rect 41061 20213 41095 20247
rect 41095 20213 41104 20247
rect 41052 20204 41104 20213
rect 41420 20247 41472 20256
rect 41420 20213 41429 20247
rect 41429 20213 41463 20247
rect 41463 20213 41472 20247
rect 41420 20204 41472 20213
rect 41696 20204 41748 20256
rect 45100 20204 45152 20256
rect 45928 20247 45980 20256
rect 45928 20213 45937 20247
rect 45937 20213 45971 20247
rect 45971 20213 45980 20247
rect 45928 20204 45980 20213
rect 46664 20247 46716 20256
rect 46664 20213 46673 20247
rect 46673 20213 46707 20247
rect 46707 20213 46716 20247
rect 46664 20204 46716 20213
rect 47308 20247 47360 20256
rect 47308 20213 47317 20247
rect 47317 20213 47351 20247
rect 47351 20213 47360 20247
rect 47308 20204 47360 20213
rect 47860 20204 47912 20256
rect 52368 20204 52420 20256
rect 55404 20451 55456 20460
rect 55404 20417 55413 20451
rect 55413 20417 55447 20451
rect 55447 20417 55456 20451
rect 55404 20408 55456 20417
rect 58072 20476 58124 20528
rect 54024 20340 54076 20392
rect 55588 20383 55640 20392
rect 55588 20349 55606 20383
rect 55606 20349 55640 20383
rect 55588 20340 55640 20349
rect 54852 20272 54904 20324
rect 54484 20204 54536 20256
rect 56048 20340 56100 20392
rect 56324 20340 56376 20392
rect 56968 20340 57020 20392
rect 57520 20408 57572 20460
rect 57428 20272 57480 20324
rect 56692 20247 56744 20256
rect 56692 20213 56701 20247
rect 56701 20213 56735 20247
rect 56735 20213 56744 20247
rect 56692 20204 56744 20213
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 22616 20102 22668 20154
rect 22680 20102 22732 20154
rect 22744 20102 22796 20154
rect 22808 20102 22860 20154
rect 22872 20102 22924 20154
rect 37060 20102 37112 20154
rect 37124 20102 37176 20154
rect 37188 20102 37240 20154
rect 37252 20102 37304 20154
rect 37316 20102 37368 20154
rect 51504 20102 51556 20154
rect 51568 20102 51620 20154
rect 51632 20102 51684 20154
rect 51696 20102 51748 20154
rect 51760 20102 51812 20154
rect 9680 20000 9732 20052
rect 16948 20000 17000 20052
rect 19064 20043 19116 20052
rect 19064 20009 19073 20043
rect 19073 20009 19107 20043
rect 19107 20009 19116 20043
rect 19064 20000 19116 20009
rect 21088 20000 21140 20052
rect 21456 20000 21508 20052
rect 7380 19864 7432 19916
rect 7840 19864 7892 19916
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 2780 19796 2832 19848
rect 3424 19839 3476 19848
rect 3424 19805 3433 19839
rect 3433 19805 3467 19839
rect 3467 19805 3476 19839
rect 3424 19796 3476 19805
rect 3516 19796 3568 19848
rect 6920 19839 6972 19848
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 9772 19796 9824 19848
rect 6276 19771 6328 19780
rect 6276 19737 6285 19771
rect 6285 19737 6319 19771
rect 6319 19737 6328 19771
rect 6276 19728 6328 19737
rect 14648 19907 14700 19916
rect 14648 19873 14657 19907
rect 14657 19873 14691 19907
rect 14691 19873 14700 19907
rect 19524 19932 19576 19984
rect 14648 19864 14700 19873
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 18604 19864 18656 19916
rect 17040 19796 17092 19848
rect 17592 19839 17644 19848
rect 17592 19805 17610 19839
rect 17610 19805 17644 19839
rect 17592 19796 17644 19805
rect 13360 19728 13412 19780
rect 2964 19660 3016 19712
rect 3976 19660 4028 19712
rect 4528 19660 4580 19712
rect 7012 19703 7064 19712
rect 7012 19669 7021 19703
rect 7021 19669 7055 19703
rect 7055 19669 7064 19703
rect 7012 19660 7064 19669
rect 7380 19660 7432 19712
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 10600 19703 10652 19712
rect 10600 19669 10609 19703
rect 10609 19669 10643 19703
rect 10643 19669 10652 19703
rect 10600 19660 10652 19669
rect 10876 19660 10928 19712
rect 13728 19660 13780 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 18052 19660 18104 19712
rect 18788 19728 18840 19780
rect 19524 19796 19576 19848
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 20536 19864 20588 19916
rect 21456 19907 21508 19916
rect 21456 19873 21465 19907
rect 21465 19873 21499 19907
rect 21499 19873 21508 19907
rect 21456 19864 21508 19873
rect 18972 19728 19024 19780
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 22468 20000 22520 20052
rect 23664 20000 23716 20052
rect 24860 20000 24912 20052
rect 26424 20000 26476 20052
rect 27528 20043 27580 20052
rect 27528 20009 27537 20043
rect 27537 20009 27571 20043
rect 27571 20009 27580 20043
rect 27528 20000 27580 20009
rect 31116 20000 31168 20052
rect 32956 20000 33008 20052
rect 35808 20000 35860 20052
rect 35992 20000 36044 20052
rect 37740 20000 37792 20052
rect 38844 20000 38896 20052
rect 39120 20000 39172 20052
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 26792 19975 26844 19984
rect 26792 19941 26801 19975
rect 26801 19941 26835 19975
rect 26835 19941 26844 19975
rect 26792 19932 26844 19941
rect 35624 19932 35676 19984
rect 19524 19660 19576 19712
rect 19892 19660 19944 19712
rect 20628 19660 20680 19712
rect 21732 19660 21784 19712
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 26056 19864 26108 19916
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 26700 19864 26752 19916
rect 26884 19864 26936 19916
rect 23204 19796 23256 19848
rect 26240 19839 26292 19848
rect 26240 19805 26249 19839
rect 26249 19805 26283 19839
rect 26283 19805 26292 19839
rect 26240 19796 26292 19805
rect 27804 19864 27856 19916
rect 33324 19907 33376 19916
rect 33324 19873 33333 19907
rect 33333 19873 33367 19907
rect 33367 19873 33376 19907
rect 33324 19864 33376 19873
rect 33508 19907 33560 19916
rect 33508 19873 33526 19907
rect 33526 19873 33560 19907
rect 33508 19864 33560 19873
rect 25044 19728 25096 19780
rect 30380 19796 30432 19848
rect 31392 19839 31444 19848
rect 31392 19805 31426 19839
rect 31426 19805 31444 19839
rect 24952 19660 25004 19712
rect 25136 19703 25188 19712
rect 25136 19669 25145 19703
rect 25145 19669 25179 19703
rect 25179 19669 25188 19703
rect 25136 19660 25188 19669
rect 26516 19660 26568 19712
rect 26976 19660 27028 19712
rect 28448 19728 28500 19780
rect 31392 19796 31444 19805
rect 33600 19839 33652 19848
rect 33600 19805 33609 19839
rect 33609 19805 33643 19839
rect 33643 19805 33652 19839
rect 33600 19796 33652 19805
rect 34520 19839 34572 19848
rect 34520 19805 34529 19839
rect 34529 19805 34563 19839
rect 34563 19805 34572 19839
rect 34520 19796 34572 19805
rect 34796 19907 34848 19916
rect 34796 19873 34805 19907
rect 34805 19873 34839 19907
rect 34839 19873 34848 19907
rect 34796 19864 34848 19873
rect 35808 19864 35860 19916
rect 38200 19864 38252 19916
rect 38660 19907 38712 19916
rect 38660 19873 38669 19907
rect 38669 19873 38703 19907
rect 38703 19873 38712 19907
rect 38660 19864 38712 19873
rect 39028 19864 39080 19916
rect 36176 19796 36228 19848
rect 36912 19796 36964 19848
rect 38476 19796 38528 19848
rect 40040 19864 40092 19916
rect 40408 19907 40460 19916
rect 40408 19873 40417 19907
rect 40417 19873 40451 19907
rect 40451 19873 40460 19907
rect 43260 20000 43312 20052
rect 45284 20000 45336 20052
rect 48596 20043 48648 20052
rect 48596 20009 48605 20043
rect 48605 20009 48639 20043
rect 48639 20009 48648 20043
rect 48596 20000 48648 20009
rect 49148 20000 49200 20052
rect 42984 19975 43036 19984
rect 42984 19941 42993 19975
rect 42993 19941 43027 19975
rect 43027 19941 43036 19975
rect 42984 19932 43036 19941
rect 40408 19864 40460 19873
rect 41052 19796 41104 19848
rect 36728 19728 36780 19780
rect 31116 19660 31168 19712
rect 32680 19703 32732 19712
rect 32680 19669 32689 19703
rect 32689 19669 32723 19703
rect 32723 19669 32732 19703
rect 32680 19660 32732 19669
rect 34888 19660 34940 19712
rect 39856 19703 39908 19712
rect 39856 19669 39865 19703
rect 39865 19669 39899 19703
rect 39899 19669 39908 19703
rect 39856 19660 39908 19669
rect 43628 19907 43680 19916
rect 43628 19873 43637 19907
rect 43637 19873 43671 19907
rect 43671 19873 43680 19907
rect 43628 19864 43680 19873
rect 43812 19907 43864 19916
rect 43812 19873 43830 19907
rect 43830 19873 43864 19907
rect 43812 19864 43864 19873
rect 43904 19907 43956 19916
rect 43904 19873 43913 19907
rect 43913 19873 43947 19907
rect 43947 19873 43956 19907
rect 43904 19864 43956 19873
rect 44916 19864 44968 19916
rect 41236 19839 41288 19848
rect 41236 19805 41245 19839
rect 41245 19805 41279 19839
rect 41279 19805 41288 19839
rect 41236 19796 41288 19805
rect 41696 19839 41748 19848
rect 41696 19805 41730 19839
rect 41730 19805 41748 19839
rect 41696 19796 41748 19805
rect 45008 19796 45060 19848
rect 47216 19907 47268 19916
rect 47216 19873 47225 19907
rect 47225 19873 47259 19907
rect 47259 19873 47268 19907
rect 47216 19864 47268 19873
rect 50160 19907 50212 19916
rect 50160 19873 50169 19907
rect 50169 19873 50203 19907
rect 50203 19873 50212 19907
rect 50160 19864 50212 19873
rect 52368 20043 52420 20052
rect 52368 20009 52377 20043
rect 52377 20009 52411 20043
rect 52411 20009 52420 20043
rect 52368 20000 52420 20009
rect 52736 20000 52788 20052
rect 55036 20043 55088 20052
rect 55036 20009 55045 20043
rect 55045 20009 55079 20043
rect 55079 20009 55088 20043
rect 55036 20000 55088 20009
rect 52000 19932 52052 19984
rect 51816 19907 51868 19916
rect 51816 19873 51825 19907
rect 51825 19873 51859 19907
rect 51859 19873 51868 19907
rect 51816 19864 51868 19873
rect 45560 19796 45612 19848
rect 45744 19796 45796 19848
rect 49056 19839 49108 19848
rect 49056 19805 49065 19839
rect 49065 19805 49099 19839
rect 49099 19805 49108 19839
rect 49056 19796 49108 19805
rect 52092 19796 52144 19848
rect 53932 19864 53984 19916
rect 58164 20000 58216 20052
rect 58440 19932 58492 19984
rect 54116 19796 54168 19848
rect 55680 19839 55732 19848
rect 55680 19805 55689 19839
rect 55689 19805 55723 19839
rect 55723 19805 55732 19839
rect 55680 19796 55732 19805
rect 56968 19796 57020 19848
rect 45928 19728 45980 19780
rect 47492 19771 47544 19780
rect 47492 19737 47526 19771
rect 47526 19737 47544 19771
rect 47492 19728 47544 19737
rect 50252 19728 50304 19780
rect 54392 19728 54444 19780
rect 55588 19728 55640 19780
rect 56508 19728 56560 19780
rect 44456 19660 44508 19712
rect 48320 19660 48372 19712
rect 49792 19660 49844 19712
rect 51264 19660 51316 19712
rect 52276 19660 52328 19712
rect 54208 19703 54260 19712
rect 54208 19669 54217 19703
rect 54217 19669 54251 19703
rect 54251 19669 54260 19703
rect 54208 19660 54260 19669
rect 54484 19660 54536 19712
rect 58072 19660 58124 19712
rect 15394 19558 15446 19610
rect 15458 19558 15510 19610
rect 15522 19558 15574 19610
rect 15586 19558 15638 19610
rect 15650 19558 15702 19610
rect 29838 19558 29890 19610
rect 29902 19558 29954 19610
rect 29966 19558 30018 19610
rect 30030 19558 30082 19610
rect 30094 19558 30146 19610
rect 44282 19558 44334 19610
rect 44346 19558 44398 19610
rect 44410 19558 44462 19610
rect 44474 19558 44526 19610
rect 44538 19558 44590 19610
rect 58726 19558 58778 19610
rect 58790 19558 58842 19610
rect 58854 19558 58906 19610
rect 58918 19558 58970 19610
rect 58982 19558 59034 19610
rect 2136 19456 2188 19508
rect 2872 19456 2924 19508
rect 3424 19499 3476 19508
rect 3424 19465 3433 19499
rect 3433 19465 3467 19499
rect 3467 19465 3476 19499
rect 3424 19456 3476 19465
rect 4528 19456 4580 19508
rect 6276 19456 6328 19508
rect 7564 19456 7616 19508
rect 13360 19456 13412 19508
rect 16672 19456 16724 19508
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 18236 19456 18288 19508
rect 19892 19456 19944 19508
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 20996 19456 21048 19508
rect 22376 19456 22428 19508
rect 23020 19456 23072 19508
rect 25780 19456 25832 19508
rect 26700 19456 26752 19508
rect 27252 19456 27304 19508
rect 28724 19456 28776 19508
rect 3884 19431 3936 19440
rect 3884 19397 3893 19431
rect 3893 19397 3927 19431
rect 3927 19397 3936 19431
rect 3884 19388 3936 19397
rect 4068 19320 4120 19372
rect 12808 19388 12860 19440
rect 9864 19320 9916 19372
rect 12532 19320 12584 19372
rect 14096 19320 14148 19372
rect 15200 19320 15252 19372
rect 15660 19320 15712 19372
rect 15844 19320 15896 19372
rect 21180 19388 21232 19440
rect 21732 19388 21784 19440
rect 19248 19320 19300 19372
rect 20720 19320 20772 19372
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 23940 19388 23992 19440
rect 21916 19320 21968 19372
rect 24400 19363 24452 19372
rect 24400 19329 24434 19363
rect 24434 19329 24452 19363
rect 24400 19320 24452 19329
rect 25136 19320 25188 19372
rect 26332 19320 26384 19372
rect 2044 19116 2096 19168
rect 3332 19116 3384 19168
rect 4160 19252 4212 19304
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 7380 19252 7432 19304
rect 7564 19252 7616 19304
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 10600 19252 10652 19304
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 31024 19456 31076 19508
rect 32680 19456 32732 19508
rect 35532 19499 35584 19508
rect 35532 19465 35541 19499
rect 35541 19465 35575 19499
rect 35575 19465 35584 19499
rect 35532 19456 35584 19465
rect 35808 19456 35860 19508
rect 27252 19363 27304 19372
rect 27252 19329 27286 19363
rect 27286 19329 27304 19363
rect 27252 19320 27304 19329
rect 27528 19320 27580 19372
rect 31116 19388 31168 19440
rect 30564 19363 30616 19372
rect 30564 19329 30573 19363
rect 30573 19329 30607 19363
rect 30607 19329 30616 19363
rect 30564 19320 30616 19329
rect 33876 19388 33928 19440
rect 37556 19456 37608 19508
rect 38384 19456 38436 19508
rect 39120 19456 39172 19508
rect 41236 19456 41288 19508
rect 44180 19456 44232 19508
rect 45928 19456 45980 19508
rect 49700 19456 49752 19508
rect 50252 19456 50304 19508
rect 51356 19456 51408 19508
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 5356 19116 5408 19168
rect 7104 19116 7156 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7656 19116 7708 19168
rect 7932 19116 7984 19168
rect 9404 19116 9456 19168
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 14556 19116 14608 19168
rect 18604 19116 18656 19168
rect 20444 19116 20496 19168
rect 20904 19116 20956 19168
rect 23388 19116 23440 19168
rect 25412 19116 25464 19168
rect 26056 19116 26108 19168
rect 30104 19252 30156 19304
rect 31392 19295 31444 19304
rect 31392 19261 31401 19295
rect 31401 19261 31435 19295
rect 31435 19261 31444 19295
rect 31392 19252 31444 19261
rect 34152 19320 34204 19372
rect 37832 19388 37884 19440
rect 36176 19320 36228 19372
rect 35624 19295 35676 19304
rect 35624 19261 35633 19295
rect 35633 19261 35667 19295
rect 35667 19261 35676 19295
rect 35624 19252 35676 19261
rect 35716 19252 35768 19304
rect 36084 19252 36136 19304
rect 37464 19320 37516 19372
rect 38476 19320 38528 19372
rect 39580 19388 39632 19440
rect 40500 19388 40552 19440
rect 41052 19388 41104 19440
rect 36452 19295 36504 19304
rect 36452 19261 36461 19295
rect 36461 19261 36495 19295
rect 36495 19261 36504 19295
rect 36452 19252 36504 19261
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 35532 19184 35584 19236
rect 30656 19116 30708 19168
rect 33600 19159 33652 19168
rect 33600 19125 33609 19159
rect 33609 19125 33643 19159
rect 33643 19125 33652 19159
rect 33600 19116 33652 19125
rect 35072 19159 35124 19168
rect 35072 19125 35081 19159
rect 35081 19125 35115 19159
rect 35115 19125 35124 19159
rect 35072 19116 35124 19125
rect 38292 19159 38344 19168
rect 38292 19125 38301 19159
rect 38301 19125 38335 19159
rect 38335 19125 38344 19159
rect 38292 19116 38344 19125
rect 40868 19320 40920 19372
rect 43076 19320 43128 19372
rect 43720 19320 43772 19372
rect 45468 19320 45520 19372
rect 45744 19320 45796 19372
rect 46112 19363 46164 19372
rect 46112 19329 46146 19363
rect 46146 19329 46164 19363
rect 46112 19320 46164 19329
rect 47216 19320 47268 19372
rect 51264 19388 51316 19440
rect 51816 19456 51868 19508
rect 52736 19456 52788 19508
rect 54300 19499 54352 19508
rect 54300 19465 54309 19499
rect 54309 19465 54343 19499
rect 54343 19465 54352 19499
rect 54300 19456 54352 19465
rect 54392 19499 54444 19508
rect 54392 19465 54401 19499
rect 54401 19465 54435 19499
rect 54435 19465 54444 19499
rect 54392 19456 54444 19465
rect 55588 19456 55640 19508
rect 56692 19456 56744 19508
rect 56968 19456 57020 19508
rect 47860 19363 47912 19372
rect 47860 19329 47894 19363
rect 47894 19329 47912 19363
rect 47860 19320 47912 19329
rect 50160 19320 50212 19372
rect 50988 19320 51040 19372
rect 54116 19388 54168 19440
rect 53196 19363 53248 19372
rect 53196 19329 53230 19363
rect 53230 19329 53248 19363
rect 53196 19320 53248 19329
rect 54208 19320 54260 19372
rect 55036 19363 55088 19372
rect 55036 19329 55045 19363
rect 55045 19329 55079 19363
rect 55079 19329 55088 19363
rect 55036 19320 55088 19329
rect 55680 19320 55732 19372
rect 56232 19363 56284 19372
rect 56232 19329 56241 19363
rect 56241 19329 56275 19363
rect 56275 19329 56284 19363
rect 56232 19320 56284 19329
rect 58440 19363 58492 19372
rect 58440 19329 58449 19363
rect 58449 19329 58483 19363
rect 58483 19329 58492 19363
rect 58440 19320 58492 19329
rect 40776 19295 40828 19304
rect 40776 19261 40785 19295
rect 40785 19261 40819 19295
rect 40819 19261 40828 19295
rect 40776 19252 40828 19261
rect 42432 19295 42484 19304
rect 42432 19261 42441 19295
rect 42441 19261 42475 19295
rect 42475 19261 42484 19295
rect 42432 19252 42484 19261
rect 43904 19252 43956 19304
rect 45008 19252 45060 19304
rect 45100 19295 45152 19304
rect 45100 19261 45109 19295
rect 45109 19261 45143 19295
rect 45143 19261 45152 19295
rect 45100 19252 45152 19261
rect 41420 19116 41472 19168
rect 41788 19116 41840 19168
rect 44640 19159 44692 19168
rect 44640 19125 44649 19159
rect 44649 19125 44683 19159
rect 44683 19125 44692 19159
rect 44640 19116 44692 19125
rect 47400 19184 47452 19236
rect 47216 19159 47268 19168
rect 47216 19125 47225 19159
rect 47225 19125 47259 19159
rect 47259 19125 47268 19159
rect 47216 19116 47268 19125
rect 47308 19116 47360 19168
rect 57612 19159 57664 19168
rect 57612 19125 57621 19159
rect 57621 19125 57655 19159
rect 57655 19125 57664 19159
rect 57612 19116 57664 19125
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 22616 19014 22668 19066
rect 22680 19014 22732 19066
rect 22744 19014 22796 19066
rect 22808 19014 22860 19066
rect 22872 19014 22924 19066
rect 37060 19014 37112 19066
rect 37124 19014 37176 19066
rect 37188 19014 37240 19066
rect 37252 19014 37304 19066
rect 37316 19014 37368 19066
rect 51504 19014 51556 19066
rect 51568 19014 51620 19066
rect 51632 19014 51684 19066
rect 51696 19014 51748 19066
rect 51760 19014 51812 19066
rect 2228 18912 2280 18964
rect 3332 18912 3384 18964
rect 5540 18912 5592 18964
rect 4160 18844 4212 18896
rect 2044 18708 2096 18760
rect 4068 18776 4120 18828
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 4528 18776 4580 18828
rect 5356 18776 5408 18828
rect 6920 18912 6972 18964
rect 7840 18912 7892 18964
rect 9680 18912 9732 18964
rect 10140 18912 10192 18964
rect 15660 18912 15712 18964
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 19248 18955 19300 18964
rect 19248 18921 19257 18955
rect 19257 18921 19291 18955
rect 19291 18921 19300 18955
rect 19248 18912 19300 18921
rect 21088 18912 21140 18964
rect 24400 18912 24452 18964
rect 26976 18912 27028 18964
rect 29092 18912 29144 18964
rect 30104 18912 30156 18964
rect 31392 18912 31444 18964
rect 36452 18912 36504 18964
rect 38660 18912 38712 18964
rect 40776 18912 40828 18964
rect 45008 18955 45060 18964
rect 45008 18921 45017 18955
rect 45017 18921 45051 18955
rect 45051 18921 45060 18955
rect 45008 18912 45060 18921
rect 46112 18912 46164 18964
rect 54116 18955 54168 18964
rect 54116 18921 54125 18955
rect 54125 18921 54159 18955
rect 54159 18921 54168 18955
rect 54116 18912 54168 18921
rect 56508 18912 56560 18964
rect 7656 18776 7708 18828
rect 15292 18776 15344 18828
rect 19524 18776 19576 18828
rect 2964 18708 3016 18760
rect 1860 18572 1912 18624
rect 3792 18640 3844 18692
rect 3700 18572 3752 18624
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 7012 18708 7064 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 10232 18708 10284 18760
rect 17408 18708 17460 18760
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 24952 18776 25004 18828
rect 27160 18776 27212 18828
rect 29460 18844 29512 18896
rect 28356 18776 28408 18828
rect 31944 18819 31996 18828
rect 31944 18785 31953 18819
rect 31953 18785 31987 18819
rect 31987 18785 31996 18819
rect 36084 18844 36136 18896
rect 31944 18776 31996 18785
rect 9220 18640 9272 18692
rect 9404 18640 9456 18692
rect 11704 18640 11756 18692
rect 26608 18708 26660 18760
rect 27804 18751 27856 18760
rect 27804 18717 27813 18751
rect 27813 18717 27847 18751
rect 27847 18717 27856 18751
rect 27804 18708 27856 18717
rect 33508 18708 33560 18760
rect 34520 18776 34572 18828
rect 35072 18776 35124 18828
rect 36176 18776 36228 18828
rect 38016 18776 38068 18828
rect 44640 18819 44692 18828
rect 44640 18785 44649 18819
rect 44649 18785 44683 18819
rect 44683 18785 44692 18819
rect 44640 18776 44692 18785
rect 46112 18776 46164 18828
rect 47308 18776 47360 18828
rect 58164 18776 58216 18828
rect 38108 18708 38160 18760
rect 42432 18708 42484 18760
rect 46664 18708 46716 18760
rect 51816 18751 51868 18760
rect 51816 18717 51825 18751
rect 51825 18717 51859 18751
rect 51859 18717 51868 18751
rect 51816 18708 51868 18717
rect 52460 18751 52512 18760
rect 52460 18717 52469 18751
rect 52469 18717 52503 18751
rect 52503 18717 52512 18751
rect 52460 18708 52512 18717
rect 52552 18708 52604 18760
rect 57152 18751 57204 18760
rect 57152 18717 57161 18751
rect 57161 18717 57195 18751
rect 57195 18717 57204 18751
rect 57152 18708 57204 18717
rect 4712 18572 4764 18624
rect 10692 18572 10744 18624
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 21456 18572 21508 18624
rect 25228 18640 25280 18692
rect 25964 18640 26016 18692
rect 32588 18640 32640 18692
rect 22192 18572 22244 18624
rect 27436 18615 27488 18624
rect 27436 18581 27445 18615
rect 27445 18581 27479 18615
rect 27479 18581 27488 18615
rect 27436 18572 27488 18581
rect 27528 18572 27580 18624
rect 34704 18615 34756 18624
rect 34704 18581 34713 18615
rect 34713 18581 34747 18615
rect 34747 18581 34756 18615
rect 34704 18572 34756 18581
rect 34888 18572 34940 18624
rect 35624 18615 35676 18624
rect 35624 18581 35633 18615
rect 35633 18581 35667 18615
rect 35667 18581 35676 18615
rect 35624 18572 35676 18581
rect 40408 18572 40460 18624
rect 46480 18615 46532 18624
rect 46480 18581 46489 18615
rect 46489 18581 46523 18615
rect 46523 18581 46532 18615
rect 46480 18572 46532 18581
rect 51172 18615 51224 18624
rect 51172 18581 51181 18615
rect 51181 18581 51215 18615
rect 51215 18581 51224 18615
rect 51172 18572 51224 18581
rect 51908 18615 51960 18624
rect 51908 18581 51917 18615
rect 51917 18581 51951 18615
rect 51951 18581 51960 18615
rect 51908 18572 51960 18581
rect 56600 18615 56652 18624
rect 56600 18581 56609 18615
rect 56609 18581 56643 18615
rect 56643 18581 56652 18615
rect 56600 18572 56652 18581
rect 15394 18470 15446 18522
rect 15458 18470 15510 18522
rect 15522 18470 15574 18522
rect 15586 18470 15638 18522
rect 15650 18470 15702 18522
rect 29838 18470 29890 18522
rect 29902 18470 29954 18522
rect 29966 18470 30018 18522
rect 30030 18470 30082 18522
rect 30094 18470 30146 18522
rect 44282 18470 44334 18522
rect 44346 18470 44398 18522
rect 44410 18470 44462 18522
rect 44474 18470 44526 18522
rect 44538 18470 44590 18522
rect 58726 18470 58778 18522
rect 58790 18470 58842 18522
rect 58854 18470 58906 18522
rect 58918 18470 58970 18522
rect 58982 18470 59034 18522
rect 3516 18368 3568 18420
rect 3700 18368 3752 18420
rect 3884 18368 3936 18420
rect 4068 18411 4120 18420
rect 4068 18377 4077 18411
rect 4077 18377 4111 18411
rect 4111 18377 4120 18411
rect 4068 18368 4120 18377
rect 8024 18368 8076 18420
rect 8116 18411 8168 18420
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 17040 18368 17092 18420
rect 20720 18368 20772 18420
rect 27252 18368 27304 18420
rect 27436 18368 27488 18420
rect 34520 18368 34572 18420
rect 35808 18368 35860 18420
rect 51816 18411 51868 18420
rect 51816 18377 51825 18411
rect 51825 18377 51859 18411
rect 51859 18377 51868 18411
rect 51816 18368 51868 18377
rect 51908 18368 51960 18420
rect 52552 18368 52604 18420
rect 57152 18368 57204 18420
rect 2780 18300 2832 18352
rect 7196 18300 7248 18352
rect 2044 18232 2096 18284
rect 4436 18232 4488 18284
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 4252 18096 4304 18148
rect 7104 18232 7156 18284
rect 5540 18164 5592 18216
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 33600 18232 33652 18284
rect 39856 18232 39908 18284
rect 50160 18232 50212 18284
rect 56968 18275 57020 18284
rect 56968 18241 56977 18275
rect 56977 18241 57011 18275
rect 57011 18241 57020 18275
rect 56968 18232 57020 18241
rect 9128 18207 9180 18216
rect 9128 18173 9146 18207
rect 9146 18173 9180 18207
rect 9128 18164 9180 18173
rect 9404 18164 9456 18216
rect 9956 18207 10008 18216
rect 9956 18173 9965 18207
rect 9965 18173 9999 18207
rect 9999 18173 10008 18207
rect 9956 18164 10008 18173
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13360 18164 13412 18216
rect 15108 18164 15160 18216
rect 15752 18164 15804 18216
rect 19156 18207 19208 18216
rect 19156 18173 19165 18207
rect 19165 18173 19199 18207
rect 19199 18173 19208 18207
rect 19156 18164 19208 18173
rect 44640 18207 44692 18216
rect 44640 18173 44649 18207
rect 44649 18173 44683 18207
rect 44683 18173 44692 18207
rect 44640 18164 44692 18173
rect 48412 18207 48464 18216
rect 48412 18173 48421 18207
rect 48421 18173 48455 18207
rect 48455 18173 48464 18207
rect 48412 18164 48464 18173
rect 48780 18207 48832 18216
rect 48780 18173 48789 18207
rect 48789 18173 48823 18207
rect 48823 18173 48832 18207
rect 48780 18164 48832 18173
rect 52552 18207 52604 18216
rect 52552 18173 52561 18207
rect 52561 18173 52595 18207
rect 52595 18173 52604 18207
rect 52552 18164 52604 18173
rect 53840 18164 53892 18216
rect 56876 18164 56928 18216
rect 1860 18028 1912 18037
rect 4344 18028 4396 18080
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 6092 18028 6144 18080
rect 7932 18028 7984 18080
rect 8760 18028 8812 18080
rect 13912 18096 13964 18148
rect 20720 18096 20772 18148
rect 22008 18096 22060 18148
rect 26700 18096 26752 18148
rect 27160 18139 27212 18148
rect 27160 18105 27169 18139
rect 27169 18105 27203 18139
rect 27203 18105 27212 18139
rect 27160 18096 27212 18105
rect 46112 18096 46164 18148
rect 56508 18139 56560 18148
rect 56508 18105 56517 18139
rect 56517 18105 56551 18139
rect 56551 18105 56560 18139
rect 57704 18164 57756 18216
rect 56508 18096 56560 18105
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 12624 18028 12676 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 14924 18028 14976 18080
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 16396 18028 16448 18080
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 20904 18028 20956 18080
rect 25228 18028 25280 18080
rect 25964 18028 26016 18080
rect 37556 18071 37608 18080
rect 37556 18037 37565 18071
rect 37565 18037 37599 18071
rect 37599 18037 37608 18071
rect 37556 18028 37608 18037
rect 38752 18071 38804 18080
rect 38752 18037 38761 18071
rect 38761 18037 38795 18071
rect 38795 18037 38804 18071
rect 38752 18028 38804 18037
rect 40040 18028 40092 18080
rect 43168 18028 43220 18080
rect 43904 18028 43956 18080
rect 44088 18071 44140 18080
rect 44088 18037 44097 18071
rect 44097 18037 44131 18071
rect 44131 18037 44140 18071
rect 44088 18028 44140 18037
rect 44180 18028 44232 18080
rect 45376 18071 45428 18080
rect 45376 18037 45385 18071
rect 45385 18037 45419 18071
rect 45419 18037 45428 18071
rect 45376 18028 45428 18037
rect 47860 18071 47912 18080
rect 47860 18037 47869 18071
rect 47869 18037 47903 18071
rect 47903 18037 47912 18071
rect 47860 18028 47912 18037
rect 49332 18071 49384 18080
rect 49332 18037 49341 18071
rect 49341 18037 49375 18071
rect 49375 18037 49384 18071
rect 49332 18028 49384 18037
rect 51908 18071 51960 18080
rect 51908 18037 51917 18071
rect 51917 18037 51951 18071
rect 51951 18037 51960 18071
rect 51908 18028 51960 18037
rect 53380 18028 53432 18080
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 22616 17926 22668 17978
rect 22680 17926 22732 17978
rect 22744 17926 22796 17978
rect 22808 17926 22860 17978
rect 22872 17926 22924 17978
rect 37060 17926 37112 17978
rect 37124 17926 37176 17978
rect 37188 17926 37240 17978
rect 37252 17926 37304 17978
rect 37316 17926 37368 17978
rect 51504 17926 51556 17978
rect 51568 17926 51620 17978
rect 51632 17926 51684 17978
rect 51696 17926 51748 17978
rect 51760 17926 51812 17978
rect 3792 17867 3844 17876
rect 3792 17833 3801 17867
rect 3801 17833 3835 17867
rect 3835 17833 3844 17867
rect 3792 17824 3844 17833
rect 4712 17824 4764 17876
rect 8576 17824 8628 17876
rect 7564 17756 7616 17808
rect 9864 17824 9916 17876
rect 9956 17824 10008 17876
rect 12992 17824 13044 17876
rect 13912 17824 13964 17876
rect 14832 17824 14884 17876
rect 15200 17824 15252 17876
rect 13084 17756 13136 17808
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 5540 17731 5592 17740
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 7748 17688 7800 17740
rect 9036 17688 9088 17740
rect 12532 17688 12584 17740
rect 13544 17688 13596 17740
rect 6276 17552 6328 17604
rect 9496 17595 9548 17604
rect 9496 17561 9530 17595
rect 9530 17561 9548 17595
rect 9496 17552 9548 17561
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 8760 17484 8812 17536
rect 13820 17620 13872 17672
rect 25228 17867 25280 17876
rect 25228 17833 25237 17867
rect 25237 17833 25271 17867
rect 25271 17833 25280 17867
rect 25228 17824 25280 17833
rect 26056 17824 26108 17876
rect 48412 17824 48464 17876
rect 37556 17756 37608 17808
rect 17316 17688 17368 17740
rect 40040 17756 40092 17808
rect 15752 17620 15804 17672
rect 16764 17663 16816 17672
rect 16764 17629 16773 17663
rect 16773 17629 16807 17663
rect 16807 17629 16816 17663
rect 16764 17620 16816 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 18972 17663 19024 17672
rect 18972 17629 18981 17663
rect 18981 17629 19015 17663
rect 19015 17629 19024 17663
rect 18972 17620 19024 17629
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 21640 17663 21692 17672
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 26240 17620 26292 17672
rect 30380 17620 30432 17672
rect 30840 17663 30892 17672
rect 30840 17629 30849 17663
rect 30849 17629 30883 17663
rect 30883 17629 30892 17663
rect 30840 17620 30892 17629
rect 33048 17663 33100 17672
rect 33048 17629 33057 17663
rect 33057 17629 33091 17663
rect 33091 17629 33100 17663
rect 33048 17620 33100 17629
rect 33784 17663 33836 17672
rect 33784 17629 33793 17663
rect 33793 17629 33827 17663
rect 33827 17629 33836 17663
rect 33784 17620 33836 17629
rect 36360 17663 36412 17672
rect 36360 17629 36369 17663
rect 36369 17629 36403 17663
rect 36403 17629 36412 17663
rect 36360 17620 36412 17629
rect 36636 17663 36688 17672
rect 36636 17629 36645 17663
rect 36645 17629 36679 17663
rect 36679 17629 36688 17663
rect 36636 17620 36688 17629
rect 38752 17620 38804 17672
rect 18052 17552 18104 17604
rect 23388 17595 23440 17604
rect 23388 17561 23397 17595
rect 23397 17561 23431 17595
rect 23431 17561 23440 17595
rect 23388 17552 23440 17561
rect 37188 17595 37240 17604
rect 37188 17561 37197 17595
rect 37197 17561 37231 17595
rect 37231 17561 37240 17595
rect 37188 17552 37240 17561
rect 40408 17663 40460 17672
rect 40408 17629 40417 17663
rect 40417 17629 40451 17663
rect 40451 17629 40460 17663
rect 40408 17620 40460 17629
rect 41144 17663 41196 17672
rect 41144 17629 41153 17663
rect 41153 17629 41187 17663
rect 41187 17629 41196 17663
rect 41144 17620 41196 17629
rect 41328 17663 41380 17672
rect 41328 17629 41337 17663
rect 41337 17629 41371 17663
rect 41371 17629 41380 17663
rect 41328 17620 41380 17629
rect 40132 17552 40184 17604
rect 42432 17663 42484 17672
rect 42432 17629 42441 17663
rect 42441 17629 42475 17663
rect 42475 17629 42484 17663
rect 42432 17620 42484 17629
rect 45376 17688 45428 17740
rect 47768 17731 47820 17740
rect 47768 17697 47777 17731
rect 47777 17697 47811 17731
rect 47811 17697 47820 17731
rect 47768 17688 47820 17697
rect 48688 17799 48740 17808
rect 48688 17765 48697 17799
rect 48697 17765 48731 17799
rect 48731 17765 48740 17799
rect 48688 17756 48740 17765
rect 44824 17620 44876 17672
rect 47676 17620 47728 17672
rect 48964 17620 49016 17672
rect 50160 17756 50212 17808
rect 49240 17731 49292 17740
rect 49240 17697 49249 17731
rect 49249 17697 49283 17731
rect 49283 17697 49292 17731
rect 49240 17688 49292 17697
rect 52552 17824 52604 17876
rect 53840 17824 53892 17876
rect 57704 17867 57756 17876
rect 57704 17833 57713 17867
rect 57713 17833 57747 17867
rect 57747 17833 57756 17867
rect 57704 17824 57756 17833
rect 49148 17620 49200 17672
rect 51908 17620 51960 17672
rect 52552 17688 52604 17740
rect 56232 17688 56284 17740
rect 54484 17663 54536 17672
rect 54484 17629 54493 17663
rect 54493 17629 54527 17663
rect 54527 17629 54536 17663
rect 54484 17620 54536 17629
rect 56600 17663 56652 17672
rect 56600 17629 56634 17663
rect 56634 17629 56652 17663
rect 56600 17620 56652 17629
rect 43260 17552 43312 17604
rect 49332 17552 49384 17604
rect 55956 17552 56008 17604
rect 13912 17484 13964 17536
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 18512 17484 18564 17536
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 20812 17484 20864 17536
rect 25320 17527 25372 17536
rect 25320 17493 25329 17527
rect 25329 17493 25363 17527
rect 25363 17493 25372 17527
rect 25320 17484 25372 17493
rect 26332 17484 26384 17536
rect 29736 17484 29788 17536
rect 31208 17484 31260 17536
rect 33140 17484 33192 17536
rect 34428 17527 34480 17536
rect 34428 17493 34437 17527
rect 34437 17493 34471 17527
rect 34471 17493 34480 17527
rect 34428 17484 34480 17493
rect 35716 17484 35768 17536
rect 37372 17484 37424 17536
rect 38384 17484 38436 17536
rect 38568 17484 38620 17536
rect 39672 17527 39724 17536
rect 39672 17493 39681 17527
rect 39681 17493 39715 17527
rect 39715 17493 39724 17527
rect 39672 17484 39724 17493
rect 39856 17527 39908 17536
rect 39856 17493 39865 17527
rect 39865 17493 39899 17527
rect 39899 17493 39908 17527
rect 39856 17484 39908 17493
rect 40592 17527 40644 17536
rect 40592 17493 40601 17527
rect 40601 17493 40635 17527
rect 40635 17493 40644 17527
rect 40592 17484 40644 17493
rect 40684 17484 40736 17536
rect 44180 17484 44232 17536
rect 44732 17484 44784 17536
rect 45284 17484 45336 17536
rect 48320 17527 48372 17536
rect 48320 17493 48329 17527
rect 48329 17493 48363 17527
rect 48363 17493 48372 17527
rect 48320 17484 48372 17493
rect 49516 17484 49568 17536
rect 50252 17484 50304 17536
rect 51908 17484 51960 17536
rect 52092 17527 52144 17536
rect 52092 17493 52101 17527
rect 52101 17493 52135 17527
rect 52135 17493 52144 17527
rect 52092 17484 52144 17493
rect 54208 17484 54260 17536
rect 55220 17484 55272 17536
rect 56600 17484 56652 17536
rect 15394 17382 15446 17434
rect 15458 17382 15510 17434
rect 15522 17382 15574 17434
rect 15586 17382 15638 17434
rect 15650 17382 15702 17434
rect 29838 17382 29890 17434
rect 29902 17382 29954 17434
rect 29966 17382 30018 17434
rect 30030 17382 30082 17434
rect 30094 17382 30146 17434
rect 44282 17382 44334 17434
rect 44346 17382 44398 17434
rect 44410 17382 44462 17434
rect 44474 17382 44526 17434
rect 44538 17382 44590 17434
rect 58726 17382 58778 17434
rect 58790 17382 58842 17434
rect 58854 17382 58906 17434
rect 58918 17382 58970 17434
rect 58982 17382 59034 17434
rect 4344 17280 4396 17332
rect 4712 17280 4764 17332
rect 6920 17280 6972 17332
rect 8760 17280 8812 17332
rect 10140 17280 10192 17332
rect 14188 17280 14240 17332
rect 14280 17280 14332 17332
rect 16764 17280 16816 17332
rect 18236 17280 18288 17332
rect 18512 17323 18564 17332
rect 18512 17289 18521 17323
rect 18521 17289 18555 17323
rect 18555 17289 18564 17323
rect 18512 17280 18564 17289
rect 20168 17280 20220 17332
rect 20260 17280 20312 17332
rect 20812 17323 20864 17332
rect 20812 17289 20821 17323
rect 20821 17289 20855 17323
rect 20855 17289 20864 17323
rect 20812 17280 20864 17289
rect 20996 17280 21048 17332
rect 23848 17280 23900 17332
rect 24768 17280 24820 17332
rect 25872 17280 25924 17332
rect 27344 17323 27396 17332
rect 27344 17289 27353 17323
rect 27353 17289 27387 17323
rect 27387 17289 27396 17323
rect 27344 17280 27396 17289
rect 29736 17280 29788 17332
rect 30840 17280 30892 17332
rect 33784 17280 33836 17332
rect 34704 17280 34756 17332
rect 36360 17280 36412 17332
rect 36728 17280 36780 17332
rect 39856 17280 39908 17332
rect 40132 17323 40184 17332
rect 40132 17289 40141 17323
rect 40141 17289 40175 17323
rect 40175 17289 40184 17323
rect 40132 17280 40184 17289
rect 41144 17280 41196 17332
rect 9128 17212 9180 17264
rect 9496 17212 9548 17264
rect 9956 17212 10008 17264
rect 10232 17144 10284 17196
rect 12532 17212 12584 17264
rect 12624 17144 12676 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 15016 17212 15068 17264
rect 17316 17212 17368 17264
rect 13912 17144 13964 17153
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 4712 17051 4764 17060
rect 4712 17017 4721 17051
rect 4721 17017 4755 17051
rect 4755 17017 4764 17051
rect 4712 17008 4764 17017
rect 5264 17008 5316 17060
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 3424 16983 3476 16992
rect 3424 16949 3433 16983
rect 3433 16949 3467 16983
rect 3467 16949 3476 16983
rect 3424 16940 3476 16949
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 7564 17008 7616 17060
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 10416 17076 10468 17128
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 14280 17076 14332 17128
rect 16120 17144 16172 17196
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 19524 17212 19576 17264
rect 19800 17144 19852 17196
rect 20628 17144 20680 17196
rect 21548 17212 21600 17264
rect 25964 17212 26016 17264
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 22100 17187 22152 17196
rect 22100 17153 22123 17187
rect 22123 17153 22152 17187
rect 22100 17144 22152 17153
rect 25412 17144 25464 17196
rect 15936 17076 15988 17128
rect 16396 17076 16448 17128
rect 13360 17051 13412 17060
rect 13360 17017 13369 17051
rect 13369 17017 13403 17051
rect 13403 17017 13412 17051
rect 13360 17008 13412 17017
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 23388 17076 23440 17128
rect 24400 17119 24452 17128
rect 24400 17085 24409 17119
rect 24409 17085 24443 17119
rect 24443 17085 24452 17119
rect 24400 17076 24452 17085
rect 24768 17076 24820 17128
rect 26976 17144 27028 17196
rect 29552 17187 29604 17196
rect 29552 17153 29561 17187
rect 29561 17153 29595 17187
rect 29595 17153 29604 17187
rect 29552 17144 29604 17153
rect 30472 17212 30524 17264
rect 35808 17212 35860 17264
rect 33140 17187 33192 17196
rect 26056 17119 26108 17128
rect 26056 17085 26065 17119
rect 26065 17085 26099 17119
rect 26099 17085 26108 17119
rect 26056 17076 26108 17085
rect 26332 17076 26384 17128
rect 27436 17119 27488 17128
rect 27436 17085 27445 17119
rect 27445 17085 27479 17119
rect 27479 17085 27488 17119
rect 27436 17076 27488 17085
rect 24952 17008 25004 17060
rect 26792 17051 26844 17060
rect 26792 17017 26801 17051
rect 26801 17017 26835 17051
rect 26835 17017 26844 17051
rect 28816 17119 28868 17128
rect 28816 17085 28825 17119
rect 28825 17085 28859 17119
rect 28859 17085 28868 17119
rect 28816 17076 28868 17085
rect 29092 17076 29144 17128
rect 31576 17119 31628 17128
rect 31576 17085 31585 17119
rect 31585 17085 31619 17119
rect 31619 17085 31628 17119
rect 31576 17076 31628 17085
rect 26792 17008 26844 17017
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 16212 16940 16264 16992
rect 16580 16940 16632 16992
rect 18052 16940 18104 16992
rect 20996 16940 21048 16992
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 21548 16940 21600 16949
rect 23940 16940 23992 16992
rect 26884 16940 26936 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 31852 17008 31904 17060
rect 33140 17153 33149 17187
rect 33149 17153 33183 17187
rect 33183 17153 33192 17187
rect 33140 17144 33192 17153
rect 37188 17144 37240 17196
rect 37372 17144 37424 17196
rect 40684 17212 40736 17264
rect 42524 17280 42576 17332
rect 44640 17280 44692 17332
rect 45284 17280 45336 17332
rect 34244 17119 34296 17128
rect 34244 17085 34253 17119
rect 34253 17085 34287 17119
rect 34287 17085 34296 17119
rect 34244 17076 34296 17085
rect 34336 17076 34388 17128
rect 29460 16940 29512 16949
rect 30932 16940 30984 16992
rect 32680 16940 32732 16992
rect 34796 17008 34848 17060
rect 34060 16940 34112 16992
rect 34704 16983 34756 16992
rect 34704 16949 34713 16983
rect 34713 16949 34747 16983
rect 34747 16949 34756 16983
rect 34704 16940 34756 16949
rect 35256 16940 35308 16992
rect 35900 16940 35952 16992
rect 36268 16940 36320 16992
rect 36452 17119 36504 17128
rect 36452 17085 36461 17119
rect 36461 17085 36495 17119
rect 36495 17085 36504 17119
rect 36452 17076 36504 17085
rect 39212 17076 39264 17128
rect 39488 17119 39540 17128
rect 39488 17085 39497 17119
rect 39497 17085 39531 17119
rect 39531 17085 39540 17119
rect 39488 17076 39540 17085
rect 39672 17076 39724 17128
rect 37464 16940 37516 16992
rect 38660 16983 38712 16992
rect 38660 16949 38669 16983
rect 38669 16949 38703 16983
rect 38703 16949 38712 16983
rect 38660 16940 38712 16949
rect 39120 16940 39172 16992
rect 39396 16940 39448 16992
rect 39488 16940 39540 16992
rect 42800 17144 42852 17196
rect 45560 17187 45612 17196
rect 45560 17153 45569 17187
rect 45569 17153 45603 17187
rect 45603 17153 45612 17187
rect 45560 17144 45612 17153
rect 41512 17076 41564 17128
rect 44180 17076 44232 17128
rect 45376 17119 45428 17128
rect 45376 17085 45385 17119
rect 45385 17085 45419 17119
rect 45419 17085 45428 17119
rect 45376 17076 45428 17085
rect 43812 16940 43864 16992
rect 46020 16983 46072 16992
rect 46020 16949 46029 16983
rect 46029 16949 46063 16983
rect 46063 16949 46072 16983
rect 46020 16940 46072 16949
rect 48780 17280 48832 17332
rect 47860 17255 47912 17264
rect 47860 17221 47894 17255
rect 47894 17221 47912 17255
rect 47860 17212 47912 17221
rect 48596 17212 48648 17264
rect 49240 17212 49292 17264
rect 49516 17212 49568 17264
rect 52092 17280 52144 17332
rect 52460 17280 52512 17332
rect 47676 17144 47728 17196
rect 50160 17187 50212 17196
rect 50160 17153 50169 17187
rect 50169 17153 50203 17187
rect 50203 17153 50212 17187
rect 50160 17144 50212 17153
rect 50436 17187 50488 17196
rect 50436 17153 50445 17187
rect 50445 17153 50479 17187
rect 50479 17153 50488 17187
rect 50436 17144 50488 17153
rect 51172 17187 51224 17196
rect 51172 17153 51181 17187
rect 51181 17153 51215 17187
rect 51215 17153 51224 17187
rect 51172 17144 51224 17153
rect 54484 17323 54536 17332
rect 54484 17289 54493 17323
rect 54493 17289 54527 17323
rect 54527 17289 54536 17323
rect 54484 17280 54536 17289
rect 56508 17280 56560 17332
rect 54944 17255 54996 17264
rect 54944 17221 54953 17255
rect 54953 17221 54987 17255
rect 54987 17221 54996 17255
rect 54944 17212 54996 17221
rect 55220 17212 55272 17264
rect 47032 17076 47084 17128
rect 49332 17076 49384 17128
rect 50620 17076 50672 17128
rect 53380 17187 53432 17196
rect 53380 17153 53414 17187
rect 53414 17153 53432 17187
rect 53380 17144 53432 17153
rect 54116 17144 54168 17196
rect 55956 17144 56008 17196
rect 56968 17144 57020 17196
rect 51356 17008 51408 17060
rect 51908 17076 51960 17128
rect 52184 17076 52236 17128
rect 55496 17076 55548 17128
rect 56324 17076 56376 17128
rect 56508 17076 56560 17128
rect 57060 17119 57112 17128
rect 57060 17085 57069 17119
rect 57069 17085 57103 17119
rect 57103 17085 57112 17119
rect 57060 17076 57112 17085
rect 48780 16940 48832 16992
rect 50252 16940 50304 16992
rect 52552 16983 52604 16992
rect 52552 16949 52561 16983
rect 52561 16949 52595 16983
rect 52595 16949 52604 16983
rect 55404 17008 55456 17060
rect 52552 16940 52604 16949
rect 56508 16940 56560 16992
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 22616 16838 22668 16890
rect 22680 16838 22732 16890
rect 22744 16838 22796 16890
rect 22808 16838 22860 16890
rect 22872 16838 22924 16890
rect 37060 16838 37112 16890
rect 37124 16838 37176 16890
rect 37188 16838 37240 16890
rect 37252 16838 37304 16890
rect 37316 16838 37368 16890
rect 51504 16838 51556 16890
rect 51568 16838 51620 16890
rect 51632 16838 51684 16890
rect 51696 16838 51748 16890
rect 51760 16838 51812 16890
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 6736 16736 6788 16788
rect 7380 16736 7432 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 4160 16600 4212 16652
rect 4712 16600 4764 16652
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 10692 16643 10744 16652
rect 10692 16609 10701 16643
rect 10701 16609 10735 16643
rect 10735 16609 10744 16643
rect 10692 16600 10744 16609
rect 10784 16600 10836 16652
rect 12532 16736 12584 16788
rect 16028 16736 16080 16788
rect 18972 16736 19024 16788
rect 19708 16736 19760 16788
rect 20812 16736 20864 16788
rect 21824 16736 21876 16788
rect 22560 16736 22612 16788
rect 26240 16779 26292 16788
rect 26240 16745 26249 16779
rect 26249 16745 26283 16779
rect 26283 16745 26292 16779
rect 26240 16736 26292 16745
rect 14096 16600 14148 16652
rect 14924 16643 14976 16652
rect 14924 16609 14942 16643
rect 14942 16609 14976 16643
rect 14924 16600 14976 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 19064 16668 19116 16720
rect 17316 16600 17368 16652
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 20444 16643 20496 16652
rect 20444 16609 20453 16643
rect 20453 16609 20487 16643
rect 20487 16609 20496 16643
rect 20444 16600 20496 16609
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 10324 16532 10376 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 17684 16575 17736 16584
rect 15752 16532 15804 16541
rect 4896 16464 4948 16516
rect 12808 16464 12860 16516
rect 17684 16541 17718 16575
rect 17718 16541 17736 16575
rect 17684 16532 17736 16541
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 19892 16532 19944 16541
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 25964 16600 26016 16652
rect 26240 16600 26292 16652
rect 26976 16736 27028 16788
rect 29644 16736 29696 16788
rect 30104 16736 30156 16788
rect 30656 16736 30708 16788
rect 30932 16736 30984 16788
rect 28448 16643 28500 16652
rect 28448 16609 28457 16643
rect 28457 16609 28491 16643
rect 28491 16609 28500 16643
rect 28448 16600 28500 16609
rect 30104 16643 30156 16652
rect 30104 16609 30113 16643
rect 30113 16609 30147 16643
rect 30147 16609 30156 16643
rect 30104 16600 30156 16609
rect 32680 16736 32732 16788
rect 33048 16736 33100 16788
rect 33876 16736 33928 16788
rect 31208 16600 31260 16652
rect 31484 16643 31536 16652
rect 31484 16609 31493 16643
rect 31493 16609 31527 16643
rect 31527 16609 31536 16643
rect 31484 16600 31536 16609
rect 31852 16643 31904 16652
rect 31852 16609 31886 16643
rect 31886 16609 31904 16643
rect 31852 16600 31904 16609
rect 32680 16643 32732 16652
rect 32680 16609 32689 16643
rect 32689 16609 32723 16643
rect 32723 16609 32732 16643
rect 32680 16600 32732 16609
rect 34336 16736 34388 16788
rect 36636 16736 36688 16788
rect 37556 16736 37608 16788
rect 38936 16736 38988 16788
rect 39212 16736 39264 16788
rect 39028 16711 39080 16720
rect 39028 16677 39037 16711
rect 39037 16677 39071 16711
rect 39071 16677 39080 16711
rect 39028 16668 39080 16677
rect 39856 16668 39908 16720
rect 36728 16600 36780 16652
rect 37464 16600 37516 16652
rect 38292 16600 38344 16652
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 11428 16396 11480 16448
rect 13268 16439 13320 16448
rect 13268 16405 13277 16439
rect 13277 16405 13311 16439
rect 13311 16405 13320 16439
rect 13268 16396 13320 16405
rect 15200 16396 15252 16448
rect 19616 16396 19668 16448
rect 23940 16575 23992 16584
rect 23940 16541 23949 16575
rect 23949 16541 23983 16575
rect 23983 16541 23992 16575
rect 23940 16532 23992 16541
rect 26884 16575 26936 16584
rect 26884 16541 26918 16575
rect 26918 16541 26936 16575
rect 26884 16532 26936 16541
rect 29460 16532 29512 16584
rect 20996 16464 21048 16516
rect 25320 16464 25372 16516
rect 30472 16532 30524 16584
rect 32036 16575 32088 16584
rect 32036 16541 32045 16575
rect 32045 16541 32079 16575
rect 32079 16541 32088 16575
rect 32036 16532 32088 16541
rect 34428 16532 34480 16584
rect 39488 16643 39540 16652
rect 39488 16609 39497 16643
rect 39497 16609 39531 16643
rect 39531 16609 39540 16643
rect 39488 16600 39540 16609
rect 42432 16736 42484 16788
rect 43812 16736 43864 16788
rect 44824 16711 44876 16720
rect 44824 16677 44833 16711
rect 44833 16677 44867 16711
rect 44867 16677 44876 16711
rect 44824 16668 44876 16677
rect 47676 16736 47728 16788
rect 48780 16736 48832 16788
rect 51356 16779 51408 16788
rect 51356 16745 51365 16779
rect 51365 16745 51399 16779
rect 51399 16745 51408 16779
rect 51356 16736 51408 16745
rect 48688 16600 48740 16652
rect 35716 16507 35768 16516
rect 35716 16473 35750 16507
rect 35750 16473 35768 16507
rect 35716 16464 35768 16473
rect 35808 16464 35860 16516
rect 38568 16532 38620 16584
rect 38752 16575 38804 16584
rect 38752 16541 38761 16575
rect 38761 16541 38795 16575
rect 38795 16541 38804 16575
rect 38752 16532 38804 16541
rect 40408 16532 40460 16584
rect 41328 16532 41380 16584
rect 44088 16532 44140 16584
rect 46020 16532 46072 16584
rect 47032 16532 47084 16584
rect 48136 16532 48188 16584
rect 50068 16668 50120 16720
rect 50712 16600 50764 16652
rect 52368 16600 52420 16652
rect 54116 16736 54168 16788
rect 55496 16736 55548 16788
rect 56140 16643 56192 16652
rect 56140 16609 56149 16643
rect 56149 16609 56183 16643
rect 56183 16609 56192 16643
rect 56140 16600 56192 16609
rect 57152 16600 57204 16652
rect 55864 16575 55916 16584
rect 55864 16541 55873 16575
rect 55873 16541 55907 16575
rect 55907 16541 55916 16575
rect 55864 16532 55916 16541
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 24768 16396 24820 16448
rect 27988 16439 28040 16448
rect 27988 16405 27997 16439
rect 27997 16405 28031 16439
rect 28031 16405 28040 16439
rect 27988 16396 28040 16405
rect 28632 16439 28684 16448
rect 28632 16405 28641 16439
rect 28641 16405 28675 16439
rect 28675 16405 28684 16439
rect 28632 16396 28684 16405
rect 30748 16439 30800 16448
rect 30748 16405 30757 16439
rect 30757 16405 30791 16439
rect 30791 16405 30800 16439
rect 30748 16396 30800 16405
rect 37648 16439 37700 16448
rect 37648 16405 37657 16439
rect 37657 16405 37691 16439
rect 37691 16405 37700 16439
rect 37648 16396 37700 16405
rect 38752 16396 38804 16448
rect 41604 16464 41656 16516
rect 43076 16439 43128 16448
rect 43076 16405 43085 16439
rect 43085 16405 43119 16439
rect 43119 16405 43128 16439
rect 43076 16396 43128 16405
rect 48688 16439 48740 16448
rect 48688 16405 48697 16439
rect 48697 16405 48731 16439
rect 48731 16405 48740 16439
rect 48688 16396 48740 16405
rect 52092 16439 52144 16448
rect 52092 16405 52101 16439
rect 52101 16405 52135 16439
rect 52135 16405 52144 16439
rect 52092 16396 52144 16405
rect 54760 16439 54812 16448
rect 54760 16405 54769 16439
rect 54769 16405 54803 16439
rect 54803 16405 54812 16439
rect 54760 16396 54812 16405
rect 57520 16439 57572 16448
rect 57520 16405 57529 16439
rect 57529 16405 57563 16439
rect 57563 16405 57572 16439
rect 57520 16396 57572 16405
rect 15394 16294 15446 16346
rect 15458 16294 15510 16346
rect 15522 16294 15574 16346
rect 15586 16294 15638 16346
rect 15650 16294 15702 16346
rect 29838 16294 29890 16346
rect 29902 16294 29954 16346
rect 29966 16294 30018 16346
rect 30030 16294 30082 16346
rect 30094 16294 30146 16346
rect 44282 16294 44334 16346
rect 44346 16294 44398 16346
rect 44410 16294 44462 16346
rect 44474 16294 44526 16346
rect 44538 16294 44590 16346
rect 58726 16294 58778 16346
rect 58790 16294 58842 16346
rect 58854 16294 58906 16346
rect 58918 16294 58970 16346
rect 58982 16294 59034 16346
rect 2964 16192 3016 16244
rect 3976 16192 4028 16244
rect 4160 16192 4212 16244
rect 4436 16192 4488 16244
rect 9312 16192 9364 16244
rect 12808 16235 12860 16244
rect 12808 16201 12817 16235
rect 12817 16201 12851 16235
rect 12851 16201 12860 16235
rect 12808 16192 12860 16201
rect 13268 16192 13320 16244
rect 13820 16192 13872 16244
rect 14924 16192 14976 16244
rect 15108 16235 15160 16244
rect 15108 16201 15117 16235
rect 15117 16201 15151 16235
rect 15151 16201 15160 16235
rect 15108 16192 15160 16201
rect 15752 16192 15804 16244
rect 16120 16192 16172 16244
rect 17316 16192 17368 16244
rect 19156 16192 19208 16244
rect 19616 16192 19668 16244
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 13176 16056 13228 16108
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 18420 16124 18472 16176
rect 20628 16192 20680 16244
rect 21640 16192 21692 16244
rect 22100 16192 22152 16244
rect 22192 16235 22244 16244
rect 22192 16201 22201 16235
rect 22201 16201 22235 16235
rect 22235 16201 22244 16235
rect 22192 16192 22244 16201
rect 23388 16192 23440 16244
rect 24400 16192 24452 16244
rect 20352 16124 20404 16176
rect 17592 16056 17644 16108
rect 19524 16056 19576 16108
rect 25320 16192 25372 16244
rect 26792 16192 26844 16244
rect 27252 16235 27304 16244
rect 27252 16201 27261 16235
rect 27261 16201 27295 16235
rect 27295 16201 27304 16235
rect 27252 16192 27304 16201
rect 28816 16192 28868 16244
rect 29552 16192 29604 16244
rect 31576 16192 31628 16244
rect 32036 16192 32088 16244
rect 37648 16192 37700 16244
rect 38752 16192 38804 16244
rect 41512 16192 41564 16244
rect 41604 16235 41656 16244
rect 41604 16201 41613 16235
rect 41613 16201 41647 16235
rect 41647 16201 41656 16235
rect 41604 16192 41656 16201
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 4344 16031 4396 16040
rect 4344 15997 4353 16031
rect 4353 15997 4387 16031
rect 4387 15997 4396 16031
rect 4344 15988 4396 15997
rect 4620 15988 4672 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 7840 15988 7892 16040
rect 14464 15988 14516 16040
rect 19616 16031 19668 16040
rect 19616 15997 19625 16031
rect 19625 15997 19659 16031
rect 19659 15997 19668 16031
rect 19616 15988 19668 15997
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 26332 16099 26384 16108
rect 26332 16065 26341 16099
rect 26341 16065 26375 16099
rect 26375 16065 26384 16099
rect 26332 16056 26384 16065
rect 26700 16099 26752 16108
rect 26700 16065 26709 16099
rect 26709 16065 26743 16099
rect 26743 16065 26752 16099
rect 26700 16056 26752 16065
rect 29368 16056 29420 16108
rect 34704 16124 34756 16176
rect 30840 16056 30892 16108
rect 35808 16056 35860 16108
rect 40592 16124 40644 16176
rect 42340 16124 42392 16176
rect 39212 16056 39264 16108
rect 42984 16056 43036 16108
rect 22560 15988 22612 16040
rect 24768 15988 24820 16040
rect 25228 15988 25280 16040
rect 27620 15988 27672 16040
rect 25688 15963 25740 15972
rect 25688 15929 25697 15963
rect 25697 15929 25731 15963
rect 25731 15929 25740 15963
rect 25688 15920 25740 15929
rect 47768 16192 47820 16244
rect 48688 16192 48740 16244
rect 50344 16192 50396 16244
rect 51264 16192 51316 16244
rect 56324 16192 56376 16244
rect 57152 16235 57204 16244
rect 57152 16201 57161 16235
rect 57161 16201 57195 16235
rect 57195 16201 57204 16235
rect 57152 16192 57204 16201
rect 57520 16192 57572 16244
rect 44272 16056 44324 16108
rect 45284 16056 45336 16108
rect 45560 16056 45612 16108
rect 47216 16056 47268 16108
rect 54760 16124 54812 16176
rect 49700 16099 49752 16108
rect 49700 16065 49709 16099
rect 49709 16065 49743 16099
rect 49743 16065 49752 16099
rect 49700 16056 49752 16065
rect 52000 16099 52052 16108
rect 52000 16065 52009 16099
rect 52009 16065 52043 16099
rect 52043 16065 52052 16099
rect 52000 16056 52052 16065
rect 56876 16056 56928 16108
rect 44180 16031 44232 16040
rect 44180 15997 44189 16031
rect 44189 15997 44223 16031
rect 44223 15997 44232 16031
rect 44180 15988 44232 15997
rect 44640 15988 44692 16040
rect 49516 15988 49568 16040
rect 50620 15988 50672 16040
rect 44824 15920 44876 15972
rect 46388 15920 46440 15972
rect 54208 16031 54260 16040
rect 54208 15997 54217 16031
rect 54217 15997 54251 16031
rect 54251 15997 54260 16031
rect 54208 15988 54260 15997
rect 55864 15988 55916 16040
rect 4068 15852 4120 15904
rect 6552 15852 6604 15904
rect 10692 15852 10744 15904
rect 14924 15852 14976 15904
rect 15292 15852 15344 15904
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 18972 15895 19024 15904
rect 18972 15861 18981 15895
rect 18981 15861 19015 15895
rect 19015 15861 19024 15895
rect 18972 15852 19024 15861
rect 19892 15852 19944 15904
rect 25964 15852 26016 15904
rect 27712 15895 27764 15904
rect 27712 15861 27721 15895
rect 27721 15861 27755 15895
rect 27755 15861 27764 15895
rect 27712 15852 27764 15861
rect 33140 15895 33192 15904
rect 33140 15861 33149 15895
rect 33149 15861 33183 15895
rect 33183 15861 33192 15895
rect 33140 15852 33192 15861
rect 34520 15852 34572 15904
rect 42800 15852 42852 15904
rect 45284 15852 45336 15904
rect 47124 15852 47176 15904
rect 48596 15852 48648 15904
rect 50344 15895 50396 15904
rect 50344 15861 50353 15895
rect 50353 15861 50387 15895
rect 50387 15861 50396 15895
rect 50344 15852 50396 15861
rect 50436 15895 50488 15904
rect 50436 15861 50445 15895
rect 50445 15861 50479 15895
rect 50479 15861 50488 15895
rect 50436 15852 50488 15861
rect 51356 15895 51408 15904
rect 51356 15861 51365 15895
rect 51365 15861 51399 15895
rect 51399 15861 51408 15895
rect 51356 15852 51408 15861
rect 55680 15852 55732 15904
rect 57060 15988 57112 16040
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 22616 15750 22668 15802
rect 22680 15750 22732 15802
rect 22744 15750 22796 15802
rect 22808 15750 22860 15802
rect 22872 15750 22924 15802
rect 37060 15750 37112 15802
rect 37124 15750 37176 15802
rect 37188 15750 37240 15802
rect 37252 15750 37304 15802
rect 37316 15750 37368 15802
rect 51504 15750 51556 15802
rect 51568 15750 51620 15802
rect 51632 15750 51684 15802
rect 51696 15750 51748 15802
rect 51760 15750 51812 15802
rect 4160 15648 4212 15700
rect 7840 15648 7892 15700
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 54024 15648 54076 15700
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 4896 15555 4948 15564
rect 4896 15521 4930 15555
rect 4930 15521 4948 15555
rect 4896 15512 4948 15521
rect 5264 15512 5316 15564
rect 6092 15512 6144 15564
rect 6460 15580 6512 15632
rect 6736 15580 6788 15632
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 2688 15444 2740 15496
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 7012 15512 7064 15564
rect 2136 15376 2188 15428
rect 4344 15308 4396 15360
rect 4436 15308 4488 15360
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 10416 15580 10468 15632
rect 13176 15580 13228 15632
rect 7656 15512 7708 15521
rect 7104 15376 7156 15428
rect 7196 15376 7248 15428
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 6920 15308 6972 15360
rect 16672 15512 16724 15564
rect 18512 15512 18564 15564
rect 22468 15512 22520 15564
rect 27620 15580 27672 15632
rect 27712 15580 27764 15632
rect 30380 15580 30432 15632
rect 30748 15580 30800 15632
rect 30840 15580 30892 15632
rect 31944 15623 31996 15632
rect 24860 15512 24912 15564
rect 28724 15555 28776 15564
rect 28724 15521 28733 15555
rect 28733 15521 28767 15555
rect 28767 15521 28776 15555
rect 28724 15512 28776 15521
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 19064 15444 19116 15496
rect 30472 15487 30524 15496
rect 30472 15453 30481 15487
rect 30481 15453 30515 15487
rect 30515 15453 30524 15487
rect 30472 15444 30524 15453
rect 30748 15444 30800 15496
rect 31944 15589 31953 15623
rect 31953 15589 31987 15623
rect 31987 15589 31996 15623
rect 31944 15580 31996 15589
rect 42340 15623 42392 15632
rect 42340 15589 42349 15623
rect 42349 15589 42383 15623
rect 42383 15589 42392 15623
rect 42340 15580 42392 15589
rect 42156 15512 42208 15564
rect 42616 15555 42668 15564
rect 42616 15521 42625 15555
rect 42625 15521 42659 15555
rect 42659 15521 42668 15555
rect 42616 15512 42668 15521
rect 43260 15623 43312 15632
rect 43260 15589 43269 15623
rect 43269 15589 43303 15623
rect 43303 15589 43312 15623
rect 43260 15580 43312 15589
rect 44824 15580 44876 15632
rect 44180 15512 44232 15564
rect 47584 15512 47636 15564
rect 48136 15580 48188 15632
rect 48044 15555 48096 15564
rect 48044 15521 48053 15555
rect 48053 15521 48087 15555
rect 48087 15521 48096 15555
rect 48044 15512 48096 15521
rect 37832 15444 37884 15496
rect 18328 15376 18380 15428
rect 20444 15376 20496 15428
rect 23204 15376 23256 15428
rect 31208 15376 31260 15428
rect 44640 15444 44692 15496
rect 48228 15487 48280 15496
rect 48228 15453 48237 15487
rect 48237 15453 48271 15487
rect 48271 15453 48280 15487
rect 48228 15444 48280 15453
rect 50252 15444 50304 15496
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 8116 15351 8168 15360
rect 8116 15317 8125 15351
rect 8125 15317 8159 15351
rect 8159 15317 8168 15351
rect 8116 15308 8168 15317
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 11980 15351 12032 15360
rect 11980 15317 11989 15351
rect 11989 15317 12023 15351
rect 12023 15317 12032 15351
rect 11980 15308 12032 15317
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 15016 15308 15068 15360
rect 17224 15308 17276 15360
rect 17960 15308 18012 15360
rect 19156 15308 19208 15360
rect 19616 15308 19668 15360
rect 20352 15308 20404 15360
rect 20904 15308 20956 15360
rect 25044 15351 25096 15360
rect 25044 15317 25053 15351
rect 25053 15317 25087 15351
rect 25087 15317 25096 15351
rect 25044 15308 25096 15317
rect 29276 15308 29328 15360
rect 38292 15308 38344 15360
rect 42800 15308 42852 15360
rect 49608 15376 49660 15428
rect 50068 15376 50120 15428
rect 51264 15512 51316 15564
rect 51908 15512 51960 15564
rect 52092 15444 52144 15496
rect 53472 15444 53524 15496
rect 57152 15512 57204 15564
rect 54116 15487 54168 15496
rect 54116 15453 54125 15487
rect 54125 15453 54159 15487
rect 54159 15453 54168 15487
rect 54116 15444 54168 15453
rect 54852 15487 54904 15496
rect 54852 15453 54861 15487
rect 54861 15453 54895 15487
rect 54895 15453 54904 15487
rect 54852 15444 54904 15453
rect 55220 15444 55272 15496
rect 48596 15308 48648 15360
rect 48688 15351 48740 15360
rect 48688 15317 48697 15351
rect 48697 15317 48731 15351
rect 48731 15317 48740 15351
rect 48688 15308 48740 15317
rect 49884 15308 49936 15360
rect 55036 15376 55088 15428
rect 55128 15376 55180 15428
rect 51264 15308 51316 15360
rect 51816 15308 51868 15360
rect 52184 15308 52236 15360
rect 52460 15351 52512 15360
rect 52460 15317 52469 15351
rect 52469 15317 52503 15351
rect 52503 15317 52512 15351
rect 52460 15308 52512 15317
rect 53380 15308 53432 15360
rect 54300 15351 54352 15360
rect 54300 15317 54309 15351
rect 54309 15317 54343 15351
rect 54343 15317 54352 15351
rect 54300 15308 54352 15317
rect 56232 15308 56284 15360
rect 56784 15351 56836 15360
rect 56784 15317 56793 15351
rect 56793 15317 56827 15351
rect 56827 15317 56836 15351
rect 56784 15308 56836 15317
rect 56876 15351 56928 15360
rect 56876 15317 56885 15351
rect 56885 15317 56919 15351
rect 56919 15317 56928 15351
rect 56876 15308 56928 15317
rect 57336 15351 57388 15360
rect 57336 15317 57345 15351
rect 57345 15317 57379 15351
rect 57379 15317 57388 15351
rect 57336 15308 57388 15317
rect 15394 15206 15446 15258
rect 15458 15206 15510 15258
rect 15522 15206 15574 15258
rect 15586 15206 15638 15258
rect 15650 15206 15702 15258
rect 29838 15206 29890 15258
rect 29902 15206 29954 15258
rect 29966 15206 30018 15258
rect 30030 15206 30082 15258
rect 30094 15206 30146 15258
rect 44282 15206 44334 15258
rect 44346 15206 44398 15258
rect 44410 15206 44462 15258
rect 44474 15206 44526 15258
rect 44538 15206 44590 15258
rect 58726 15206 58778 15258
rect 58790 15206 58842 15258
rect 58854 15206 58906 15258
rect 58918 15206 58970 15258
rect 58982 15206 59034 15258
rect 2136 15147 2188 15156
rect 2136 15113 2145 15147
rect 2145 15113 2179 15147
rect 2179 15113 2188 15147
rect 2136 15104 2188 15113
rect 5080 15104 5132 15156
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 6736 15147 6788 15156
rect 6736 15113 6745 15147
rect 6745 15113 6779 15147
rect 6779 15113 6788 15147
rect 6736 15104 6788 15113
rect 7472 15104 7524 15156
rect 7840 15104 7892 15156
rect 9128 15104 9180 15156
rect 12532 15104 12584 15156
rect 13912 15104 13964 15156
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 14648 15104 14700 15156
rect 2688 15036 2740 15088
rect 3424 15036 3476 15088
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 7196 14968 7248 15020
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 7012 14900 7064 14952
rect 8116 15036 8168 15088
rect 8484 15036 8536 15088
rect 12440 15036 12492 15088
rect 7472 14968 7524 15020
rect 7564 14900 7616 14952
rect 13452 14968 13504 15020
rect 9220 14832 9272 14884
rect 10416 14900 10468 14952
rect 10968 14900 11020 14952
rect 12440 14832 12492 14884
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 17592 15147 17644 15156
rect 17592 15113 17601 15147
rect 17601 15113 17635 15147
rect 17635 15113 17644 15147
rect 17592 15104 17644 15113
rect 19064 15104 19116 15156
rect 25044 15104 25096 15156
rect 25688 15104 25740 15156
rect 29368 15147 29420 15156
rect 29368 15113 29377 15147
rect 29377 15113 29411 15147
rect 29411 15113 29420 15147
rect 29368 15104 29420 15113
rect 30104 15147 30156 15156
rect 30104 15113 30113 15147
rect 30113 15113 30147 15147
rect 30147 15113 30156 15147
rect 30104 15104 30156 15113
rect 32312 15104 32364 15156
rect 36728 15104 36780 15156
rect 37556 15104 37608 15156
rect 42984 15104 43036 15156
rect 44088 15104 44140 15156
rect 49608 15104 49660 15156
rect 50620 15147 50672 15156
rect 50620 15113 50629 15147
rect 50629 15113 50663 15147
rect 50663 15113 50672 15147
rect 50620 15104 50672 15113
rect 50712 15147 50764 15156
rect 50712 15113 50721 15147
rect 50721 15113 50755 15147
rect 50755 15113 50764 15147
rect 50712 15104 50764 15113
rect 23848 15079 23900 15088
rect 23848 15045 23857 15079
rect 23857 15045 23891 15079
rect 23891 15045 23900 15079
rect 23848 15036 23900 15045
rect 24216 15036 24268 15088
rect 30472 15036 30524 15088
rect 31484 15036 31536 15088
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 15292 15011 15344 15020
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 17960 14968 18012 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 18512 14968 18564 15020
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 17776 14900 17828 14952
rect 21456 14900 21508 14952
rect 28448 14968 28500 15020
rect 28632 14968 28684 15020
rect 30196 15011 30248 15020
rect 30196 14977 30205 15011
rect 30205 14977 30239 15011
rect 30239 14977 30248 15011
rect 30196 14968 30248 14977
rect 4804 14764 4856 14816
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6920 14764 6972 14816
rect 8024 14764 8076 14816
rect 8116 14764 8168 14816
rect 9864 14764 9916 14816
rect 10324 14764 10376 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 14924 14832 14976 14884
rect 15200 14832 15252 14884
rect 15660 14875 15712 14884
rect 15660 14841 15669 14875
rect 15669 14841 15703 14875
rect 15703 14841 15712 14875
rect 15660 14832 15712 14841
rect 18052 14832 18104 14884
rect 19248 14832 19300 14884
rect 15844 14764 15896 14816
rect 23388 14807 23440 14816
rect 23388 14773 23397 14807
rect 23397 14773 23431 14807
rect 23431 14773 23440 14807
rect 23388 14764 23440 14773
rect 31484 14807 31536 14816
rect 31484 14773 31493 14807
rect 31493 14773 31527 14807
rect 31527 14773 31536 14807
rect 31484 14764 31536 14773
rect 36544 15036 36596 15088
rect 48688 15036 48740 15088
rect 52184 15104 52236 15156
rect 54116 15104 54168 15156
rect 54852 15104 54904 15156
rect 55036 15104 55088 15156
rect 57796 15104 57848 15156
rect 43076 15011 43128 15020
rect 43076 14977 43085 15011
rect 43085 14977 43119 15011
rect 43119 14977 43128 15011
rect 43076 14968 43128 14977
rect 47676 14968 47728 15020
rect 48412 14968 48464 15020
rect 49332 14968 49384 15020
rect 52460 15036 52512 15088
rect 54208 15036 54260 15088
rect 56232 15036 56284 15088
rect 57336 15036 57388 15088
rect 52368 14968 52420 15020
rect 33140 14832 33192 14884
rect 35624 14900 35676 14952
rect 35992 14900 36044 14952
rect 43352 14900 43404 14952
rect 38108 14832 38160 14884
rect 50068 14943 50120 14952
rect 50068 14909 50077 14943
rect 50077 14909 50111 14943
rect 50111 14909 50120 14943
rect 50068 14900 50120 14909
rect 50896 14900 50948 14952
rect 49608 14832 49660 14884
rect 51080 14832 51132 14884
rect 52092 14832 52144 14884
rect 52368 14832 52420 14884
rect 55128 14968 55180 15020
rect 56140 14968 56192 15020
rect 57612 14968 57664 15020
rect 54208 14943 54260 14952
rect 54208 14909 54217 14943
rect 54217 14909 54251 14943
rect 54251 14909 54260 14943
rect 54208 14900 54260 14909
rect 55036 14943 55088 14952
rect 55036 14909 55045 14943
rect 55045 14909 55079 14943
rect 55079 14909 55088 14943
rect 55036 14900 55088 14909
rect 55312 14943 55364 14952
rect 55312 14909 55321 14943
rect 55321 14909 55355 14943
rect 55355 14909 55364 14943
rect 55312 14900 55364 14909
rect 56048 14832 56100 14884
rect 32772 14764 32824 14816
rect 33232 14764 33284 14816
rect 33600 14807 33652 14816
rect 33600 14773 33609 14807
rect 33609 14773 33643 14807
rect 33643 14773 33652 14807
rect 33600 14764 33652 14773
rect 37740 14764 37792 14816
rect 38200 14764 38252 14816
rect 41788 14807 41840 14816
rect 41788 14773 41797 14807
rect 41797 14773 41831 14807
rect 41831 14773 41840 14807
rect 41788 14764 41840 14773
rect 42432 14764 42484 14816
rect 43812 14764 43864 14816
rect 45008 14807 45060 14816
rect 45008 14773 45017 14807
rect 45017 14773 45051 14807
rect 45051 14773 45060 14807
rect 45008 14764 45060 14773
rect 45376 14807 45428 14816
rect 45376 14773 45385 14807
rect 45385 14773 45419 14807
rect 45419 14773 45428 14807
rect 45376 14764 45428 14773
rect 49516 14764 49568 14816
rect 53840 14764 53892 14816
rect 54208 14764 54260 14816
rect 57704 14807 57756 14816
rect 57704 14773 57713 14807
rect 57713 14773 57747 14807
rect 57747 14773 57756 14807
rect 57704 14764 57756 14773
rect 58532 14807 58584 14816
rect 58532 14773 58541 14807
rect 58541 14773 58575 14807
rect 58575 14773 58584 14807
rect 58532 14764 58584 14773
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 22616 14662 22668 14714
rect 22680 14662 22732 14714
rect 22744 14662 22796 14714
rect 22808 14662 22860 14714
rect 22872 14662 22924 14714
rect 37060 14662 37112 14714
rect 37124 14662 37176 14714
rect 37188 14662 37240 14714
rect 37252 14662 37304 14714
rect 37316 14662 37368 14714
rect 51504 14662 51556 14714
rect 51568 14662 51620 14714
rect 51632 14662 51684 14714
rect 51696 14662 51748 14714
rect 51760 14662 51812 14714
rect 2780 14560 2832 14612
rect 5356 14560 5408 14612
rect 4252 14424 4304 14476
rect 7564 14560 7616 14612
rect 8024 14560 8076 14612
rect 9680 14560 9732 14612
rect 10508 14560 10560 14612
rect 12440 14560 12492 14612
rect 13176 14560 13228 14612
rect 15292 14560 15344 14612
rect 23204 14603 23256 14612
rect 23204 14569 23213 14603
rect 23213 14569 23247 14603
rect 23247 14569 23256 14603
rect 23204 14560 23256 14569
rect 23388 14560 23440 14612
rect 23572 14560 23624 14612
rect 24216 14603 24268 14612
rect 24216 14569 24225 14603
rect 24225 14569 24259 14603
rect 24259 14569 24268 14603
rect 24216 14560 24268 14569
rect 26056 14560 26108 14612
rect 29736 14560 29788 14612
rect 30104 14560 30156 14612
rect 35532 14560 35584 14612
rect 8760 14492 8812 14544
rect 9220 14492 9272 14544
rect 7196 14424 7248 14476
rect 8024 14424 8076 14476
rect 9128 14424 9180 14476
rect 4988 14356 5040 14408
rect 6000 14356 6052 14408
rect 7748 14399 7800 14408
rect 7748 14365 7766 14399
rect 7766 14365 7800 14399
rect 7748 14356 7800 14365
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8852 14356 8904 14408
rect 4436 14288 4488 14340
rect 5540 14288 5592 14340
rect 10600 14424 10652 14476
rect 11060 14467 11112 14476
rect 11060 14433 11069 14467
rect 11069 14433 11103 14467
rect 11103 14433 11112 14467
rect 11060 14424 11112 14433
rect 15200 14492 15252 14544
rect 18696 14492 18748 14544
rect 22928 14535 22980 14544
rect 22928 14501 22937 14535
rect 22937 14501 22971 14535
rect 22971 14501 22980 14535
rect 22928 14492 22980 14501
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 13820 14424 13872 14476
rect 16120 14424 16172 14476
rect 19800 14467 19852 14476
rect 19800 14433 19809 14467
rect 19809 14433 19843 14467
rect 19843 14433 19852 14467
rect 19800 14424 19852 14433
rect 13912 14356 13964 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 14832 14356 14884 14408
rect 15844 14356 15896 14408
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 19708 14356 19760 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 21456 14356 21508 14408
rect 24952 14467 25004 14476
rect 24952 14433 24961 14467
rect 24961 14433 24995 14467
rect 24995 14433 25004 14467
rect 24952 14424 25004 14433
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 12440 14288 12492 14340
rect 19340 14288 19392 14340
rect 26424 14356 26476 14408
rect 29736 14356 29788 14408
rect 30288 14356 30340 14408
rect 30932 14356 30984 14408
rect 31208 14399 31260 14408
rect 31208 14365 31217 14399
rect 31217 14365 31251 14399
rect 31251 14365 31260 14399
rect 31208 14356 31260 14365
rect 31024 14288 31076 14340
rect 32404 14424 32456 14476
rect 37740 14560 37792 14612
rect 39028 14560 39080 14612
rect 39396 14560 39448 14612
rect 40040 14535 40092 14544
rect 40040 14501 40049 14535
rect 40049 14501 40083 14535
rect 40083 14501 40092 14535
rect 40040 14492 40092 14501
rect 32680 14356 32732 14408
rect 36728 14399 36780 14408
rect 36728 14365 36737 14399
rect 36737 14365 36771 14399
rect 36771 14365 36780 14399
rect 36728 14356 36780 14365
rect 38752 14424 38804 14476
rect 39120 14424 39172 14476
rect 42432 14467 42484 14476
rect 42432 14433 42441 14467
rect 42441 14433 42475 14467
rect 42475 14433 42484 14467
rect 42432 14424 42484 14433
rect 42708 14424 42760 14476
rect 37280 14399 37332 14408
rect 37280 14365 37289 14399
rect 37289 14365 37323 14399
rect 37323 14365 37332 14399
rect 37280 14356 37332 14365
rect 37464 14356 37516 14408
rect 38476 14356 38528 14408
rect 40224 14399 40276 14408
rect 40224 14365 40233 14399
rect 40233 14365 40267 14399
rect 40267 14365 40276 14399
rect 40224 14356 40276 14365
rect 43904 14424 43956 14476
rect 51264 14560 51316 14612
rect 45284 14467 45336 14476
rect 45284 14433 45293 14467
rect 45293 14433 45327 14467
rect 45327 14433 45336 14467
rect 45284 14424 45336 14433
rect 55312 14560 55364 14612
rect 43536 14399 43588 14408
rect 43536 14365 43545 14399
rect 43545 14365 43579 14399
rect 43579 14365 43588 14399
rect 43536 14356 43588 14365
rect 33232 14288 33284 14340
rect 36636 14288 36688 14340
rect 37648 14288 37700 14340
rect 40776 14288 40828 14340
rect 42800 14288 42852 14340
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 10968 14220 11020 14272
rect 12532 14220 12584 14272
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 13452 14220 13504 14272
rect 14832 14220 14884 14272
rect 20076 14220 20128 14272
rect 20168 14263 20220 14272
rect 20168 14229 20177 14263
rect 20177 14229 20211 14263
rect 20211 14229 20220 14263
rect 20168 14220 20220 14229
rect 21180 14220 21232 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 22928 14220 22980 14272
rect 23664 14220 23716 14272
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 25596 14263 25648 14272
rect 25596 14229 25605 14263
rect 25605 14229 25639 14263
rect 25639 14229 25648 14263
rect 25596 14220 25648 14229
rect 25688 14220 25740 14272
rect 26148 14220 26200 14272
rect 28724 14263 28776 14272
rect 28724 14229 28733 14263
rect 28733 14229 28767 14263
rect 28767 14229 28776 14263
rect 28724 14220 28776 14229
rect 30288 14220 30340 14272
rect 30656 14263 30708 14272
rect 30656 14229 30665 14263
rect 30665 14229 30699 14263
rect 30699 14229 30708 14263
rect 30656 14220 30708 14229
rect 32496 14263 32548 14272
rect 32496 14229 32505 14263
rect 32505 14229 32539 14263
rect 32539 14229 32548 14263
rect 32496 14220 32548 14229
rect 33508 14220 33560 14272
rect 33784 14263 33836 14272
rect 33784 14229 33793 14263
rect 33793 14229 33827 14263
rect 33827 14229 33836 14263
rect 33784 14220 33836 14229
rect 35348 14263 35400 14272
rect 35348 14229 35357 14263
rect 35357 14229 35391 14263
rect 35391 14229 35400 14263
rect 35348 14220 35400 14229
rect 35900 14220 35952 14272
rect 37372 14220 37424 14272
rect 37924 14220 37976 14272
rect 38292 14220 38344 14272
rect 38660 14220 38712 14272
rect 40868 14263 40920 14272
rect 40868 14229 40877 14263
rect 40877 14229 40911 14263
rect 40911 14229 40920 14263
rect 40868 14220 40920 14229
rect 41144 14263 41196 14272
rect 41144 14229 41153 14263
rect 41153 14229 41187 14263
rect 41187 14229 41196 14263
rect 41144 14220 41196 14229
rect 42892 14220 42944 14272
rect 43812 14288 43864 14340
rect 49332 14467 49384 14476
rect 49332 14433 49341 14467
rect 49341 14433 49375 14467
rect 49375 14433 49384 14467
rect 49332 14424 49384 14433
rect 49516 14467 49568 14476
rect 49516 14433 49525 14467
rect 49525 14433 49559 14467
rect 49559 14433 49568 14467
rect 49516 14424 49568 14433
rect 48320 14288 48372 14340
rect 49700 14424 49752 14476
rect 51080 14467 51132 14476
rect 51080 14433 51089 14467
rect 51089 14433 51123 14467
rect 51123 14433 51132 14467
rect 51080 14424 51132 14433
rect 51264 14424 51316 14476
rect 54944 14492 54996 14544
rect 52368 14424 52420 14476
rect 55588 14424 55640 14476
rect 56048 14424 56100 14476
rect 56232 14467 56284 14476
rect 56232 14433 56241 14467
rect 56241 14433 56275 14467
rect 56275 14433 56284 14467
rect 56232 14424 56284 14433
rect 56508 14560 56560 14612
rect 56784 14424 56836 14476
rect 49884 14356 49936 14408
rect 50804 14399 50856 14408
rect 50804 14365 50813 14399
rect 50813 14365 50847 14399
rect 50847 14365 50856 14399
rect 50804 14356 50856 14365
rect 52000 14399 52052 14408
rect 52000 14365 52009 14399
rect 52009 14365 52043 14399
rect 52043 14365 52052 14399
rect 52000 14356 52052 14365
rect 53380 14399 53432 14408
rect 53380 14365 53414 14399
rect 53414 14365 53432 14399
rect 53380 14356 53432 14365
rect 56968 14399 57020 14408
rect 56968 14365 56977 14399
rect 56977 14365 57011 14399
rect 57011 14365 57020 14399
rect 56968 14356 57020 14365
rect 57796 14467 57848 14476
rect 57796 14433 57805 14467
rect 57805 14433 57839 14467
rect 57839 14433 57848 14467
rect 57796 14424 57848 14433
rect 57888 14356 57940 14408
rect 43444 14220 43496 14272
rect 45468 14220 45520 14272
rect 45744 14263 45796 14272
rect 45744 14229 45753 14263
rect 45753 14229 45787 14263
rect 45787 14229 45796 14263
rect 45744 14220 45796 14229
rect 47308 14263 47360 14272
rect 47308 14229 47317 14263
rect 47317 14229 47351 14263
rect 47351 14229 47360 14263
rect 47308 14220 47360 14229
rect 48780 14263 48832 14272
rect 48780 14229 48789 14263
rect 48789 14229 48823 14263
rect 48823 14229 48832 14263
rect 48780 14220 48832 14229
rect 48872 14263 48924 14272
rect 48872 14229 48881 14263
rect 48881 14229 48915 14263
rect 48915 14229 48924 14263
rect 48872 14220 48924 14229
rect 49976 14263 50028 14272
rect 49976 14229 49985 14263
rect 49985 14229 50019 14263
rect 50019 14229 50028 14263
rect 53012 14263 53064 14272
rect 49976 14220 50028 14229
rect 53012 14229 53021 14263
rect 53021 14229 53055 14263
rect 53055 14229 53064 14263
rect 53012 14220 53064 14229
rect 55036 14220 55088 14272
rect 57244 14263 57296 14272
rect 57244 14229 57253 14263
rect 57253 14229 57287 14263
rect 57287 14229 57296 14263
rect 57244 14220 57296 14229
rect 15394 14118 15446 14170
rect 15458 14118 15510 14170
rect 15522 14118 15574 14170
rect 15586 14118 15638 14170
rect 15650 14118 15702 14170
rect 29838 14118 29890 14170
rect 29902 14118 29954 14170
rect 29966 14118 30018 14170
rect 30030 14118 30082 14170
rect 30094 14118 30146 14170
rect 44282 14118 44334 14170
rect 44346 14118 44398 14170
rect 44410 14118 44462 14170
rect 44474 14118 44526 14170
rect 44538 14118 44590 14170
rect 58726 14118 58778 14170
rect 58790 14118 58842 14170
rect 58854 14118 58906 14170
rect 58918 14118 58970 14170
rect 58982 14118 59034 14170
rect 6920 14016 6972 14068
rect 7104 13948 7156 14000
rect 7104 13812 7156 13864
rect 7288 13812 7340 13864
rect 7840 13812 7892 13864
rect 8668 14016 8720 14068
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 8116 13948 8168 14000
rect 9496 13948 9548 14000
rect 11060 13948 11112 14000
rect 11980 13948 12032 14000
rect 12348 13880 12400 13932
rect 14832 14016 14884 14068
rect 15752 14016 15804 14068
rect 16948 14016 17000 14068
rect 13636 13948 13688 14000
rect 13820 13923 13872 13932
rect 13820 13889 13854 13923
rect 13854 13889 13872 13923
rect 13820 13880 13872 13889
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 15200 13880 15252 13932
rect 18328 14016 18380 14068
rect 19340 14016 19392 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 18788 13948 18840 14000
rect 19524 13880 19576 13932
rect 19708 13923 19760 13932
rect 19708 13889 19742 13923
rect 19742 13889 19760 13923
rect 19708 13880 19760 13889
rect 25412 14016 25464 14068
rect 25596 14016 25648 14068
rect 26148 14016 26200 14068
rect 10324 13812 10376 13864
rect 10416 13812 10468 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 21456 13855 21508 13864
rect 21456 13821 21465 13855
rect 21465 13821 21499 13855
rect 21499 13821 21508 13855
rect 21456 13812 21508 13821
rect 23572 13948 23624 14000
rect 23848 13948 23900 14000
rect 24308 13948 24360 14000
rect 19156 13744 19208 13796
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8852 13676 8904 13728
rect 12256 13676 12308 13728
rect 13268 13676 13320 13728
rect 17408 13676 17460 13728
rect 17868 13676 17920 13728
rect 17960 13676 18012 13728
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 21916 13744 21968 13796
rect 20444 13676 20496 13728
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 22468 13676 22520 13728
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 25872 13880 25924 13932
rect 29736 14016 29788 14068
rect 28724 13991 28776 14000
rect 28724 13957 28758 13991
rect 28758 13957 28776 13991
rect 28724 13948 28776 13957
rect 30656 14016 30708 14068
rect 30840 14016 30892 14068
rect 32496 14016 32548 14068
rect 32128 13948 32180 14000
rect 33416 14016 33468 14068
rect 33508 14016 33560 14068
rect 33600 14016 33652 14068
rect 35900 14016 35952 14068
rect 35992 14059 36044 14068
rect 35992 14025 36001 14059
rect 36001 14025 36035 14059
rect 36035 14025 36044 14059
rect 35992 14016 36044 14025
rect 36728 14016 36780 14068
rect 27252 13812 27304 13864
rect 26240 13744 26292 13796
rect 27620 13744 27672 13796
rect 31024 13923 31076 13932
rect 31024 13889 31033 13923
rect 31033 13889 31067 13923
rect 31067 13889 31076 13923
rect 31024 13880 31076 13889
rect 30840 13812 30892 13864
rect 31116 13855 31168 13864
rect 31116 13821 31150 13855
rect 31150 13821 31168 13855
rect 31116 13812 31168 13821
rect 32036 13812 32088 13864
rect 30472 13744 30524 13796
rect 38200 14016 38252 14068
rect 38936 14016 38988 14068
rect 40224 14016 40276 14068
rect 40868 14016 40920 14068
rect 43536 14016 43588 14068
rect 43628 14016 43680 14068
rect 45008 14016 45060 14068
rect 45468 14016 45520 14068
rect 45744 14016 45796 14068
rect 47032 14016 47084 14068
rect 48320 14059 48372 14068
rect 48320 14025 48329 14059
rect 48329 14025 48363 14059
rect 48363 14025 48372 14059
rect 48320 14016 48372 14025
rect 49516 14016 49568 14068
rect 40040 13948 40092 14000
rect 41144 13991 41196 14000
rect 34612 13923 34664 13932
rect 34612 13889 34621 13923
rect 34621 13889 34655 13923
rect 34655 13889 34664 13923
rect 34612 13880 34664 13889
rect 37188 13880 37240 13932
rect 37372 13880 37424 13932
rect 37648 13880 37700 13932
rect 38200 13923 38252 13932
rect 38200 13889 38209 13923
rect 38209 13889 38243 13923
rect 38243 13889 38252 13923
rect 38200 13880 38252 13889
rect 36544 13812 36596 13864
rect 36728 13812 36780 13864
rect 38660 13812 38712 13864
rect 39396 13855 39448 13864
rect 39396 13821 39405 13855
rect 39405 13821 39439 13855
rect 39439 13821 39448 13855
rect 39396 13812 39448 13821
rect 39764 13812 39816 13864
rect 40500 13855 40552 13864
rect 40500 13821 40509 13855
rect 40509 13821 40543 13855
rect 40543 13821 40552 13855
rect 40500 13812 40552 13821
rect 41144 13957 41167 13991
rect 41167 13957 41196 13991
rect 41144 13948 41196 13957
rect 43812 13923 43864 13932
rect 43812 13889 43821 13923
rect 43821 13889 43855 13923
rect 43855 13889 43864 13923
rect 43812 13880 43864 13889
rect 43904 13923 43956 13932
rect 43904 13889 43938 13923
rect 43938 13889 43956 13923
rect 43904 13880 43956 13889
rect 44088 13923 44140 13932
rect 44088 13889 44097 13923
rect 44097 13889 44131 13923
rect 44131 13889 44140 13923
rect 44088 13880 44140 13889
rect 45376 13880 45428 13932
rect 45836 13880 45888 13932
rect 47308 13948 47360 14000
rect 48872 13923 48924 13932
rect 48872 13889 48881 13923
rect 48881 13889 48915 13923
rect 48915 13889 48924 13923
rect 48872 13880 48924 13889
rect 49976 13948 50028 14000
rect 50436 13948 50488 14000
rect 50896 14016 50948 14068
rect 52000 14016 52052 14068
rect 55220 14016 55272 14068
rect 58440 14016 58492 14068
rect 57704 13948 57756 14000
rect 57888 13991 57940 14000
rect 57888 13957 57897 13991
rect 57897 13957 57931 13991
rect 57931 13957 57940 13991
rect 57888 13948 57940 13957
rect 51908 13880 51960 13932
rect 54300 13880 54352 13932
rect 54944 13923 54996 13932
rect 54944 13889 54953 13923
rect 54953 13889 54987 13923
rect 54987 13889 54996 13923
rect 54944 13880 54996 13889
rect 23848 13676 23900 13728
rect 27712 13676 27764 13728
rect 28080 13719 28132 13728
rect 28080 13685 28089 13719
rect 28089 13685 28123 13719
rect 28123 13685 28132 13719
rect 28080 13676 28132 13685
rect 29920 13676 29972 13728
rect 33600 13719 33652 13728
rect 33600 13685 33609 13719
rect 33609 13685 33643 13719
rect 33643 13685 33652 13719
rect 33600 13676 33652 13685
rect 37832 13744 37884 13796
rect 42708 13855 42760 13864
rect 42708 13821 42717 13855
rect 42717 13821 42751 13855
rect 42751 13821 42760 13855
rect 42708 13812 42760 13821
rect 42984 13812 43036 13864
rect 45008 13812 45060 13864
rect 51080 13812 51132 13864
rect 52000 13812 52052 13864
rect 52276 13812 52328 13864
rect 53012 13812 53064 13864
rect 39948 13676 40000 13728
rect 40040 13719 40092 13728
rect 40040 13685 40049 13719
rect 40049 13685 40083 13719
rect 40083 13685 40092 13719
rect 40040 13676 40092 13685
rect 43628 13744 43680 13796
rect 41604 13676 41656 13728
rect 44088 13676 44140 13728
rect 46572 13676 46624 13728
rect 46756 13719 46808 13728
rect 46756 13685 46765 13719
rect 46765 13685 46799 13719
rect 46799 13685 46808 13719
rect 46756 13676 46808 13685
rect 50436 13676 50488 13728
rect 51264 13676 51316 13728
rect 55496 13855 55548 13864
rect 55496 13821 55505 13855
rect 55505 13821 55539 13855
rect 55539 13821 55548 13855
rect 55496 13812 55548 13821
rect 56140 13855 56192 13864
rect 56140 13821 56149 13855
rect 56149 13821 56183 13855
rect 56183 13821 56192 13855
rect 56140 13812 56192 13821
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 22616 13574 22668 13626
rect 22680 13574 22732 13626
rect 22744 13574 22796 13626
rect 22808 13574 22860 13626
rect 22872 13574 22924 13626
rect 37060 13574 37112 13626
rect 37124 13574 37176 13626
rect 37188 13574 37240 13626
rect 37252 13574 37304 13626
rect 37316 13574 37368 13626
rect 51504 13574 51556 13626
rect 51568 13574 51620 13626
rect 51632 13574 51684 13626
rect 51696 13574 51748 13626
rect 51760 13574 51812 13626
rect 10876 13472 10928 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13268 13472 13320 13524
rect 8852 13336 8904 13388
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 3884 13268 3936 13320
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6828 13268 6880 13320
rect 12348 13268 12400 13320
rect 14924 13336 14976 13388
rect 16028 13336 16080 13388
rect 17040 13404 17092 13456
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 18512 13472 18564 13524
rect 20168 13472 20220 13524
rect 21456 13472 21508 13524
rect 22468 13404 22520 13456
rect 23940 13472 23992 13524
rect 26424 13515 26476 13524
rect 26424 13481 26433 13515
rect 26433 13481 26467 13515
rect 26467 13481 26476 13515
rect 26424 13472 26476 13481
rect 29920 13472 29972 13524
rect 30380 13472 30432 13524
rect 31484 13472 31536 13524
rect 31208 13404 31260 13456
rect 32404 13404 32456 13456
rect 34520 13404 34572 13456
rect 20444 13379 20496 13388
rect 20444 13345 20453 13379
rect 20453 13345 20487 13379
rect 20487 13345 20496 13379
rect 20444 13336 20496 13345
rect 20720 13336 20772 13388
rect 15844 13268 15896 13320
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 17408 13268 17460 13320
rect 19064 13268 19116 13320
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 20076 13311 20128 13320
rect 20076 13277 20094 13311
rect 20094 13277 20128 13311
rect 20076 13268 20128 13277
rect 20168 13311 20220 13320
rect 20168 13277 20177 13311
rect 20177 13277 20211 13311
rect 20211 13277 20220 13311
rect 20168 13268 20220 13277
rect 6460 13200 6512 13252
rect 8760 13200 8812 13252
rect 13912 13200 13964 13252
rect 15108 13200 15160 13252
rect 17040 13200 17092 13252
rect 18420 13200 18472 13252
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 21364 13268 21416 13320
rect 2964 13175 3016 13184
rect 2964 13141 2973 13175
rect 2973 13141 3007 13175
rect 3007 13141 3016 13175
rect 2964 13132 3016 13141
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 10876 13132 10928 13184
rect 13636 13132 13688 13184
rect 14372 13132 14424 13184
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 15844 13132 15896 13184
rect 16028 13132 16080 13184
rect 16764 13132 16816 13184
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 17868 13132 17920 13184
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 21456 13200 21508 13252
rect 22376 13336 22428 13388
rect 24768 13336 24820 13388
rect 25596 13336 25648 13388
rect 25780 13336 25832 13388
rect 26148 13379 26200 13388
rect 26148 13345 26157 13379
rect 26157 13345 26191 13379
rect 26191 13345 26200 13379
rect 26148 13336 26200 13345
rect 25320 13311 25372 13320
rect 25320 13277 25338 13311
rect 25338 13277 25372 13311
rect 25320 13268 25372 13277
rect 26240 13268 26292 13320
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 28080 13268 28132 13320
rect 29736 13268 29788 13320
rect 34612 13336 34664 13388
rect 45836 13515 45888 13524
rect 45836 13481 45845 13515
rect 45845 13481 45879 13515
rect 45879 13481 45888 13515
rect 45836 13472 45888 13481
rect 43352 13404 43404 13456
rect 41604 13336 41656 13388
rect 45192 13379 45244 13388
rect 45192 13345 45201 13379
rect 45201 13345 45235 13379
rect 45235 13345 45244 13379
rect 45192 13336 45244 13345
rect 49700 13515 49752 13524
rect 49700 13481 49709 13515
rect 49709 13481 49743 13515
rect 49743 13481 49752 13515
rect 49700 13472 49752 13481
rect 55496 13472 55548 13524
rect 55588 13515 55640 13524
rect 55588 13481 55597 13515
rect 55597 13481 55631 13515
rect 55631 13481 55640 13515
rect 55588 13472 55640 13481
rect 56140 13472 56192 13524
rect 46204 13404 46256 13456
rect 27712 13200 27764 13252
rect 28632 13200 28684 13252
rect 30472 13200 30524 13252
rect 30932 13200 30984 13252
rect 19892 13132 19944 13184
rect 21548 13175 21600 13184
rect 21548 13141 21557 13175
rect 21557 13141 21591 13175
rect 21591 13141 21600 13175
rect 21548 13132 21600 13141
rect 21916 13132 21968 13184
rect 25688 13132 25740 13184
rect 31024 13132 31076 13184
rect 32128 13175 32180 13184
rect 32128 13141 32137 13175
rect 32137 13141 32171 13175
rect 32171 13141 32180 13175
rect 32128 13132 32180 13141
rect 32680 13200 32732 13252
rect 32864 13243 32916 13252
rect 32864 13209 32898 13243
rect 32898 13209 32916 13243
rect 32864 13200 32916 13209
rect 35808 13268 35860 13320
rect 39764 13268 39816 13320
rect 39856 13311 39908 13320
rect 39856 13277 39865 13311
rect 39865 13277 39899 13311
rect 39899 13277 39908 13311
rect 39856 13268 39908 13277
rect 44640 13268 44692 13320
rect 45376 13268 45428 13320
rect 35164 13200 35216 13252
rect 35440 13200 35492 13252
rect 32956 13132 33008 13184
rect 34336 13175 34388 13184
rect 34336 13141 34345 13175
rect 34345 13141 34379 13175
rect 34379 13141 34388 13175
rect 39396 13200 39448 13252
rect 42340 13200 42392 13252
rect 44732 13200 44784 13252
rect 45008 13200 45060 13252
rect 46112 13336 46164 13388
rect 46572 13336 46624 13388
rect 48136 13336 48188 13388
rect 46756 13268 46808 13320
rect 47216 13311 47268 13320
rect 47216 13277 47225 13311
rect 47225 13277 47259 13311
rect 47259 13277 47268 13311
rect 47216 13268 47268 13277
rect 48780 13336 48832 13388
rect 56692 13336 56744 13388
rect 56784 13379 56836 13388
rect 56784 13345 56793 13379
rect 56793 13345 56827 13379
rect 56827 13345 56836 13379
rect 56784 13336 56836 13345
rect 58440 13379 58492 13388
rect 58440 13345 58449 13379
rect 58449 13345 58483 13379
rect 58483 13345 58492 13379
rect 58440 13336 58492 13345
rect 50804 13268 50856 13320
rect 56968 13268 57020 13320
rect 34336 13132 34388 13141
rect 36084 13175 36136 13184
rect 36084 13141 36093 13175
rect 36093 13141 36127 13175
rect 36127 13141 36136 13175
rect 36084 13132 36136 13141
rect 37740 13175 37792 13184
rect 37740 13141 37749 13175
rect 37749 13141 37783 13175
rect 37783 13141 37792 13175
rect 37740 13132 37792 13141
rect 37924 13132 37976 13184
rect 39304 13175 39356 13184
rect 39304 13141 39313 13175
rect 39313 13141 39347 13175
rect 39347 13141 39356 13175
rect 39304 13132 39356 13141
rect 42524 13132 42576 13184
rect 43168 13175 43220 13184
rect 43168 13141 43177 13175
rect 43177 13141 43211 13175
rect 43211 13141 43220 13175
rect 43168 13132 43220 13141
rect 45284 13175 45336 13184
rect 45284 13141 45293 13175
rect 45293 13141 45327 13175
rect 45327 13141 45336 13175
rect 45284 13132 45336 13141
rect 46296 13175 46348 13184
rect 46296 13141 46305 13175
rect 46305 13141 46339 13175
rect 46339 13141 46348 13175
rect 46296 13132 46348 13141
rect 47400 13175 47452 13184
rect 47400 13141 47409 13175
rect 47409 13141 47443 13175
rect 47443 13141 47452 13175
rect 47400 13132 47452 13141
rect 50436 13175 50488 13184
rect 50436 13141 50445 13175
rect 50445 13141 50479 13175
rect 50479 13141 50488 13175
rect 50436 13132 50488 13141
rect 56876 13132 56928 13184
rect 57520 13132 57572 13184
rect 15394 13030 15446 13082
rect 15458 13030 15510 13082
rect 15522 13030 15574 13082
rect 15586 13030 15638 13082
rect 15650 13030 15702 13082
rect 29838 13030 29890 13082
rect 29902 13030 29954 13082
rect 29966 13030 30018 13082
rect 30030 13030 30082 13082
rect 30094 13030 30146 13082
rect 44282 13030 44334 13082
rect 44346 13030 44398 13082
rect 44410 13030 44462 13082
rect 44474 13030 44526 13082
rect 44538 13030 44590 13082
rect 58726 13030 58778 13082
rect 58790 13030 58842 13082
rect 58854 13030 58906 13082
rect 58918 13030 58970 13082
rect 58982 13030 59034 13082
rect 7748 12928 7800 12980
rect 8116 12928 8168 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12716 12928 12768 12980
rect 13636 12928 13688 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 13820 12928 13872 12980
rect 2964 12903 3016 12912
rect 2964 12869 2998 12903
rect 2998 12869 3016 12903
rect 2964 12860 3016 12869
rect 7012 12903 7064 12912
rect 7012 12869 7021 12903
rect 7021 12869 7055 12903
rect 7055 12869 7064 12903
rect 7012 12860 7064 12869
rect 7656 12860 7708 12912
rect 20996 12928 21048 12980
rect 21456 12971 21508 12980
rect 21456 12937 21465 12971
rect 21465 12937 21499 12971
rect 21499 12937 21508 12971
rect 21456 12928 21508 12937
rect 22100 12928 22152 12980
rect 25320 12971 25372 12980
rect 25320 12937 25329 12971
rect 25329 12937 25363 12971
rect 25363 12937 25372 12971
rect 25320 12928 25372 12937
rect 26240 12928 26292 12980
rect 29000 12928 29052 12980
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 30932 12928 30984 12980
rect 31024 12928 31076 12980
rect 32036 12928 32088 12980
rect 32864 12971 32916 12980
rect 32864 12937 32873 12971
rect 32873 12937 32907 12971
rect 32907 12937 32916 12971
rect 32864 12928 32916 12937
rect 33784 12928 33836 12980
rect 33968 12971 34020 12980
rect 33968 12937 33977 12971
rect 33977 12937 34011 12971
rect 34011 12937 34020 12971
rect 33968 12928 34020 12937
rect 34244 12928 34296 12980
rect 35164 12971 35216 12980
rect 35164 12937 35173 12971
rect 35173 12937 35207 12971
rect 35207 12937 35216 12971
rect 35164 12928 35216 12937
rect 35808 12928 35860 12980
rect 10232 12792 10284 12844
rect 14372 12860 14424 12912
rect 15016 12860 15068 12912
rect 15200 12860 15252 12912
rect 15752 12860 15804 12912
rect 19984 12903 20036 12912
rect 19984 12869 19993 12903
rect 19993 12869 20027 12903
rect 20027 12869 20036 12903
rect 19984 12860 20036 12869
rect 30380 12860 30432 12912
rect 7380 12724 7432 12776
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 17592 12792 17644 12844
rect 19064 12792 19116 12844
rect 20904 12792 20956 12844
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 23020 12792 23072 12844
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 26424 12792 26476 12844
rect 14832 12724 14884 12776
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 6828 12656 6880 12708
rect 13912 12656 13964 12708
rect 14556 12656 14608 12708
rect 23848 12724 23900 12776
rect 25412 12767 25464 12776
rect 25412 12733 25421 12767
rect 25421 12733 25455 12767
rect 25455 12733 25464 12767
rect 25412 12724 25464 12733
rect 27988 12792 28040 12844
rect 34980 12860 35032 12912
rect 29184 12724 29236 12776
rect 26884 12656 26936 12708
rect 28908 12656 28960 12708
rect 35348 12792 35400 12844
rect 36084 12860 36136 12912
rect 36636 12903 36688 12912
rect 36636 12869 36645 12903
rect 36645 12869 36679 12903
rect 36679 12869 36688 12903
rect 36636 12860 36688 12869
rect 37556 12903 37608 12912
rect 37556 12869 37565 12903
rect 37565 12869 37599 12903
rect 37599 12869 37608 12903
rect 37556 12860 37608 12869
rect 37740 12860 37792 12912
rect 39856 12928 39908 12980
rect 41604 12928 41656 12980
rect 42984 12928 43036 12980
rect 43444 12928 43496 12980
rect 45284 12928 45336 12980
rect 45376 12971 45428 12980
rect 45376 12937 45385 12971
rect 45385 12937 45419 12971
rect 45419 12937 45428 12971
rect 45376 12928 45428 12937
rect 47216 12928 47268 12980
rect 47400 12928 47452 12980
rect 49976 12928 50028 12980
rect 40040 12860 40092 12912
rect 40776 12903 40828 12912
rect 40776 12869 40785 12903
rect 40785 12869 40819 12903
rect 40819 12869 40828 12903
rect 40776 12860 40828 12869
rect 42524 12860 42576 12912
rect 43720 12860 43772 12912
rect 45192 12792 45244 12844
rect 54944 12928 54996 12980
rect 55128 12928 55180 12980
rect 55588 12928 55640 12980
rect 58072 12860 58124 12912
rect 50528 12835 50580 12844
rect 50528 12801 50562 12835
rect 50562 12801 50580 12835
rect 50528 12792 50580 12801
rect 56968 12835 57020 12844
rect 56968 12801 56977 12835
rect 56977 12801 57011 12835
rect 57011 12801 57020 12835
rect 56968 12792 57020 12801
rect 58440 12835 58492 12844
rect 58440 12801 58449 12835
rect 58449 12801 58483 12835
rect 58483 12801 58492 12835
rect 58440 12792 58492 12801
rect 29644 12767 29696 12776
rect 29644 12733 29653 12767
rect 29653 12733 29687 12767
rect 29687 12733 29696 12767
rect 29644 12724 29696 12733
rect 31300 12724 31352 12776
rect 33968 12724 34020 12776
rect 31116 12656 31168 12708
rect 40960 12767 41012 12776
rect 40960 12733 40969 12767
rect 40969 12733 41003 12767
rect 41003 12733 41012 12767
rect 40960 12724 41012 12733
rect 43076 12767 43128 12776
rect 43076 12733 43085 12767
rect 43085 12733 43119 12767
rect 43119 12733 43128 12767
rect 43076 12724 43128 12733
rect 48320 12767 48372 12776
rect 48320 12733 48329 12767
rect 48329 12733 48363 12767
rect 48363 12733 48372 12767
rect 48320 12724 48372 12733
rect 54668 12767 54720 12776
rect 54668 12733 54677 12767
rect 54677 12733 54711 12767
rect 54711 12733 54720 12767
rect 54668 12724 54720 12733
rect 2964 12588 3016 12640
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 7012 12588 7064 12640
rect 8024 12588 8076 12640
rect 10324 12588 10376 12640
rect 14740 12631 14792 12640
rect 14740 12597 14749 12631
rect 14749 12597 14783 12631
rect 14783 12597 14792 12631
rect 14740 12588 14792 12597
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 21088 12588 21140 12640
rect 21272 12588 21324 12640
rect 23848 12631 23900 12640
rect 23848 12597 23857 12631
rect 23857 12597 23891 12631
rect 23891 12597 23900 12631
rect 23848 12588 23900 12597
rect 28448 12588 28500 12640
rect 29000 12631 29052 12640
rect 29000 12597 29009 12631
rect 29009 12597 29043 12631
rect 29043 12597 29052 12631
rect 29000 12588 29052 12597
rect 29736 12588 29788 12640
rect 30656 12588 30708 12640
rect 32680 12631 32732 12640
rect 32680 12597 32689 12631
rect 32689 12597 32723 12631
rect 32723 12597 32732 12631
rect 32680 12588 32732 12597
rect 38476 12588 38528 12640
rect 40316 12631 40368 12640
rect 40316 12597 40325 12631
rect 40325 12597 40359 12631
rect 40359 12597 40368 12631
rect 40316 12588 40368 12597
rect 40408 12631 40460 12640
rect 40408 12597 40417 12631
rect 40417 12597 40451 12631
rect 40451 12597 40460 12631
rect 40408 12588 40460 12597
rect 42432 12588 42484 12640
rect 42616 12588 42668 12640
rect 44088 12588 44140 12640
rect 50068 12656 50120 12708
rect 57060 12767 57112 12776
rect 57060 12733 57069 12767
rect 57069 12733 57103 12767
rect 57103 12733 57112 12767
rect 57060 12724 57112 12733
rect 57152 12767 57204 12776
rect 57152 12733 57161 12767
rect 57161 12733 57195 12767
rect 57195 12733 57204 12767
rect 57152 12724 57204 12733
rect 47768 12631 47820 12640
rect 47768 12597 47777 12631
rect 47777 12597 47811 12631
rect 47811 12597 47820 12631
rect 47768 12588 47820 12597
rect 52276 12588 52328 12640
rect 54116 12631 54168 12640
rect 54116 12597 54125 12631
rect 54125 12597 54159 12631
rect 54159 12597 54168 12631
rect 54116 12588 54168 12597
rect 56692 12588 56744 12640
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 22616 12486 22668 12538
rect 22680 12486 22732 12538
rect 22744 12486 22796 12538
rect 22808 12486 22860 12538
rect 22872 12486 22924 12538
rect 37060 12486 37112 12538
rect 37124 12486 37176 12538
rect 37188 12486 37240 12538
rect 37252 12486 37304 12538
rect 37316 12486 37368 12538
rect 51504 12486 51556 12538
rect 51568 12486 51620 12538
rect 51632 12486 51684 12538
rect 51696 12486 51748 12538
rect 51760 12486 51812 12538
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 7564 12384 7616 12436
rect 10784 12384 10836 12436
rect 13912 12384 13964 12436
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 7748 12316 7800 12368
rect 13544 12316 13596 12368
rect 15936 12384 15988 12436
rect 16764 12384 16816 12436
rect 17592 12427 17644 12436
rect 17592 12393 17601 12427
rect 17601 12393 17635 12427
rect 17635 12393 17644 12427
rect 17592 12384 17644 12393
rect 18880 12384 18932 12436
rect 19984 12384 20036 12436
rect 21088 12384 21140 12436
rect 21548 12427 21600 12436
rect 21548 12393 21557 12427
rect 21557 12393 21591 12427
rect 21591 12393 21600 12427
rect 21548 12384 21600 12393
rect 23020 12384 23072 12436
rect 23388 12384 23440 12436
rect 2964 12248 3016 12257
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 2964 12112 3016 12164
rect 3884 12180 3936 12232
rect 6644 12180 6696 12232
rect 9496 12248 9548 12300
rect 10508 12248 10560 12300
rect 12164 12248 12216 12300
rect 14096 12248 14148 12300
rect 8024 12180 8076 12232
rect 10232 12180 10284 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 12256 12180 12308 12232
rect 13912 12180 13964 12232
rect 14280 12180 14332 12232
rect 14740 12180 14792 12232
rect 17316 12180 17368 12232
rect 20168 12248 20220 12300
rect 20812 12248 20864 12300
rect 4252 12112 4304 12164
rect 11428 12112 11480 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 3056 12087 3108 12096
rect 3056 12053 3065 12087
rect 3065 12053 3099 12087
rect 3099 12053 3108 12087
rect 3056 12044 3108 12053
rect 3332 12044 3384 12096
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 5080 12044 5132 12096
rect 7564 12087 7616 12096
rect 7564 12053 7573 12087
rect 7573 12053 7607 12087
rect 7607 12053 7616 12087
rect 7564 12044 7616 12053
rect 8668 12044 8720 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 10968 12044 11020 12096
rect 12716 12044 12768 12096
rect 15752 12155 15804 12164
rect 15752 12121 15761 12155
rect 15761 12121 15795 12155
rect 15795 12121 15804 12155
rect 15752 12112 15804 12121
rect 20076 12180 20128 12232
rect 18788 12155 18840 12164
rect 18788 12121 18797 12155
rect 18797 12121 18831 12155
rect 18831 12121 18840 12155
rect 18788 12112 18840 12121
rect 13912 12044 13964 12096
rect 16120 12044 16172 12096
rect 16396 12044 16448 12096
rect 18328 12044 18380 12096
rect 19892 12087 19944 12096
rect 19892 12053 19901 12087
rect 19901 12053 19935 12087
rect 19935 12053 19944 12087
rect 19892 12044 19944 12053
rect 20904 12155 20956 12164
rect 20904 12121 20913 12155
rect 20913 12121 20947 12155
rect 20947 12121 20956 12155
rect 20904 12112 20956 12121
rect 20720 12044 20772 12096
rect 20996 12044 21048 12096
rect 21456 12316 21508 12368
rect 22100 12291 22152 12300
rect 22100 12257 22109 12291
rect 22109 12257 22143 12291
rect 22143 12257 22152 12291
rect 22100 12248 22152 12257
rect 23848 12291 23900 12300
rect 23848 12257 23857 12291
rect 23857 12257 23891 12291
rect 23891 12257 23900 12291
rect 23848 12248 23900 12257
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 25136 12180 25188 12232
rect 26424 12384 26476 12436
rect 28632 12427 28684 12436
rect 28632 12393 28641 12427
rect 28641 12393 28675 12427
rect 28675 12393 28684 12427
rect 28632 12384 28684 12393
rect 29184 12384 29236 12436
rect 29460 12384 29512 12436
rect 29736 12427 29788 12436
rect 29736 12393 29745 12427
rect 29745 12393 29779 12427
rect 29779 12393 29788 12427
rect 29736 12384 29788 12393
rect 30288 12384 30340 12436
rect 40776 12384 40828 12436
rect 42340 12427 42392 12436
rect 42340 12393 42349 12427
rect 42349 12393 42383 12427
rect 42383 12393 42392 12427
rect 42340 12384 42392 12393
rect 42984 12384 43036 12436
rect 44732 12427 44784 12436
rect 44732 12393 44741 12427
rect 44741 12393 44775 12427
rect 44775 12393 44784 12427
rect 44732 12384 44784 12393
rect 45192 12384 45244 12436
rect 45560 12427 45612 12436
rect 45560 12393 45569 12427
rect 45569 12393 45603 12427
rect 45603 12393 45612 12427
rect 45560 12384 45612 12393
rect 46112 12384 46164 12436
rect 45100 12316 45152 12368
rect 46480 12316 46532 12368
rect 50528 12384 50580 12436
rect 52000 12427 52052 12436
rect 52000 12393 52009 12427
rect 52009 12393 52043 12427
rect 52043 12393 52052 12427
rect 52000 12384 52052 12393
rect 53840 12384 53892 12436
rect 26240 12248 26292 12300
rect 29184 12291 29236 12300
rect 29184 12257 29193 12291
rect 29193 12257 29227 12291
rect 29227 12257 29236 12291
rect 29184 12248 29236 12257
rect 30656 12291 30708 12300
rect 30656 12257 30665 12291
rect 30665 12257 30699 12291
rect 30699 12257 30708 12291
rect 30656 12248 30708 12257
rect 39304 12248 39356 12300
rect 40408 12248 40460 12300
rect 42892 12291 42944 12300
rect 42892 12257 42901 12291
rect 42901 12257 42935 12291
rect 42935 12257 42944 12291
rect 42892 12248 42944 12257
rect 43168 12248 43220 12300
rect 44088 12291 44140 12300
rect 44088 12257 44097 12291
rect 44097 12257 44131 12291
rect 44131 12257 44140 12291
rect 44088 12248 44140 12257
rect 47308 12291 47360 12300
rect 25872 12112 25924 12164
rect 23020 12044 23072 12096
rect 23388 12044 23440 12096
rect 24492 12044 24544 12096
rect 24860 12044 24912 12096
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 25228 12044 25280 12096
rect 27620 12180 27672 12232
rect 28264 12180 28316 12232
rect 37648 12180 37700 12232
rect 39396 12180 39448 12232
rect 44640 12180 44692 12232
rect 46756 12180 46808 12232
rect 47308 12257 47317 12291
rect 47317 12257 47351 12291
rect 47351 12257 47360 12291
rect 47308 12248 47360 12257
rect 54668 12384 54720 12436
rect 55312 12384 55364 12436
rect 56600 12384 56652 12436
rect 47216 12223 47268 12232
rect 47216 12189 47225 12223
rect 47225 12189 47259 12223
rect 47259 12189 47268 12223
rect 47216 12180 47268 12189
rect 51080 12223 51132 12232
rect 51080 12189 51089 12223
rect 51089 12189 51123 12223
rect 51123 12189 51132 12223
rect 51080 12180 51132 12189
rect 52368 12180 52420 12232
rect 55312 12223 55364 12232
rect 55312 12189 55321 12223
rect 55321 12189 55355 12223
rect 55355 12189 55364 12223
rect 55312 12180 55364 12189
rect 56232 12180 56284 12232
rect 56692 12223 56744 12232
rect 56692 12189 56726 12223
rect 56726 12189 56744 12223
rect 56692 12180 56744 12189
rect 42616 12112 42668 12164
rect 27620 12087 27672 12096
rect 27620 12053 27629 12087
rect 27629 12053 27663 12087
rect 27663 12053 27672 12087
rect 27620 12044 27672 12053
rect 27804 12044 27856 12096
rect 31116 12087 31168 12096
rect 31116 12053 31125 12087
rect 31125 12053 31159 12087
rect 31159 12053 31168 12087
rect 31116 12044 31168 12053
rect 36084 12044 36136 12096
rect 36912 12044 36964 12096
rect 38292 12044 38344 12096
rect 41788 12044 41840 12096
rect 43076 12044 43128 12096
rect 45560 12112 45612 12164
rect 46480 12044 46532 12096
rect 49056 12112 49108 12164
rect 52092 12155 52144 12164
rect 52092 12121 52101 12155
rect 52101 12121 52135 12155
rect 52135 12121 52144 12155
rect 52092 12112 52144 12121
rect 56140 12112 56192 12164
rect 48596 12044 48648 12096
rect 48780 12087 48832 12096
rect 48780 12053 48789 12087
rect 48789 12053 48823 12087
rect 48823 12053 48832 12087
rect 48780 12044 48832 12053
rect 51356 12044 51408 12096
rect 52920 12044 52972 12096
rect 54668 12044 54720 12096
rect 57060 12044 57112 12096
rect 15394 11942 15446 11994
rect 15458 11942 15510 11994
rect 15522 11942 15574 11994
rect 15586 11942 15638 11994
rect 15650 11942 15702 11994
rect 29838 11942 29890 11994
rect 29902 11942 29954 11994
rect 29966 11942 30018 11994
rect 30030 11942 30082 11994
rect 30094 11942 30146 11994
rect 44282 11942 44334 11994
rect 44346 11942 44398 11994
rect 44410 11942 44462 11994
rect 44474 11942 44526 11994
rect 44538 11942 44590 11994
rect 58726 11942 58778 11994
rect 58790 11942 58842 11994
rect 58854 11942 58906 11994
rect 58918 11942 58970 11994
rect 58982 11942 59034 11994
rect 1584 11840 1636 11892
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3056 11840 3108 11892
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 7288 11772 7340 11824
rect 11244 11840 11296 11892
rect 16488 11840 16540 11892
rect 19708 11840 19760 11892
rect 23756 11883 23808 11892
rect 23756 11849 23765 11883
rect 23765 11849 23799 11883
rect 23799 11849 23808 11883
rect 23756 11840 23808 11849
rect 24952 11840 25004 11892
rect 29736 11840 29788 11892
rect 34888 11840 34940 11892
rect 38568 11840 38620 11892
rect 41604 11840 41656 11892
rect 44456 11840 44508 11892
rect 46756 11883 46808 11892
rect 46756 11849 46765 11883
rect 46765 11849 46799 11883
rect 46799 11849 46808 11883
rect 46756 11840 46808 11849
rect 48320 11840 48372 11892
rect 49056 11883 49108 11892
rect 49056 11849 49065 11883
rect 49065 11849 49099 11883
rect 49099 11849 49108 11883
rect 49056 11840 49108 11849
rect 55312 11840 55364 11892
rect 4712 11704 4764 11756
rect 7472 11747 7524 11756
rect 7472 11713 7490 11747
rect 7490 11713 7524 11747
rect 7472 11704 7524 11713
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 4804 11679 4856 11688
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 8024 11636 8076 11688
rect 3148 11568 3200 11620
rect 4068 11568 4120 11620
rect 23664 11772 23716 11824
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11612 11704 11664 11756
rect 12072 11704 12124 11756
rect 12348 11704 12400 11756
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10324 11636 10376 11688
rect 10968 11636 11020 11688
rect 13728 11704 13780 11756
rect 16304 11704 16356 11756
rect 3424 11500 3476 11552
rect 6000 11500 6052 11552
rect 6644 11500 6696 11552
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 10876 11500 10928 11552
rect 10968 11543 11020 11552
rect 10968 11509 10977 11543
rect 10977 11509 11011 11543
rect 11011 11509 11020 11543
rect 10968 11500 11020 11509
rect 11060 11500 11112 11552
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 18144 11704 18196 11756
rect 19800 11704 19852 11756
rect 19892 11704 19944 11756
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 20076 11636 20128 11688
rect 20168 11636 20220 11688
rect 29644 11772 29696 11824
rect 31668 11772 31720 11824
rect 35440 11815 35492 11824
rect 35440 11781 35449 11815
rect 35449 11781 35483 11815
rect 35483 11781 35492 11815
rect 35440 11772 35492 11781
rect 54116 11772 54168 11824
rect 29184 11747 29236 11756
rect 29184 11713 29193 11747
rect 29193 11713 29227 11747
rect 29227 11713 29236 11747
rect 29184 11704 29236 11713
rect 35072 11747 35124 11756
rect 35072 11713 35081 11747
rect 35081 11713 35115 11747
rect 35115 11713 35124 11747
rect 35072 11704 35124 11713
rect 38108 11747 38160 11756
rect 38108 11713 38117 11747
rect 38117 11713 38151 11747
rect 38151 11713 38160 11747
rect 38108 11704 38160 11713
rect 46940 11747 46992 11756
rect 46940 11713 46949 11747
rect 46949 11713 46983 11747
rect 46983 11713 46992 11747
rect 46940 11704 46992 11713
rect 48872 11704 48924 11756
rect 49976 11704 50028 11756
rect 50436 11747 50488 11756
rect 50436 11713 50445 11747
rect 50445 11713 50479 11747
rect 50479 11713 50488 11747
rect 50436 11704 50488 11713
rect 51172 11747 51224 11756
rect 51172 11713 51181 11747
rect 51181 11713 51215 11747
rect 51215 11713 51224 11747
rect 51172 11704 51224 11713
rect 56232 11840 56284 11892
rect 57060 11840 57112 11892
rect 56140 11704 56192 11756
rect 58532 11747 58584 11756
rect 58532 11713 58541 11747
rect 58541 11713 58575 11747
rect 58575 11713 58584 11747
rect 58532 11704 58584 11713
rect 26516 11636 26568 11688
rect 28724 11636 28776 11688
rect 30104 11636 30156 11688
rect 31576 11679 31628 11688
rect 31576 11645 31585 11679
rect 31585 11645 31619 11679
rect 31619 11645 31628 11679
rect 31576 11636 31628 11645
rect 33600 11679 33652 11688
rect 33600 11645 33609 11679
rect 33609 11645 33643 11679
rect 33643 11645 33652 11679
rect 33600 11636 33652 11645
rect 33784 11679 33836 11688
rect 33784 11645 33793 11679
rect 33793 11645 33827 11679
rect 33827 11645 33836 11679
rect 33784 11636 33836 11645
rect 34796 11679 34848 11688
rect 34796 11645 34805 11679
rect 34805 11645 34839 11679
rect 34839 11645 34848 11679
rect 34796 11636 34848 11645
rect 36084 11636 36136 11688
rect 36176 11679 36228 11688
rect 36176 11645 36185 11679
rect 36185 11645 36219 11679
rect 36219 11645 36228 11679
rect 36176 11636 36228 11645
rect 36360 11679 36412 11688
rect 36360 11645 36369 11679
rect 36369 11645 36403 11679
rect 36403 11645 36412 11679
rect 36360 11636 36412 11645
rect 37832 11679 37884 11688
rect 37832 11645 37841 11679
rect 37841 11645 37875 11679
rect 37875 11645 37884 11679
rect 37832 11636 37884 11645
rect 40868 11679 40920 11688
rect 40868 11645 40877 11679
rect 40877 11645 40911 11679
rect 40911 11645 40920 11679
rect 40868 11636 40920 11645
rect 42984 11679 43036 11688
rect 42984 11645 42993 11679
rect 42993 11645 43027 11679
rect 43027 11645 43036 11679
rect 42984 11636 43036 11645
rect 45468 11636 45520 11688
rect 45652 11679 45704 11688
rect 45652 11645 45661 11679
rect 45661 11645 45695 11679
rect 45695 11645 45704 11679
rect 45652 11636 45704 11645
rect 45928 11679 45980 11688
rect 45928 11645 45937 11679
rect 45937 11645 45971 11679
rect 45971 11645 45980 11679
rect 45928 11636 45980 11645
rect 49608 11679 49660 11688
rect 49608 11645 49617 11679
rect 49617 11645 49651 11679
rect 49651 11645 49660 11679
rect 49608 11636 49660 11645
rect 52460 11679 52512 11688
rect 52460 11645 52469 11679
rect 52469 11645 52503 11679
rect 52503 11645 52512 11679
rect 52460 11636 52512 11645
rect 53288 11679 53340 11688
rect 53288 11645 53297 11679
rect 53297 11645 53331 11679
rect 53331 11645 53340 11679
rect 53288 11636 53340 11645
rect 53748 11679 53800 11688
rect 53748 11645 53757 11679
rect 53757 11645 53791 11679
rect 53791 11645 53800 11679
rect 53748 11636 53800 11645
rect 14924 11568 14976 11620
rect 16856 11568 16908 11620
rect 20444 11568 20496 11620
rect 25412 11568 25464 11620
rect 32128 11568 32180 11620
rect 32680 11568 32732 11620
rect 36820 11568 36872 11620
rect 56508 11636 56560 11688
rect 57060 11679 57112 11688
rect 57060 11645 57069 11679
rect 57069 11645 57103 11679
rect 57103 11645 57112 11679
rect 57060 11636 57112 11645
rect 55588 11568 55640 11620
rect 56600 11611 56652 11620
rect 56600 11577 56609 11611
rect 56609 11577 56643 11611
rect 56643 11577 56652 11611
rect 56600 11568 56652 11577
rect 56876 11568 56928 11620
rect 11704 11500 11756 11552
rect 13820 11500 13872 11552
rect 13912 11500 13964 11552
rect 14372 11500 14424 11552
rect 14556 11500 14608 11552
rect 14740 11500 14792 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 18328 11500 18380 11552
rect 19524 11500 19576 11552
rect 21272 11500 21324 11552
rect 24492 11500 24544 11552
rect 25504 11500 25556 11552
rect 25964 11543 26016 11552
rect 25964 11509 25973 11543
rect 25973 11509 26007 11543
rect 26007 11509 26016 11543
rect 25964 11500 26016 11509
rect 27712 11500 27764 11552
rect 29092 11500 29144 11552
rect 30564 11500 30616 11552
rect 30840 11543 30892 11552
rect 30840 11509 30849 11543
rect 30849 11509 30883 11543
rect 30883 11509 30892 11543
rect 30840 11500 30892 11509
rect 31024 11543 31076 11552
rect 31024 11509 31033 11543
rect 31033 11509 31067 11543
rect 31067 11509 31076 11543
rect 31024 11500 31076 11509
rect 33048 11543 33100 11552
rect 33048 11509 33057 11543
rect 33057 11509 33091 11543
rect 33091 11509 33100 11543
rect 33048 11500 33100 11509
rect 34428 11543 34480 11552
rect 34428 11509 34437 11543
rect 34437 11509 34471 11543
rect 34471 11509 34480 11543
rect 34428 11500 34480 11509
rect 35624 11543 35676 11552
rect 35624 11509 35633 11543
rect 35633 11509 35667 11543
rect 35667 11509 35676 11543
rect 35624 11500 35676 11509
rect 36636 11500 36688 11552
rect 40040 11500 40092 11552
rect 42156 11500 42208 11552
rect 42800 11500 42852 11552
rect 43720 11543 43772 11552
rect 43720 11509 43729 11543
rect 43729 11509 43763 11543
rect 43763 11509 43772 11543
rect 43720 11500 43772 11509
rect 45100 11543 45152 11552
rect 45100 11509 45109 11543
rect 45109 11509 45143 11543
rect 45143 11509 45152 11543
rect 45100 11500 45152 11509
rect 45560 11500 45612 11552
rect 47308 11500 47360 11552
rect 48320 11500 48372 11552
rect 49424 11500 49476 11552
rect 50712 11500 50764 11552
rect 50988 11543 51040 11552
rect 50988 11509 50997 11543
rect 50997 11509 51031 11543
rect 51031 11509 51040 11543
rect 50988 11500 51040 11509
rect 51908 11543 51960 11552
rect 51908 11509 51917 11543
rect 51917 11509 51951 11543
rect 51951 11509 51960 11543
rect 51908 11500 51960 11509
rect 52736 11543 52788 11552
rect 52736 11509 52745 11543
rect 52745 11509 52779 11543
rect 52779 11509 52788 11543
rect 52736 11500 52788 11509
rect 56692 11500 56744 11552
rect 57428 11500 57480 11552
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 22616 11398 22668 11450
rect 22680 11398 22732 11450
rect 22744 11398 22796 11450
rect 22808 11398 22860 11450
rect 22872 11398 22924 11450
rect 37060 11398 37112 11450
rect 37124 11398 37176 11450
rect 37188 11398 37240 11450
rect 37252 11398 37304 11450
rect 37316 11398 37368 11450
rect 51504 11398 51556 11450
rect 51568 11398 51620 11450
rect 51632 11398 51684 11450
rect 51696 11398 51748 11450
rect 51760 11398 51812 11450
rect 4804 11296 4856 11348
rect 7564 11296 7616 11348
rect 7932 11296 7984 11348
rect 9956 11296 10008 11348
rect 2872 11228 2924 11280
rect 4436 11228 4488 11280
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 3424 11092 3476 11144
rect 3792 11135 3844 11144
rect 3792 11101 3821 11135
rect 3821 11101 3844 11135
rect 3792 11092 3844 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 2872 10956 2924 11008
rect 3516 10956 3568 11008
rect 3792 10956 3844 11008
rect 4252 10956 4304 11008
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 7748 11160 7800 11212
rect 6920 11092 6972 11144
rect 7288 11024 7340 11076
rect 8944 11092 8996 11144
rect 10508 11160 10560 11212
rect 11704 11296 11756 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 13360 11228 13412 11280
rect 15200 11228 15252 11280
rect 16212 11228 16264 11280
rect 16856 11228 16908 11280
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 23480 11296 23532 11348
rect 23664 11296 23716 11348
rect 24492 11296 24544 11348
rect 27528 11296 27580 11348
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11704 11160 11756 11212
rect 13544 11160 13596 11212
rect 21456 11228 21508 11280
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 11888 11092 11940 11144
rect 9956 11024 10008 11076
rect 10232 11024 10284 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 12532 11092 12584 11144
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 20352 11135 20404 11144
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 20444 11092 20496 11144
rect 6828 10999 6880 11008
rect 6828 10965 6837 10999
rect 6837 10965 6871 10999
rect 6871 10965 6880 10999
rect 6828 10956 6880 10965
rect 10968 10956 11020 11008
rect 11244 10956 11296 11008
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 19800 11067 19852 11076
rect 19800 11033 19809 11067
rect 19809 11033 19843 11067
rect 19843 11033 19852 11067
rect 19800 11024 19852 11033
rect 21180 11135 21232 11144
rect 21180 11101 21189 11135
rect 21189 11101 21223 11135
rect 21223 11101 21232 11135
rect 21180 11092 21232 11101
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 22376 11228 22428 11280
rect 23296 11228 23348 11280
rect 14372 10999 14424 11008
rect 14372 10965 14381 10999
rect 14381 10965 14415 10999
rect 14415 10965 14424 10999
rect 14372 10956 14424 10965
rect 14556 10999 14608 11008
rect 14556 10965 14565 10999
rect 14565 10965 14599 10999
rect 14599 10965 14608 10999
rect 14556 10956 14608 10965
rect 15292 10956 15344 11008
rect 17132 10956 17184 11008
rect 17684 10956 17736 11008
rect 17960 10956 18012 11008
rect 19248 10956 19300 11008
rect 20536 10956 20588 11008
rect 21548 10956 21600 11008
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 28724 11228 28776 11280
rect 28908 11228 28960 11280
rect 30104 11339 30156 11348
rect 30104 11305 30113 11339
rect 30113 11305 30147 11339
rect 30147 11305 30156 11339
rect 30104 11296 30156 11305
rect 37832 11296 37884 11348
rect 42984 11296 43036 11348
rect 44456 11339 44508 11348
rect 44456 11305 44465 11339
rect 44465 11305 44499 11339
rect 44499 11305 44508 11339
rect 44456 11296 44508 11305
rect 44640 11296 44692 11348
rect 45652 11296 45704 11348
rect 26424 11092 26476 11144
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 23204 11024 23256 11076
rect 22008 10999 22060 11008
rect 22008 10965 22017 10999
rect 22017 10965 22051 10999
rect 22051 10965 22060 10999
rect 22008 10956 22060 10965
rect 22928 10999 22980 11008
rect 22928 10965 22937 10999
rect 22937 10965 22971 10999
rect 22971 10965 22980 10999
rect 22928 10956 22980 10965
rect 23664 10956 23716 11008
rect 26516 11024 26568 11076
rect 26700 11067 26752 11076
rect 26700 11033 26709 11067
rect 26709 11033 26743 11067
rect 26743 11033 26752 11067
rect 26700 11024 26752 11033
rect 27896 11067 27948 11076
rect 27896 11033 27905 11067
rect 27905 11033 27939 11067
rect 27939 11033 27948 11067
rect 27896 11024 27948 11033
rect 29184 11024 29236 11076
rect 27252 10956 27304 11008
rect 29000 10999 29052 11008
rect 29000 10965 29009 10999
rect 29009 10965 29043 10999
rect 29043 10965 29052 10999
rect 29000 10956 29052 10965
rect 35532 11228 35584 11280
rect 37648 11228 37700 11280
rect 44180 11228 44232 11280
rect 30748 11203 30800 11212
rect 30748 11169 30757 11203
rect 30757 11169 30791 11203
rect 30791 11169 30800 11203
rect 30748 11160 30800 11169
rect 31668 11203 31720 11212
rect 31668 11169 31677 11203
rect 31677 11169 31711 11203
rect 31711 11169 31720 11203
rect 31668 11160 31720 11169
rect 30472 11067 30524 11076
rect 30472 11033 30481 11067
rect 30481 11033 30515 11067
rect 30515 11033 30524 11067
rect 30472 11024 30524 11033
rect 31024 11024 31076 11076
rect 32404 11160 32456 11212
rect 34796 11160 34848 11212
rect 35440 11160 35492 11212
rect 37740 11160 37792 11212
rect 33508 11024 33560 11076
rect 34060 11024 34112 11076
rect 34336 11067 34388 11076
rect 34336 11033 34345 11067
rect 34345 11033 34379 11067
rect 34379 11033 34388 11067
rect 34336 11024 34388 11033
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 37556 11092 37608 11144
rect 39028 11135 39080 11144
rect 39028 11101 39037 11135
rect 39037 11101 39071 11135
rect 39071 11101 39080 11135
rect 39028 11092 39080 11101
rect 39856 11203 39908 11212
rect 39856 11169 39865 11203
rect 39865 11169 39899 11203
rect 39899 11169 39908 11203
rect 39856 11160 39908 11169
rect 41604 11160 41656 11212
rect 42064 11203 42116 11212
rect 42064 11169 42073 11203
rect 42073 11169 42107 11203
rect 42107 11169 42116 11203
rect 42064 11160 42116 11169
rect 46480 11296 46532 11348
rect 48136 11296 48188 11348
rect 48780 11296 48832 11348
rect 48872 11296 48924 11348
rect 49608 11296 49660 11348
rect 50528 11296 50580 11348
rect 52368 11339 52420 11348
rect 52368 11305 52377 11339
rect 52377 11305 52411 11339
rect 52411 11305 52420 11339
rect 52368 11296 52420 11305
rect 52460 11339 52512 11348
rect 52460 11305 52469 11339
rect 52469 11305 52503 11339
rect 52503 11305 52512 11339
rect 52460 11296 52512 11305
rect 53472 11339 53524 11348
rect 53472 11305 53481 11339
rect 53481 11305 53515 11339
rect 53515 11305 53524 11339
rect 53472 11296 53524 11305
rect 47676 11271 47728 11280
rect 47676 11237 47685 11271
rect 47685 11237 47719 11271
rect 47719 11237 47728 11271
rect 47676 11228 47728 11237
rect 48228 11228 48280 11280
rect 47768 11160 47820 11212
rect 48596 11203 48648 11212
rect 48596 11169 48605 11203
rect 48605 11169 48639 11203
rect 48639 11169 48648 11203
rect 48596 11160 48648 11169
rect 35992 11024 36044 11076
rect 36820 11024 36872 11076
rect 38384 11067 38436 11076
rect 38384 11033 38393 11067
rect 38393 11033 38427 11067
rect 38427 11033 38436 11067
rect 38384 11024 38436 11033
rect 40224 11024 40276 11076
rect 41328 11135 41380 11144
rect 41328 11101 41337 11135
rect 41337 11101 41371 11135
rect 41371 11101 41380 11135
rect 41328 11092 41380 11101
rect 44088 11135 44140 11144
rect 44088 11101 44097 11135
rect 44097 11101 44131 11135
rect 44131 11101 44140 11135
rect 44088 11092 44140 11101
rect 45560 11135 45612 11144
rect 45560 11101 45569 11135
rect 45569 11101 45603 11135
rect 45603 11101 45612 11135
rect 45560 11092 45612 11101
rect 47283 11135 47335 11144
rect 47283 11101 47305 11135
rect 47305 11101 47335 11135
rect 47283 11092 47335 11101
rect 47400 11135 47452 11144
rect 47400 11101 47409 11135
rect 47409 11101 47443 11135
rect 47443 11101 47452 11135
rect 47400 11092 47452 11101
rect 52920 11203 52972 11212
rect 52920 11169 52929 11203
rect 52929 11169 52963 11203
rect 52963 11169 52972 11203
rect 52920 11160 52972 11169
rect 58440 11228 58492 11280
rect 53748 11203 53800 11212
rect 53748 11169 53757 11203
rect 53757 11169 53791 11203
rect 53791 11169 53800 11203
rect 53748 11160 53800 11169
rect 56232 11203 56284 11212
rect 56232 11169 56241 11203
rect 56241 11169 56275 11203
rect 56275 11169 56284 11203
rect 56232 11160 56284 11169
rect 49700 11092 49752 11144
rect 41788 11024 41840 11076
rect 43904 11024 43956 11076
rect 46480 11067 46532 11076
rect 46480 11033 46489 11067
rect 46489 11033 46523 11067
rect 46523 11033 46532 11067
rect 46480 11024 46532 11033
rect 55864 11135 55916 11144
rect 55864 11101 55873 11135
rect 55873 11101 55907 11135
rect 55907 11101 55916 11135
rect 55864 11092 55916 11101
rect 57336 11092 57388 11144
rect 51908 11024 51960 11076
rect 32220 10999 32272 11008
rect 32220 10965 32229 10999
rect 32229 10965 32263 10999
rect 32263 10965 32272 10999
rect 32220 10956 32272 10965
rect 35808 10956 35860 11008
rect 37924 10999 37976 11008
rect 37924 10965 37933 10999
rect 37933 10965 37967 10999
rect 37967 10965 37976 10999
rect 37924 10956 37976 10965
rect 38016 10999 38068 11008
rect 38016 10965 38025 10999
rect 38025 10965 38059 10999
rect 38059 10965 38068 10999
rect 38016 10956 38068 10965
rect 39304 10999 39356 11008
rect 39304 10965 39313 10999
rect 39313 10965 39347 10999
rect 39347 10965 39356 10999
rect 39304 10956 39356 10965
rect 41972 10999 42024 11008
rect 41972 10965 41981 10999
rect 41981 10965 42015 10999
rect 42015 10965 42024 10999
rect 41972 10956 42024 10965
rect 43536 10999 43588 11008
rect 43536 10965 43545 10999
rect 43545 10965 43579 10999
rect 43579 10965 43588 10999
rect 43536 10956 43588 10965
rect 45652 10999 45704 11008
rect 45652 10965 45661 10999
rect 45661 10965 45695 10999
rect 45695 10965 45704 10999
rect 45652 10956 45704 10965
rect 46572 10956 46624 11008
rect 47124 10956 47176 11008
rect 48688 10999 48740 11008
rect 48688 10965 48697 10999
rect 48697 10965 48731 10999
rect 48731 10965 48740 10999
rect 48688 10956 48740 10965
rect 51172 10956 51224 11008
rect 52828 10999 52880 11008
rect 52828 10965 52837 10999
rect 52837 10965 52871 10999
rect 52871 10965 52880 10999
rect 52828 10956 52880 10965
rect 55128 10999 55180 11008
rect 55128 10965 55137 10999
rect 55137 10965 55171 10999
rect 55171 10965 55180 10999
rect 55128 10956 55180 10965
rect 15394 10854 15446 10906
rect 15458 10854 15510 10906
rect 15522 10854 15574 10906
rect 15586 10854 15638 10906
rect 15650 10854 15702 10906
rect 29838 10854 29890 10906
rect 29902 10854 29954 10906
rect 29966 10854 30018 10906
rect 30030 10854 30082 10906
rect 30094 10854 30146 10906
rect 44282 10854 44334 10906
rect 44346 10854 44398 10906
rect 44410 10854 44462 10906
rect 44474 10854 44526 10906
rect 44538 10854 44590 10906
rect 58726 10854 58778 10906
rect 58790 10854 58842 10906
rect 58854 10854 58906 10906
rect 58918 10854 58970 10906
rect 58982 10854 59034 10906
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 3976 10752 4028 10804
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 3332 10616 3384 10668
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 3792 10684 3844 10736
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 7472 10752 7524 10804
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 9956 10752 10008 10804
rect 10600 10752 10652 10804
rect 10968 10752 11020 10804
rect 8576 10684 8628 10736
rect 11704 10684 11756 10736
rect 3148 10548 3200 10600
rect 3056 10480 3108 10532
rect 3792 10548 3844 10600
rect 4160 10616 4212 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 10600 10616 10652 10668
rect 11336 10616 11388 10668
rect 12072 10616 12124 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 9772 10548 9824 10600
rect 10968 10548 11020 10600
rect 11152 10548 11204 10600
rect 11428 10548 11480 10600
rect 9864 10523 9916 10532
rect 9864 10489 9873 10523
rect 9873 10489 9907 10523
rect 9907 10489 9916 10523
rect 9864 10480 9916 10489
rect 10324 10480 10376 10532
rect 15200 10752 15252 10804
rect 17500 10752 17552 10804
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 20352 10752 20404 10804
rect 21456 10752 21508 10804
rect 27988 10752 28040 10804
rect 14372 10684 14424 10736
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 16764 10616 16816 10668
rect 17960 10616 18012 10668
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 20536 10659 20588 10668
rect 20536 10625 20570 10659
rect 20570 10625 20588 10659
rect 20536 10616 20588 10625
rect 15752 10548 15804 10600
rect 15844 10591 15896 10600
rect 15844 10557 15853 10591
rect 15853 10557 15887 10591
rect 15887 10557 15896 10591
rect 15844 10548 15896 10557
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 18972 10548 19024 10600
rect 16580 10480 16632 10532
rect 3240 10412 3292 10464
rect 4068 10412 4120 10464
rect 6460 10412 6512 10464
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 10968 10412 11020 10464
rect 12532 10412 12584 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13176 10455 13228 10464
rect 13176 10421 13185 10455
rect 13185 10421 13219 10455
rect 13219 10421 13228 10455
rect 13176 10412 13228 10421
rect 14740 10412 14792 10464
rect 18144 10455 18196 10464
rect 18144 10421 18153 10455
rect 18153 10421 18187 10455
rect 18187 10421 18196 10455
rect 18144 10412 18196 10421
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 21456 10548 21508 10600
rect 22928 10616 22980 10668
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 26332 10616 26384 10668
rect 23756 10591 23808 10600
rect 23756 10557 23765 10591
rect 23765 10557 23799 10591
rect 23799 10557 23808 10591
rect 23756 10548 23808 10557
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 27620 10684 27672 10736
rect 29736 10684 29788 10736
rect 30748 10727 30800 10736
rect 30748 10693 30757 10727
rect 30757 10693 30791 10727
rect 30791 10693 30800 10727
rect 30748 10684 30800 10693
rect 27252 10616 27304 10668
rect 27712 10616 27764 10668
rect 33600 10795 33652 10804
rect 33600 10761 33609 10795
rect 33609 10761 33643 10795
rect 33643 10761 33652 10795
rect 33600 10752 33652 10761
rect 34428 10752 34480 10804
rect 35072 10752 35124 10804
rect 35716 10752 35768 10804
rect 35900 10752 35952 10804
rect 36176 10795 36228 10804
rect 36176 10761 36185 10795
rect 36185 10761 36219 10795
rect 36219 10761 36228 10795
rect 36176 10752 36228 10761
rect 36636 10795 36688 10804
rect 36636 10761 36645 10795
rect 36645 10761 36679 10795
rect 36679 10761 36688 10795
rect 36636 10752 36688 10761
rect 39304 10752 39356 10804
rect 33048 10684 33100 10736
rect 35624 10684 35676 10736
rect 37556 10684 37608 10736
rect 30932 10659 30984 10668
rect 30932 10625 30941 10659
rect 30941 10625 30975 10659
rect 30975 10625 30984 10659
rect 30932 10616 30984 10625
rect 32128 10659 32180 10668
rect 32128 10625 32137 10659
rect 32137 10625 32171 10659
rect 32171 10625 32180 10659
rect 32128 10616 32180 10625
rect 33968 10659 34020 10668
rect 33968 10625 33977 10659
rect 33977 10625 34011 10659
rect 34011 10625 34020 10659
rect 33968 10616 34020 10625
rect 34796 10616 34848 10668
rect 21272 10412 21324 10464
rect 22100 10412 22152 10464
rect 33784 10548 33836 10600
rect 36360 10548 36412 10600
rect 36544 10548 36596 10600
rect 38568 10616 38620 10668
rect 40040 10684 40092 10736
rect 40868 10795 40920 10804
rect 40868 10761 40877 10795
rect 40877 10761 40911 10795
rect 40911 10761 40920 10795
rect 40868 10752 40920 10761
rect 41328 10752 41380 10804
rect 41328 10591 41380 10600
rect 41328 10557 41337 10591
rect 41337 10557 41371 10591
rect 41371 10557 41380 10591
rect 41328 10548 41380 10557
rect 42616 10752 42668 10804
rect 43904 10795 43956 10804
rect 43904 10761 43913 10795
rect 43913 10761 43947 10795
rect 43947 10761 43956 10795
rect 43904 10752 43956 10761
rect 45928 10752 45980 10804
rect 47768 10752 47820 10804
rect 43536 10684 43588 10736
rect 45100 10684 45152 10736
rect 47400 10684 47452 10736
rect 42064 10616 42116 10668
rect 44640 10659 44692 10668
rect 44640 10625 44649 10659
rect 44649 10625 44683 10659
rect 44683 10625 44692 10659
rect 44640 10616 44692 10625
rect 45652 10616 45704 10668
rect 48688 10752 48740 10804
rect 49792 10752 49844 10804
rect 48136 10684 48188 10736
rect 48596 10727 48648 10736
rect 48596 10693 48605 10727
rect 48605 10693 48639 10727
rect 48639 10693 48648 10727
rect 52000 10752 52052 10804
rect 53380 10752 53432 10804
rect 55864 10752 55916 10804
rect 56508 10752 56560 10804
rect 57060 10752 57112 10804
rect 57336 10795 57388 10804
rect 57336 10761 57345 10795
rect 57345 10761 57379 10795
rect 57379 10761 57388 10795
rect 57336 10752 57388 10761
rect 48596 10684 48648 10693
rect 52736 10684 52788 10736
rect 44456 10591 44508 10600
rect 44456 10557 44465 10591
rect 44465 10557 44499 10591
rect 44499 10557 44508 10591
rect 44456 10548 44508 10557
rect 41972 10480 42024 10532
rect 23848 10412 23900 10464
rect 25136 10455 25188 10464
rect 25136 10421 25145 10455
rect 25145 10421 25179 10455
rect 25179 10421 25188 10455
rect 25136 10412 25188 10421
rect 27160 10412 27212 10464
rect 28540 10455 28592 10464
rect 28540 10421 28549 10455
rect 28549 10421 28583 10455
rect 28583 10421 28592 10455
rect 28540 10412 28592 10421
rect 29552 10412 29604 10464
rect 34152 10412 34204 10464
rect 38844 10455 38896 10464
rect 38844 10421 38853 10455
rect 38853 10421 38887 10455
rect 38887 10421 38896 10455
rect 38844 10412 38896 10421
rect 40776 10412 40828 10464
rect 42708 10412 42760 10464
rect 43812 10455 43864 10464
rect 43812 10421 43821 10455
rect 43821 10421 43855 10455
rect 43855 10421 43864 10455
rect 43812 10412 43864 10421
rect 46112 10455 46164 10464
rect 46112 10421 46121 10455
rect 46121 10421 46155 10455
rect 46155 10421 46164 10455
rect 46112 10412 46164 10421
rect 47952 10548 48004 10600
rect 48228 10616 48280 10668
rect 49700 10548 49752 10600
rect 49884 10659 49936 10668
rect 49884 10625 49893 10659
rect 49893 10625 49927 10659
rect 49927 10625 49936 10659
rect 49884 10616 49936 10625
rect 50528 10616 50580 10668
rect 51172 10659 51224 10668
rect 51172 10625 51181 10659
rect 51181 10625 51215 10659
rect 51215 10625 51224 10659
rect 51172 10616 51224 10625
rect 53104 10659 53156 10668
rect 53104 10625 53113 10659
rect 53113 10625 53147 10659
rect 53147 10625 53156 10659
rect 53104 10616 53156 10625
rect 50252 10591 50304 10600
rect 50252 10557 50261 10591
rect 50261 10557 50295 10591
rect 50295 10557 50304 10591
rect 50252 10548 50304 10557
rect 52736 10548 52788 10600
rect 53380 10591 53432 10600
rect 53380 10557 53389 10591
rect 53389 10557 53423 10591
rect 53423 10557 53432 10591
rect 53380 10548 53432 10557
rect 54668 10659 54720 10668
rect 54668 10625 54677 10659
rect 54677 10625 54711 10659
rect 54711 10625 54720 10659
rect 54668 10616 54720 10625
rect 56968 10616 57020 10668
rect 58440 10659 58492 10668
rect 58440 10625 58449 10659
rect 58449 10625 58483 10659
rect 58483 10625 58492 10659
rect 58440 10616 58492 10625
rect 54300 10548 54352 10600
rect 55036 10548 55088 10600
rect 55128 10548 55180 10600
rect 56784 10591 56836 10600
rect 56784 10557 56793 10591
rect 56793 10557 56827 10591
rect 56827 10557 56836 10591
rect 56784 10548 56836 10557
rect 48044 10412 48096 10464
rect 50804 10455 50856 10464
rect 50804 10421 50813 10455
rect 50813 10421 50847 10455
rect 50847 10421 50856 10455
rect 50804 10412 50856 10421
rect 53288 10412 53340 10464
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 22616 10310 22668 10362
rect 22680 10310 22732 10362
rect 22744 10310 22796 10362
rect 22808 10310 22860 10362
rect 22872 10310 22924 10362
rect 37060 10310 37112 10362
rect 37124 10310 37176 10362
rect 37188 10310 37240 10362
rect 37252 10310 37304 10362
rect 37316 10310 37368 10362
rect 51504 10310 51556 10362
rect 51568 10310 51620 10362
rect 51632 10310 51684 10362
rect 51696 10310 51748 10362
rect 51760 10310 51812 10362
rect 3332 10208 3384 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 8024 10208 8076 10260
rect 9864 10208 9916 10260
rect 10048 10208 10100 10260
rect 10232 10208 10284 10260
rect 10692 10208 10744 10260
rect 12072 10208 12124 10260
rect 13176 10208 13228 10260
rect 15844 10208 15896 10260
rect 3056 10140 3108 10192
rect 3056 9979 3108 9988
rect 3056 9945 3065 9979
rect 3065 9945 3099 9979
rect 3099 9945 3108 9979
rect 3056 9936 3108 9945
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 4252 10072 4304 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 6368 10140 6420 10192
rect 7012 10183 7064 10192
rect 7012 10149 7021 10183
rect 7021 10149 7055 10183
rect 7055 10149 7064 10183
rect 7012 10140 7064 10149
rect 8944 10183 8996 10192
rect 8944 10149 8953 10183
rect 8953 10149 8987 10183
rect 8987 10149 8996 10183
rect 8944 10140 8996 10149
rect 9404 10140 9456 10192
rect 6736 10072 6788 10124
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 6460 10004 6512 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 11888 10115 11940 10124
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 15292 10140 15344 10192
rect 16028 10140 16080 10192
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 17868 10208 17920 10260
rect 18696 10208 18748 10260
rect 21456 10251 21508 10260
rect 21456 10217 21465 10251
rect 21465 10217 21499 10251
rect 21499 10217 21508 10251
rect 21456 10208 21508 10217
rect 16764 10115 16816 10124
rect 16764 10081 16773 10115
rect 16773 10081 16807 10115
rect 16807 10081 16816 10115
rect 16764 10072 16816 10081
rect 16948 10072 17000 10124
rect 17132 10072 17184 10124
rect 10876 10004 10928 10056
rect 11704 10004 11756 10056
rect 6552 9936 6604 9988
rect 12256 9936 12308 9988
rect 16580 10004 16632 10056
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 18420 10072 18472 10124
rect 22468 10208 22520 10260
rect 26424 10208 26476 10260
rect 30932 10208 30984 10260
rect 31576 10208 31628 10260
rect 34152 10208 34204 10260
rect 36544 10208 36596 10260
rect 23572 10140 23624 10192
rect 14556 9936 14608 9988
rect 20260 10004 20312 10056
rect 22652 10072 22704 10124
rect 23112 10072 23164 10124
rect 23204 10115 23256 10124
rect 23204 10081 23213 10115
rect 23213 10081 23247 10115
rect 23247 10081 23256 10115
rect 23204 10072 23256 10081
rect 22284 10004 22336 10056
rect 23388 10047 23440 10056
rect 23388 10013 23397 10047
rect 23397 10013 23431 10047
rect 23431 10013 23440 10047
rect 23388 10004 23440 10013
rect 23664 10115 23716 10124
rect 23664 10081 23673 10115
rect 23673 10081 23707 10115
rect 23707 10081 23716 10115
rect 23664 10072 23716 10081
rect 32680 10183 32732 10192
rect 32680 10149 32689 10183
rect 32689 10149 32723 10183
rect 32723 10149 32732 10183
rect 32680 10140 32732 10149
rect 25044 10004 25096 10056
rect 25964 10004 26016 10056
rect 27160 10072 27212 10124
rect 27988 10072 28040 10124
rect 28172 10072 28224 10124
rect 29000 10072 29052 10124
rect 29736 10072 29788 10124
rect 31944 10072 31996 10124
rect 32404 10115 32456 10124
rect 32404 10081 32413 10115
rect 32413 10081 32447 10115
rect 32447 10081 32456 10115
rect 32404 10072 32456 10081
rect 37924 10140 37976 10192
rect 33968 10072 34020 10124
rect 34336 10072 34388 10124
rect 34428 10072 34480 10124
rect 35992 10072 36044 10124
rect 37372 10072 37424 10124
rect 37832 10072 37884 10124
rect 38016 10072 38068 10124
rect 38292 10115 38344 10124
rect 38292 10081 38301 10115
rect 38301 10081 38335 10115
rect 38335 10081 38344 10115
rect 38292 10072 38344 10081
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 27712 10047 27764 10056
rect 27712 10013 27730 10047
rect 27730 10013 27764 10047
rect 27712 10004 27764 10013
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 30840 10004 30892 10056
rect 32128 10047 32180 10056
rect 32128 10013 32137 10047
rect 32137 10013 32171 10047
rect 32171 10013 32180 10047
rect 32128 10004 32180 10013
rect 3332 9868 3384 9920
rect 4160 9868 4212 9920
rect 6368 9868 6420 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8760 9868 8812 9920
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 13820 9868 13872 9920
rect 17960 9868 18012 9920
rect 19892 9936 19944 9988
rect 23204 9936 23256 9988
rect 25136 9936 25188 9988
rect 34796 10004 34848 10056
rect 36912 10047 36964 10056
rect 36912 10013 36921 10047
rect 36921 10013 36955 10047
rect 36955 10013 36964 10047
rect 36912 10004 36964 10013
rect 37188 10047 37240 10056
rect 37188 10013 37197 10047
rect 37197 10013 37231 10047
rect 37231 10013 37240 10047
rect 37188 10004 37240 10013
rect 38844 10208 38896 10260
rect 42156 10208 42208 10260
rect 44456 10208 44508 10260
rect 47400 10208 47452 10260
rect 47952 10251 48004 10260
rect 47952 10217 47961 10251
rect 47961 10217 47995 10251
rect 47995 10217 48004 10251
rect 47952 10208 48004 10217
rect 48044 10208 48096 10260
rect 40776 10115 40828 10124
rect 40776 10081 40785 10115
rect 40785 10081 40819 10115
rect 40819 10081 40828 10115
rect 40776 10072 40828 10081
rect 41972 10072 42024 10124
rect 42156 10115 42208 10124
rect 42156 10081 42165 10115
rect 42165 10081 42199 10115
rect 42199 10081 42208 10115
rect 42156 10072 42208 10081
rect 42432 10115 42484 10124
rect 42432 10081 42441 10115
rect 42441 10081 42475 10115
rect 42475 10081 42484 10115
rect 42432 10072 42484 10081
rect 43260 10115 43312 10124
rect 43260 10081 43269 10115
rect 43269 10081 43303 10115
rect 43303 10081 43312 10115
rect 43260 10072 43312 10081
rect 44180 10072 44232 10124
rect 44640 10072 44692 10124
rect 45100 10072 45152 10124
rect 50252 10251 50304 10260
rect 50252 10217 50261 10251
rect 50261 10217 50295 10251
rect 50295 10217 50304 10251
rect 50252 10208 50304 10217
rect 54300 10208 54352 10260
rect 55404 10208 55456 10260
rect 56324 10251 56376 10260
rect 56324 10217 56333 10251
rect 56333 10217 56367 10251
rect 56367 10217 56376 10251
rect 56324 10208 56376 10217
rect 53104 10140 53156 10192
rect 53380 10140 53432 10192
rect 33600 9936 33652 9988
rect 35256 9936 35308 9988
rect 41880 10047 41932 10056
rect 41880 10013 41889 10047
rect 41889 10013 41923 10047
rect 41923 10013 41932 10047
rect 41880 10004 41932 10013
rect 18236 9868 18288 9920
rect 18972 9911 19024 9920
rect 18972 9877 18981 9911
rect 18981 9877 19015 9911
rect 19015 9877 19024 9911
rect 18972 9868 19024 9877
rect 20812 9911 20864 9920
rect 20812 9877 20821 9911
rect 20821 9877 20855 9911
rect 20855 9877 20864 9911
rect 20812 9868 20864 9877
rect 23664 9868 23716 9920
rect 24400 9911 24452 9920
rect 24400 9877 24409 9911
rect 24409 9877 24443 9911
rect 24443 9877 24452 9911
rect 24400 9868 24452 9877
rect 26608 9911 26660 9920
rect 26608 9877 26617 9911
rect 26617 9877 26651 9911
rect 26651 9877 26660 9911
rect 26608 9868 26660 9877
rect 28080 9868 28132 9920
rect 32956 9868 33008 9920
rect 34152 9911 34204 9920
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 34428 9868 34480 9920
rect 36084 9911 36136 9920
rect 36084 9877 36093 9911
rect 36093 9877 36127 9911
rect 36127 9877 36136 9911
rect 36084 9868 36136 9877
rect 36268 9911 36320 9920
rect 36268 9877 36277 9911
rect 36277 9877 36311 9911
rect 36311 9877 36320 9911
rect 36268 9868 36320 9877
rect 41328 9936 41380 9988
rect 43352 10004 43404 10056
rect 49700 10004 49752 10056
rect 50620 10047 50672 10056
rect 50620 10013 50629 10047
rect 50629 10013 50663 10047
rect 50663 10013 50672 10047
rect 50620 10004 50672 10013
rect 45836 9936 45888 9988
rect 48136 9936 48188 9988
rect 51724 10047 51776 10056
rect 51724 10013 51733 10047
rect 51733 10013 51767 10047
rect 51767 10013 51776 10047
rect 51724 10004 51776 10013
rect 51908 10047 51960 10056
rect 51908 10013 51926 10047
rect 51926 10013 51960 10047
rect 51908 10004 51960 10013
rect 57244 10072 57296 10124
rect 38292 9868 38344 9920
rect 38936 9911 38988 9920
rect 38936 9877 38945 9911
rect 38945 9877 38979 9911
rect 38979 9877 38988 9911
rect 38936 9868 38988 9877
rect 40500 9868 40552 9920
rect 42892 9868 42944 9920
rect 43444 9911 43496 9920
rect 43444 9877 43453 9911
rect 43453 9877 43487 9911
rect 43487 9877 43496 9911
rect 43444 9868 43496 9877
rect 47860 9868 47912 9920
rect 51172 9936 51224 9988
rect 52920 10047 52972 10056
rect 52920 10013 52929 10047
rect 52929 10013 52963 10047
rect 52963 10013 52972 10047
rect 52920 10004 52972 10013
rect 55312 9936 55364 9988
rect 52000 9868 52052 9920
rect 56968 9911 57020 9920
rect 56968 9877 56977 9911
rect 56977 9877 57011 9911
rect 57011 9877 57020 9911
rect 56968 9868 57020 9877
rect 15394 9766 15446 9818
rect 15458 9766 15510 9818
rect 15522 9766 15574 9818
rect 15586 9766 15638 9818
rect 15650 9766 15702 9818
rect 29838 9766 29890 9818
rect 29902 9766 29954 9818
rect 29966 9766 30018 9818
rect 30030 9766 30082 9818
rect 30094 9766 30146 9818
rect 44282 9766 44334 9818
rect 44346 9766 44398 9818
rect 44410 9766 44462 9818
rect 44474 9766 44526 9818
rect 44538 9766 44590 9818
rect 58726 9766 58778 9818
rect 58790 9766 58842 9818
rect 58854 9766 58906 9818
rect 58918 9766 58970 9818
rect 58982 9766 59034 9818
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 6368 9664 6420 9716
rect 10876 9664 10928 9716
rect 11704 9664 11756 9716
rect 11980 9664 12032 9716
rect 13544 9664 13596 9716
rect 15200 9664 15252 9716
rect 16028 9664 16080 9716
rect 16580 9664 16632 9716
rect 7012 9596 7064 9648
rect 6184 9528 6236 9580
rect 6368 9528 6420 9580
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 11244 9596 11296 9648
rect 11612 9596 11664 9648
rect 13728 9596 13780 9648
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 10140 9528 10192 9580
rect 11428 9528 11480 9580
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 7104 9392 7156 9444
rect 3240 9324 3292 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 8944 9324 8996 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 10048 9392 10100 9444
rect 12900 9528 12952 9580
rect 14372 9528 14424 9580
rect 18144 9596 18196 9648
rect 19800 9596 19852 9648
rect 22284 9664 22336 9716
rect 22192 9596 22244 9648
rect 22468 9664 22520 9716
rect 16948 9528 17000 9580
rect 10232 9392 10284 9444
rect 15844 9460 15896 9512
rect 16488 9460 16540 9512
rect 15476 9392 15528 9444
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 22008 9528 22060 9580
rect 24400 9596 24452 9648
rect 24768 9664 24820 9716
rect 31944 9707 31996 9716
rect 31944 9673 31953 9707
rect 31953 9673 31987 9707
rect 31987 9673 31996 9707
rect 31944 9664 31996 9673
rect 32128 9664 32180 9716
rect 21272 9392 21324 9444
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 22192 9392 22244 9444
rect 11060 9324 11112 9376
rect 13820 9324 13872 9376
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 15568 9324 15620 9376
rect 15752 9324 15804 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 17684 9324 17736 9376
rect 18052 9324 18104 9376
rect 18420 9324 18472 9376
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 20444 9324 20496 9376
rect 21180 9324 21232 9376
rect 21640 9324 21692 9376
rect 23848 9528 23900 9580
rect 25044 9571 25096 9580
rect 25044 9537 25053 9571
rect 25053 9537 25087 9571
rect 25087 9537 25096 9571
rect 25044 9528 25096 9537
rect 25596 9528 25648 9580
rect 23756 9503 23808 9512
rect 23756 9469 23765 9503
rect 23765 9469 23799 9503
rect 23799 9469 23808 9503
rect 23756 9460 23808 9469
rect 27160 9596 27212 9648
rect 27896 9571 27948 9580
rect 27896 9537 27930 9571
rect 27930 9537 27948 9571
rect 27896 9528 27948 9537
rect 29000 9528 29052 9580
rect 33600 9664 33652 9716
rect 35256 9707 35308 9716
rect 35256 9673 35265 9707
rect 35265 9673 35299 9707
rect 35299 9673 35308 9707
rect 35256 9664 35308 9673
rect 35992 9664 36044 9716
rect 38016 9664 38068 9716
rect 38568 9707 38620 9716
rect 38568 9673 38577 9707
rect 38577 9673 38611 9707
rect 38611 9673 38620 9707
rect 38568 9664 38620 9673
rect 33508 9596 33560 9648
rect 38292 9596 38344 9648
rect 40960 9664 41012 9716
rect 40224 9639 40276 9648
rect 40224 9605 40233 9639
rect 40233 9605 40267 9639
rect 40267 9605 40276 9639
rect 40224 9596 40276 9605
rect 32220 9528 32272 9580
rect 33416 9528 33468 9580
rect 34152 9528 34204 9580
rect 34704 9528 34756 9580
rect 34980 9528 35032 9580
rect 35532 9528 35584 9580
rect 36084 9571 36136 9580
rect 36084 9537 36093 9571
rect 36093 9537 36127 9571
rect 36127 9537 36136 9571
rect 36084 9528 36136 9537
rect 37648 9528 37700 9580
rect 38936 9528 38988 9580
rect 40500 9528 40552 9580
rect 41328 9664 41380 9716
rect 43444 9664 43496 9716
rect 45100 9707 45152 9716
rect 45100 9673 45109 9707
rect 45109 9673 45143 9707
rect 45143 9673 45152 9707
rect 45100 9664 45152 9673
rect 45836 9707 45888 9716
rect 45836 9673 45845 9707
rect 45845 9673 45879 9707
rect 45879 9673 45888 9707
rect 45836 9664 45888 9673
rect 49700 9707 49752 9716
rect 49700 9673 49709 9707
rect 49709 9673 49743 9707
rect 49743 9673 49752 9707
rect 49700 9664 49752 9673
rect 50620 9664 50672 9716
rect 41788 9596 41840 9648
rect 32680 9503 32732 9512
rect 32680 9469 32689 9503
rect 32689 9469 32723 9503
rect 32723 9469 32732 9503
rect 32680 9460 32732 9469
rect 37280 9392 37332 9444
rect 23388 9324 23440 9376
rect 26424 9367 26476 9376
rect 26424 9333 26433 9367
rect 26433 9333 26467 9367
rect 26467 9333 26476 9367
rect 26424 9324 26476 9333
rect 26516 9324 26568 9376
rect 27528 9324 27580 9376
rect 36728 9324 36780 9376
rect 37372 9324 37424 9376
rect 37648 9324 37700 9376
rect 40132 9324 40184 9376
rect 42432 9460 42484 9512
rect 43352 9639 43404 9648
rect 43352 9605 43361 9639
rect 43361 9605 43395 9639
rect 43395 9605 43404 9639
rect 43352 9596 43404 9605
rect 50804 9639 50856 9648
rect 50804 9605 50822 9639
rect 50822 9605 50856 9639
rect 50804 9596 50856 9605
rect 43812 9528 43864 9580
rect 46112 9528 46164 9580
rect 54668 9664 54720 9716
rect 57060 9664 57112 9716
rect 51908 9596 51960 9648
rect 47952 9460 48004 9512
rect 48136 9503 48188 9512
rect 48136 9469 48145 9503
rect 48145 9469 48179 9503
rect 48179 9469 48188 9503
rect 48136 9460 48188 9469
rect 51080 9503 51132 9512
rect 51080 9469 51089 9503
rect 51089 9469 51123 9503
rect 51123 9469 51132 9503
rect 51080 9460 51132 9469
rect 51264 9503 51316 9512
rect 51264 9469 51273 9503
rect 51273 9469 51307 9503
rect 51307 9469 51316 9503
rect 51264 9460 51316 9469
rect 51724 9528 51776 9580
rect 55588 9596 55640 9648
rect 56140 9571 56192 9580
rect 56140 9537 56149 9571
rect 56149 9537 56183 9571
rect 56183 9537 56192 9571
rect 56140 9528 56192 9537
rect 52736 9460 52788 9512
rect 53288 9503 53340 9512
rect 53288 9469 53297 9503
rect 53297 9469 53331 9503
rect 53331 9469 53340 9503
rect 53288 9460 53340 9469
rect 41604 9367 41656 9376
rect 41604 9333 41613 9367
rect 41613 9333 41647 9367
rect 41647 9333 41656 9367
rect 41604 9324 41656 9333
rect 44088 9392 44140 9444
rect 43260 9324 43312 9376
rect 47216 9367 47268 9376
rect 47216 9333 47225 9367
rect 47225 9333 47259 9367
rect 47259 9333 47268 9367
rect 47216 9324 47268 9333
rect 48044 9367 48096 9376
rect 48044 9333 48053 9367
rect 48053 9333 48087 9367
rect 48087 9333 48096 9367
rect 48044 9324 48096 9333
rect 48228 9324 48280 9376
rect 50160 9324 50212 9376
rect 51172 9392 51224 9444
rect 51724 9392 51776 9444
rect 55496 9503 55548 9512
rect 55496 9469 55505 9503
rect 55505 9469 55539 9503
rect 55539 9469 55548 9503
rect 55496 9460 55548 9469
rect 56324 9460 56376 9512
rect 57152 9392 57204 9444
rect 51908 9367 51960 9376
rect 51908 9333 51917 9367
rect 51917 9333 51951 9367
rect 51951 9333 51960 9367
rect 51908 9324 51960 9333
rect 53840 9367 53892 9376
rect 53840 9333 53849 9367
rect 53849 9333 53883 9367
rect 53883 9333 53892 9367
rect 53840 9324 53892 9333
rect 54760 9367 54812 9376
rect 54760 9333 54769 9367
rect 54769 9333 54803 9367
rect 54803 9333 54812 9367
rect 54760 9324 54812 9333
rect 56232 9324 56284 9376
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 22616 9222 22668 9274
rect 22680 9222 22732 9274
rect 22744 9222 22796 9274
rect 22808 9222 22860 9274
rect 22872 9222 22924 9274
rect 37060 9222 37112 9274
rect 37124 9222 37176 9274
rect 37188 9222 37240 9274
rect 37252 9222 37304 9274
rect 37316 9222 37368 9274
rect 51504 9222 51556 9274
rect 51568 9222 51620 9274
rect 51632 9222 51684 9274
rect 51696 9222 51748 9274
rect 51760 9222 51812 9274
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 4068 9120 4120 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 7380 9120 7432 9172
rect 7656 9120 7708 9172
rect 10048 9120 10100 9172
rect 6184 9095 6236 9104
rect 6184 9061 6193 9095
rect 6193 9061 6227 9095
rect 6227 9061 6236 9095
rect 6184 9052 6236 9061
rect 7196 9052 7248 9104
rect 3148 8984 3200 9036
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3792 8916 3844 8968
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 6920 8984 6972 9036
rect 2320 8780 2372 8832
rect 5264 8848 5316 8900
rect 8576 9052 8628 9104
rect 9220 9052 9272 9104
rect 14372 9120 14424 9172
rect 15292 9120 15344 9172
rect 12348 8984 12400 9036
rect 13820 8984 13872 9036
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 7748 8891 7800 8900
rect 7748 8857 7757 8891
rect 7757 8857 7791 8891
rect 7791 8857 7800 8891
rect 7748 8848 7800 8857
rect 6368 8780 6420 8832
rect 7656 8780 7708 8832
rect 8208 8780 8260 8832
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 8668 8891 8720 8900
rect 8668 8857 8677 8891
rect 8677 8857 8711 8891
rect 8711 8857 8720 8891
rect 8668 8848 8720 8857
rect 8760 8848 8812 8900
rect 10508 8848 10560 8900
rect 11244 8780 11296 8832
rect 12440 8848 12492 8900
rect 14464 8848 14516 8900
rect 15476 9120 15528 9172
rect 16580 9120 16632 9172
rect 16672 9120 16724 9172
rect 18236 9120 18288 9172
rect 18420 9120 18472 9172
rect 20260 9120 20312 9172
rect 20444 9120 20496 9172
rect 22284 9120 22336 9172
rect 22376 9163 22428 9172
rect 22376 9129 22385 9163
rect 22385 9129 22419 9163
rect 22419 9129 22428 9163
rect 22376 9120 22428 9129
rect 23296 9163 23348 9172
rect 23296 9129 23305 9163
rect 23305 9129 23339 9163
rect 23339 9129 23348 9163
rect 23296 9120 23348 9129
rect 23756 9120 23808 9172
rect 27804 9120 27856 9172
rect 29736 9163 29788 9172
rect 29736 9129 29745 9163
rect 29745 9129 29779 9163
rect 29779 9129 29788 9163
rect 29736 9120 29788 9129
rect 32680 9120 32732 9172
rect 34428 9163 34480 9172
rect 34428 9129 34437 9163
rect 34437 9129 34471 9163
rect 34471 9129 34480 9163
rect 34428 9120 34480 9129
rect 34796 9120 34848 9172
rect 36544 9120 36596 9172
rect 38292 9120 38344 9172
rect 38476 9163 38528 9172
rect 38476 9129 38485 9163
rect 38485 9129 38519 9163
rect 38519 9129 38528 9163
rect 38476 9120 38528 9129
rect 19892 9095 19944 9104
rect 19892 9061 19901 9095
rect 19901 9061 19935 9095
rect 19935 9061 19944 9095
rect 19892 9052 19944 9061
rect 43260 9052 43312 9104
rect 20812 9027 20864 9036
rect 20812 8993 20821 9027
rect 20821 8993 20855 9027
rect 20855 8993 20864 9027
rect 20812 8984 20864 8993
rect 22376 8984 22428 9036
rect 23388 8984 23440 9036
rect 16304 8848 16356 8900
rect 23112 8916 23164 8968
rect 16488 8848 16540 8900
rect 20628 8848 20680 8900
rect 26608 8984 26660 9036
rect 27988 8984 28040 9036
rect 28264 9027 28316 9036
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 27712 8916 27764 8968
rect 27896 8916 27948 8968
rect 28264 8993 28273 9027
rect 28273 8993 28307 9027
rect 28307 8993 28316 9027
rect 28264 8984 28316 8993
rect 28540 9027 28592 9036
rect 28540 8993 28549 9027
rect 28549 8993 28583 9027
rect 28583 8993 28592 9027
rect 28540 8984 28592 8993
rect 30472 8984 30524 9036
rect 31668 9027 31720 9036
rect 31668 8993 31677 9027
rect 31677 8993 31711 9027
rect 31711 8993 31720 9027
rect 31668 8984 31720 8993
rect 33232 8984 33284 9036
rect 34888 8984 34940 9036
rect 35992 8984 36044 9036
rect 36912 8984 36964 9036
rect 28724 8916 28776 8968
rect 32956 8959 33008 8968
rect 32956 8925 32965 8959
rect 32965 8925 32999 8959
rect 32999 8925 33008 8959
rect 32956 8916 33008 8925
rect 33324 8916 33376 8968
rect 34336 8916 34388 8968
rect 27068 8848 27120 8900
rect 28264 8848 28316 8900
rect 31944 8848 31996 8900
rect 22284 8780 22336 8832
rect 23204 8780 23256 8832
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 26332 8780 26384 8832
rect 28632 8780 28684 8832
rect 29184 8780 29236 8832
rect 31668 8780 31720 8832
rect 34612 8848 34664 8900
rect 36360 8959 36412 8968
rect 36360 8925 36369 8959
rect 36369 8925 36403 8959
rect 36403 8925 36412 8959
rect 36360 8916 36412 8925
rect 36820 8916 36872 8968
rect 39672 8916 39724 8968
rect 42248 8984 42300 9036
rect 48044 9052 48096 9104
rect 47032 9027 47084 9036
rect 47032 8993 47041 9027
rect 47041 8993 47075 9027
rect 47075 8993 47084 9027
rect 47032 8984 47084 8993
rect 47860 8984 47912 9036
rect 50068 9052 50120 9104
rect 48688 8984 48740 9036
rect 50160 9027 50212 9036
rect 50160 8993 50169 9027
rect 50169 8993 50203 9027
rect 50203 8993 50212 9027
rect 50160 8984 50212 8993
rect 45652 8916 45704 8968
rect 46296 8916 46348 8968
rect 46664 8916 46716 8968
rect 53288 9120 53340 9172
rect 55588 9163 55640 9172
rect 55588 9129 55597 9163
rect 55597 9129 55631 9163
rect 55631 9129 55640 9163
rect 55588 9120 55640 9129
rect 56232 9120 56284 9172
rect 56600 9120 56652 9172
rect 51908 8984 51960 9036
rect 37556 8848 37608 8900
rect 39488 8848 39540 8900
rect 47216 8848 47268 8900
rect 33416 8780 33468 8832
rect 34152 8780 34204 8832
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 36544 8780 36596 8832
rect 37832 8823 37884 8832
rect 37832 8789 37841 8823
rect 37841 8789 37875 8823
rect 37875 8789 37884 8823
rect 37832 8780 37884 8789
rect 44916 8780 44968 8832
rect 45376 8823 45428 8832
rect 45376 8789 45385 8823
rect 45385 8789 45419 8823
rect 45419 8789 45428 8823
rect 45376 8780 45428 8789
rect 46296 8823 46348 8832
rect 46296 8789 46305 8823
rect 46305 8789 46339 8823
rect 46339 8789 46348 8823
rect 46296 8780 46348 8789
rect 46664 8780 46716 8832
rect 47768 8780 47820 8832
rect 48228 8780 48280 8832
rect 55956 8916 56008 8968
rect 56232 8916 56284 8968
rect 57152 8916 57204 8968
rect 58440 8959 58492 8968
rect 58440 8925 58449 8959
rect 58449 8925 58483 8959
rect 58483 8925 58492 8959
rect 58440 8916 58492 8925
rect 49148 8823 49200 8832
rect 49148 8789 49157 8823
rect 49157 8789 49191 8823
rect 49191 8789 49200 8823
rect 49148 8780 49200 8789
rect 53196 8823 53248 8832
rect 53196 8789 53205 8823
rect 53205 8789 53239 8823
rect 53239 8789 53248 8823
rect 54300 8848 54352 8900
rect 57244 8848 57296 8900
rect 53196 8780 53248 8789
rect 57796 8823 57848 8832
rect 57796 8789 57805 8823
rect 57805 8789 57839 8823
rect 57839 8789 57848 8823
rect 57796 8780 57848 8789
rect 15394 8678 15446 8730
rect 15458 8678 15510 8730
rect 15522 8678 15574 8730
rect 15586 8678 15638 8730
rect 15650 8678 15702 8730
rect 29838 8678 29890 8730
rect 29902 8678 29954 8730
rect 29966 8678 30018 8730
rect 30030 8678 30082 8730
rect 30094 8678 30146 8730
rect 44282 8678 44334 8730
rect 44346 8678 44398 8730
rect 44410 8678 44462 8730
rect 44474 8678 44526 8730
rect 44538 8678 44590 8730
rect 58726 8678 58778 8730
rect 58790 8678 58842 8730
rect 58854 8678 58906 8730
rect 58918 8678 58970 8730
rect 58982 8678 59034 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 4252 8619 4304 8628
rect 4252 8585 4261 8619
rect 4261 8585 4295 8619
rect 4295 8585 4304 8619
rect 4252 8576 4304 8585
rect 7840 8576 7892 8628
rect 8484 8576 8536 8628
rect 9496 8576 9548 8628
rect 3884 8551 3936 8560
rect 3884 8517 3893 8551
rect 3893 8517 3927 8551
rect 3927 8517 3936 8551
rect 3884 8508 3936 8517
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 5264 8440 5316 8492
rect 6368 8440 6420 8492
rect 6736 8508 6788 8560
rect 8208 8508 8260 8560
rect 7196 8440 7248 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 9864 8508 9916 8560
rect 10048 8576 10100 8628
rect 10968 8576 11020 8628
rect 11060 8508 11112 8560
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 6184 8372 6236 8424
rect 8944 8440 8996 8492
rect 12348 8576 12400 8628
rect 14280 8576 14332 8628
rect 15844 8576 15896 8628
rect 16212 8576 16264 8628
rect 17776 8576 17828 8628
rect 18052 8576 18104 8628
rect 20260 8576 20312 8628
rect 21548 8576 21600 8628
rect 25228 8576 25280 8628
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 27160 8576 27212 8628
rect 27712 8576 27764 8628
rect 27896 8619 27948 8628
rect 27896 8585 27905 8619
rect 27905 8585 27939 8619
rect 27939 8585 27948 8619
rect 27896 8576 27948 8585
rect 7840 8372 7892 8424
rect 7656 8236 7708 8288
rect 10232 8372 10284 8424
rect 10508 8372 10560 8424
rect 10876 8372 10928 8424
rect 14188 8508 14240 8560
rect 12808 8440 12860 8492
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 33048 8508 33100 8560
rect 34888 8508 34940 8560
rect 35808 8551 35860 8560
rect 35808 8517 35817 8551
rect 35817 8517 35851 8551
rect 35851 8517 35860 8551
rect 35808 8508 35860 8517
rect 35992 8508 36044 8560
rect 36176 8508 36228 8560
rect 13268 8440 13320 8449
rect 14188 8372 14240 8424
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 16120 8440 16172 8492
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 25504 8440 25556 8449
rect 25780 8440 25832 8492
rect 26424 8440 26476 8492
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 18328 8372 18380 8424
rect 8576 8236 8628 8288
rect 10876 8236 10928 8288
rect 13820 8304 13872 8356
rect 14464 8304 14516 8356
rect 21180 8372 21232 8424
rect 22100 8347 22152 8356
rect 22100 8313 22109 8347
rect 22109 8313 22143 8347
rect 22143 8313 22152 8347
rect 22100 8304 22152 8313
rect 22468 8372 22520 8424
rect 23388 8415 23440 8424
rect 23388 8381 23397 8415
rect 23397 8381 23431 8415
rect 23431 8381 23440 8415
rect 23388 8372 23440 8381
rect 28908 8372 28960 8424
rect 30104 8372 30156 8424
rect 25964 8304 26016 8356
rect 30472 8304 30524 8356
rect 30656 8415 30708 8424
rect 30656 8381 30665 8415
rect 30665 8381 30699 8415
rect 30699 8381 30708 8415
rect 30656 8372 30708 8381
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 31944 8304 31996 8356
rect 16304 8236 16356 8288
rect 17592 8236 17644 8288
rect 21824 8236 21876 8288
rect 22376 8236 22428 8288
rect 24768 8236 24820 8288
rect 26148 8236 26200 8288
rect 27436 8236 27488 8288
rect 28724 8236 28776 8288
rect 30288 8236 30340 8288
rect 30932 8236 30984 8288
rect 32680 8279 32732 8288
rect 32680 8245 32689 8279
rect 32689 8245 32723 8279
rect 32723 8245 32732 8279
rect 34336 8483 34388 8492
rect 34336 8449 34345 8483
rect 34345 8449 34379 8483
rect 34379 8449 34388 8483
rect 34336 8440 34388 8449
rect 34520 8483 34572 8492
rect 34520 8449 34529 8483
rect 34529 8449 34563 8483
rect 34563 8449 34572 8483
rect 34520 8440 34572 8449
rect 33232 8372 33284 8424
rect 33416 8372 33468 8424
rect 33876 8304 33928 8356
rect 35164 8347 35216 8356
rect 35164 8313 35173 8347
rect 35173 8313 35207 8347
rect 35207 8313 35216 8347
rect 35164 8304 35216 8313
rect 36452 8440 36504 8492
rect 37004 8440 37056 8492
rect 44916 8508 44968 8560
rect 40408 8483 40460 8492
rect 40408 8449 40417 8483
rect 40417 8449 40451 8483
rect 40451 8449 40460 8483
rect 40408 8440 40460 8449
rect 42984 8440 43036 8492
rect 45376 8576 45428 8628
rect 48136 8576 48188 8628
rect 49148 8576 49200 8628
rect 51264 8576 51316 8628
rect 52184 8576 52236 8628
rect 54760 8576 54812 8628
rect 55496 8576 55548 8628
rect 35440 8372 35492 8424
rect 37096 8372 37148 8424
rect 37556 8372 37608 8424
rect 37924 8372 37976 8424
rect 36912 8304 36964 8356
rect 37004 8304 37056 8356
rect 32680 8236 32732 8245
rect 37096 8236 37148 8288
rect 38936 8372 38988 8424
rect 39120 8415 39172 8424
rect 39120 8381 39129 8415
rect 39129 8381 39163 8415
rect 39163 8381 39172 8415
rect 39120 8372 39172 8381
rect 43076 8415 43128 8424
rect 43076 8381 43085 8415
rect 43085 8381 43119 8415
rect 43119 8381 43128 8415
rect 43076 8372 43128 8381
rect 44732 8415 44784 8424
rect 44732 8381 44741 8415
rect 44741 8381 44775 8415
rect 44775 8381 44784 8415
rect 44732 8372 44784 8381
rect 40224 8304 40276 8356
rect 40500 8304 40552 8356
rect 39304 8279 39356 8288
rect 39304 8245 39313 8279
rect 39313 8245 39347 8279
rect 39347 8245 39356 8279
rect 39304 8236 39356 8245
rect 42064 8236 42116 8288
rect 42432 8279 42484 8288
rect 42432 8245 42441 8279
rect 42441 8245 42475 8279
rect 42475 8245 42484 8279
rect 42432 8236 42484 8245
rect 43904 8236 43956 8288
rect 44180 8304 44232 8356
rect 46296 8440 46348 8492
rect 47676 8508 47728 8560
rect 50160 8372 50212 8424
rect 50436 8415 50488 8424
rect 50436 8381 50445 8415
rect 50445 8381 50479 8415
rect 50479 8381 50488 8415
rect 50436 8372 50488 8381
rect 51908 8440 51960 8492
rect 53656 8440 53708 8492
rect 56784 8576 56836 8628
rect 57152 8576 57204 8628
rect 57244 8576 57296 8628
rect 54300 8440 54352 8492
rect 56140 8440 56192 8492
rect 53380 8415 53432 8424
rect 53380 8381 53389 8415
rect 53389 8381 53423 8415
rect 53423 8381 53432 8415
rect 53380 8372 53432 8381
rect 55680 8372 55732 8424
rect 56508 8372 56560 8424
rect 55312 8347 55364 8356
rect 55312 8313 55321 8347
rect 55321 8313 55355 8347
rect 55355 8313 55364 8347
rect 55312 8304 55364 8313
rect 46480 8236 46532 8288
rect 49884 8279 49936 8288
rect 49884 8245 49893 8279
rect 49893 8245 49927 8279
rect 49927 8245 49936 8279
rect 49884 8236 49936 8245
rect 50068 8236 50120 8288
rect 52644 8236 52696 8288
rect 52828 8279 52880 8288
rect 52828 8245 52837 8279
rect 52837 8245 52871 8279
rect 52871 8245 52880 8279
rect 52828 8236 52880 8245
rect 56876 8304 56928 8356
rect 57888 8372 57940 8424
rect 58164 8304 58216 8356
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 22616 8134 22668 8186
rect 22680 8134 22732 8186
rect 22744 8134 22796 8186
rect 22808 8134 22860 8186
rect 22872 8134 22924 8186
rect 37060 8134 37112 8186
rect 37124 8134 37176 8186
rect 37188 8134 37240 8186
rect 37252 8134 37304 8186
rect 37316 8134 37368 8186
rect 51504 8134 51556 8186
rect 51568 8134 51620 8186
rect 51632 8134 51684 8186
rect 51696 8134 51748 8186
rect 51760 8134 51812 8186
rect 3516 8032 3568 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8576 8032 8628 8084
rect 3792 8007 3844 8016
rect 3792 7973 3801 8007
rect 3801 7973 3835 8007
rect 3835 7973 3844 8007
rect 3792 7964 3844 7973
rect 13268 8032 13320 8084
rect 15752 8032 15804 8084
rect 19432 8032 19484 8084
rect 20996 8075 21048 8084
rect 20996 8041 21005 8075
rect 21005 8041 21039 8075
rect 21039 8041 21048 8075
rect 20996 8032 21048 8041
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 10508 7964 10560 8016
rect 22468 8032 22520 8084
rect 23020 8032 23072 8084
rect 23480 8032 23532 8084
rect 24768 8032 24820 8084
rect 25136 8032 25188 8084
rect 25872 8032 25924 8084
rect 3700 7828 3752 7880
rect 3792 7692 3844 7744
rect 7840 7896 7892 7948
rect 10968 7896 11020 7948
rect 5264 7828 5316 7880
rect 6184 7828 6236 7880
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6920 7828 6972 7880
rect 7288 7828 7340 7880
rect 8668 7828 8720 7880
rect 10416 7828 10468 7880
rect 8116 7760 8168 7812
rect 6092 7692 6144 7744
rect 7656 7692 7708 7744
rect 11060 7760 11112 7812
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 15476 7896 15528 7948
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 17684 7896 17736 7948
rect 18052 7896 18104 7948
rect 18512 7896 18564 7948
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 14004 7828 14056 7880
rect 14188 7828 14240 7880
rect 15200 7828 15252 7880
rect 15016 7760 15068 7812
rect 16672 7803 16724 7812
rect 16672 7769 16681 7803
rect 16681 7769 16715 7803
rect 16715 7769 16724 7803
rect 16672 7760 16724 7769
rect 16948 7760 17000 7812
rect 17960 7828 18012 7880
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 12992 7692 13044 7744
rect 15752 7692 15804 7744
rect 16304 7692 16356 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 20168 7692 20220 7744
rect 20812 7760 20864 7812
rect 24860 8007 24912 8016
rect 24860 7973 24869 8007
rect 24869 7973 24903 8007
rect 24903 7973 24912 8007
rect 24860 7964 24912 7973
rect 28908 8032 28960 8084
rect 29644 8032 29696 8084
rect 30656 8032 30708 8084
rect 25780 7896 25832 7948
rect 25964 7896 26016 7948
rect 26148 7939 26200 7948
rect 26148 7905 26157 7939
rect 26157 7905 26191 7939
rect 26191 7905 26200 7939
rect 26148 7896 26200 7905
rect 22376 7871 22428 7880
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 25596 7871 25648 7880
rect 25596 7837 25605 7871
rect 25605 7837 25639 7871
rect 25639 7837 25648 7871
rect 25596 7828 25648 7837
rect 26976 7828 27028 7880
rect 27988 7939 28040 7948
rect 27988 7905 27997 7939
rect 27997 7905 28031 7939
rect 28031 7905 28040 7939
rect 27988 7896 28040 7905
rect 30748 7964 30800 8016
rect 28540 7828 28592 7880
rect 29644 7896 29696 7948
rect 35440 8032 35492 8084
rect 36176 8075 36228 8084
rect 36176 8041 36185 8075
rect 36185 8041 36219 8075
rect 36219 8041 36228 8075
rect 36176 8032 36228 8041
rect 36360 8032 36412 8084
rect 39120 8032 39172 8084
rect 33232 7964 33284 8016
rect 44732 8032 44784 8084
rect 31760 7896 31812 7948
rect 32312 7939 32364 7948
rect 32312 7905 32321 7939
rect 32321 7905 32355 7939
rect 32355 7905 32364 7939
rect 32312 7896 32364 7905
rect 42984 7896 43036 7948
rect 45284 7964 45336 8016
rect 47676 7964 47728 8016
rect 49792 7964 49844 8016
rect 30472 7828 30524 7880
rect 23940 7760 23992 7812
rect 25044 7803 25096 7812
rect 25044 7769 25053 7803
rect 25053 7769 25087 7803
rect 25087 7769 25096 7803
rect 25044 7760 25096 7769
rect 26424 7803 26476 7812
rect 22008 7692 22060 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 23204 7692 23256 7744
rect 26424 7769 26433 7803
rect 26433 7769 26467 7803
rect 26467 7769 26476 7803
rect 26424 7760 26476 7769
rect 28632 7760 28684 7812
rect 30932 7760 30984 7812
rect 31944 7871 31996 7880
rect 31944 7837 31953 7871
rect 31953 7837 31987 7871
rect 31987 7837 31996 7871
rect 31944 7828 31996 7837
rect 32312 7760 32364 7812
rect 26332 7735 26384 7744
rect 26332 7701 26341 7735
rect 26341 7701 26375 7735
rect 26375 7701 26384 7735
rect 26332 7692 26384 7701
rect 26608 7692 26660 7744
rect 26792 7735 26844 7744
rect 26792 7701 26801 7735
rect 26801 7701 26835 7735
rect 26835 7701 26844 7735
rect 26792 7692 26844 7701
rect 26884 7692 26936 7744
rect 30104 7692 30156 7744
rect 30564 7692 30616 7744
rect 30748 7692 30800 7744
rect 34888 7828 34940 7880
rect 39120 7871 39172 7880
rect 39120 7837 39129 7871
rect 39129 7837 39163 7871
rect 39163 7837 39172 7871
rect 39120 7828 39172 7837
rect 39304 7828 39356 7880
rect 41052 7871 41104 7880
rect 41052 7837 41061 7871
rect 41061 7837 41095 7871
rect 41095 7837 41104 7871
rect 41052 7828 41104 7837
rect 35256 7760 35308 7812
rect 36360 7760 36412 7812
rect 36544 7760 36596 7812
rect 37832 7760 37884 7812
rect 40960 7760 41012 7812
rect 41512 7828 41564 7880
rect 42432 7760 42484 7812
rect 47768 7939 47820 7948
rect 47768 7905 47777 7939
rect 47777 7905 47811 7939
rect 47811 7905 47820 7939
rect 47768 7896 47820 7905
rect 50436 8032 50488 8084
rect 51080 8032 51132 8084
rect 51356 8032 51408 8084
rect 45376 7871 45428 7880
rect 45376 7837 45385 7871
rect 45385 7837 45419 7871
rect 45419 7837 45428 7871
rect 45376 7828 45428 7837
rect 46756 7871 46808 7880
rect 46756 7837 46765 7871
rect 46765 7837 46799 7871
rect 46799 7837 46808 7871
rect 46756 7828 46808 7837
rect 46848 7828 46900 7880
rect 47032 7871 47084 7880
rect 47032 7837 47041 7871
rect 47041 7837 47075 7871
rect 47075 7837 47084 7871
rect 47032 7828 47084 7837
rect 47952 7871 48004 7880
rect 47952 7837 47961 7871
rect 47961 7837 47995 7871
rect 47995 7837 48004 7871
rect 47952 7828 48004 7837
rect 48412 7871 48464 7880
rect 48412 7837 48421 7871
rect 48421 7837 48455 7871
rect 48455 7837 48464 7871
rect 48412 7828 48464 7837
rect 45836 7760 45888 7812
rect 36176 7692 36228 7744
rect 38752 7692 38804 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 40500 7735 40552 7744
rect 40500 7701 40509 7735
rect 40509 7701 40543 7735
rect 40543 7701 40552 7735
rect 40500 7692 40552 7701
rect 41788 7692 41840 7744
rect 42340 7692 42392 7744
rect 42984 7692 43036 7744
rect 44640 7692 44692 7744
rect 45560 7692 45612 7744
rect 50988 7871 51040 7880
rect 50988 7837 50997 7871
rect 50997 7837 51031 7871
rect 51031 7837 51040 7871
rect 50988 7828 51040 7837
rect 51356 7760 51408 7812
rect 52276 7939 52328 7948
rect 52276 7905 52285 7939
rect 52285 7905 52319 7939
rect 52319 7905 52328 7939
rect 52276 7896 52328 7905
rect 52644 7939 52696 7948
rect 52644 7905 52653 7939
rect 52653 7905 52687 7939
rect 52687 7905 52696 7939
rect 52644 7896 52696 7905
rect 52828 7871 52880 7880
rect 52828 7837 52837 7871
rect 52837 7837 52871 7871
rect 52871 7837 52880 7871
rect 52828 7828 52880 7837
rect 57888 8032 57940 8084
rect 58440 8032 58492 8084
rect 57888 7896 57940 7948
rect 54300 7828 54352 7880
rect 53748 7760 53800 7812
rect 54208 7760 54260 7812
rect 48044 7735 48096 7744
rect 48044 7701 48053 7735
rect 48053 7701 48087 7735
rect 48087 7701 48096 7735
rect 48044 7692 48096 7701
rect 48596 7692 48648 7744
rect 50620 7735 50672 7744
rect 50620 7701 50629 7735
rect 50629 7701 50663 7735
rect 50663 7701 50672 7735
rect 50620 7692 50672 7701
rect 52736 7735 52788 7744
rect 52736 7701 52745 7735
rect 52745 7701 52779 7735
rect 52779 7701 52788 7735
rect 52736 7692 52788 7701
rect 56232 7828 56284 7880
rect 56600 7871 56652 7880
rect 56600 7837 56634 7871
rect 56634 7837 56652 7871
rect 56600 7828 56652 7837
rect 58164 7871 58216 7880
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 55036 7760 55088 7812
rect 55128 7735 55180 7744
rect 55128 7701 55137 7735
rect 55137 7701 55171 7735
rect 55171 7701 55180 7735
rect 55128 7692 55180 7701
rect 57060 7692 57112 7744
rect 15394 7590 15446 7642
rect 15458 7590 15510 7642
rect 15522 7590 15574 7642
rect 15586 7590 15638 7642
rect 15650 7590 15702 7642
rect 29838 7590 29890 7642
rect 29902 7590 29954 7642
rect 29966 7590 30018 7642
rect 30030 7590 30082 7642
rect 30094 7590 30146 7642
rect 44282 7590 44334 7642
rect 44346 7590 44398 7642
rect 44410 7590 44462 7642
rect 44474 7590 44526 7642
rect 44538 7590 44590 7642
rect 58726 7590 58778 7642
rect 58790 7590 58842 7642
rect 58854 7590 58906 7642
rect 58918 7590 58970 7642
rect 58982 7590 59034 7642
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 6368 7488 6420 7540
rect 7564 7488 7616 7540
rect 9404 7488 9456 7540
rect 9772 7488 9824 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 10508 7420 10560 7472
rect 5448 7352 5500 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7380 7352 7432 7404
rect 5540 7284 5592 7336
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 7840 7352 7892 7404
rect 8116 7352 8168 7404
rect 8760 7284 8812 7336
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 3792 7216 3844 7268
rect 7656 7216 7708 7268
rect 10876 7284 10928 7336
rect 11244 7488 11296 7540
rect 12992 7488 13044 7540
rect 14004 7488 14056 7540
rect 14556 7488 14608 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 15752 7488 15804 7540
rect 15936 7488 15988 7540
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 12532 7420 12584 7472
rect 12808 7463 12860 7472
rect 12808 7429 12817 7463
rect 12817 7429 12851 7463
rect 12851 7429 12860 7463
rect 12808 7420 12860 7429
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 12164 7284 12216 7336
rect 12440 7284 12492 7336
rect 15384 7352 15436 7404
rect 16948 7352 17000 7404
rect 18236 7352 18288 7404
rect 20168 7531 20220 7540
rect 20168 7497 20177 7531
rect 20177 7497 20211 7531
rect 20211 7497 20220 7531
rect 20168 7488 20220 7497
rect 21916 7488 21968 7540
rect 23848 7488 23900 7540
rect 25596 7488 25648 7540
rect 26424 7488 26476 7540
rect 20536 7420 20588 7472
rect 21272 7352 21324 7404
rect 24676 7420 24728 7472
rect 26792 7420 26844 7472
rect 8852 7148 8904 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 15292 7284 15344 7336
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 20352 7327 20404 7336
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 24952 7352 25004 7404
rect 27528 7352 27580 7404
rect 27988 7352 28040 7404
rect 28724 7395 28776 7404
rect 28724 7361 28742 7395
rect 28742 7361 28776 7395
rect 28724 7352 28776 7361
rect 31392 7488 31444 7540
rect 36268 7488 36320 7540
rect 36360 7531 36412 7540
rect 36360 7497 36369 7531
rect 36369 7497 36403 7531
rect 36403 7497 36412 7531
rect 36360 7488 36412 7497
rect 37924 7488 37976 7540
rect 39120 7488 39172 7540
rect 40500 7488 40552 7540
rect 40960 7531 41012 7540
rect 40960 7497 40969 7531
rect 40969 7497 41003 7531
rect 41003 7497 41012 7531
rect 40960 7488 41012 7497
rect 41052 7531 41104 7540
rect 41052 7497 41061 7531
rect 41061 7497 41095 7531
rect 41095 7497 41104 7531
rect 41052 7488 41104 7497
rect 41420 7488 41472 7540
rect 42984 7488 43036 7540
rect 43076 7488 43128 7540
rect 45652 7531 45704 7540
rect 45652 7497 45661 7531
rect 45661 7497 45695 7531
rect 45695 7497 45704 7531
rect 45652 7488 45704 7497
rect 45836 7488 45888 7540
rect 47216 7488 47268 7540
rect 47860 7488 47912 7540
rect 50988 7488 51040 7540
rect 52000 7488 52052 7540
rect 53380 7488 53432 7540
rect 30288 7420 30340 7472
rect 32220 7352 32272 7404
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 16672 7148 16724 7200
rect 17408 7148 17460 7200
rect 17684 7148 17736 7200
rect 19340 7148 19392 7200
rect 20996 7148 21048 7200
rect 23020 7284 23072 7336
rect 23940 7327 23992 7336
rect 23940 7293 23949 7327
rect 23949 7293 23983 7327
rect 23983 7293 23992 7327
rect 23940 7284 23992 7293
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24400 7284 24452 7293
rect 22468 7148 22520 7200
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 25872 7148 25924 7200
rect 31852 7327 31904 7336
rect 31852 7293 31861 7327
rect 31861 7293 31895 7327
rect 31895 7293 31904 7327
rect 31852 7284 31904 7293
rect 33600 7395 33652 7404
rect 33600 7361 33609 7395
rect 33609 7361 33643 7395
rect 33643 7361 33652 7395
rect 33600 7352 33652 7361
rect 33876 7352 33928 7404
rect 33692 7284 33744 7336
rect 29092 7191 29144 7200
rect 29092 7157 29101 7191
rect 29101 7157 29135 7191
rect 29135 7157 29144 7191
rect 29092 7148 29144 7157
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 33508 7191 33560 7200
rect 33508 7157 33517 7191
rect 33517 7157 33551 7191
rect 33551 7157 33560 7191
rect 33508 7148 33560 7157
rect 35072 7327 35124 7336
rect 35072 7293 35081 7327
rect 35081 7293 35115 7327
rect 35115 7293 35124 7327
rect 35072 7284 35124 7293
rect 36176 7327 36228 7336
rect 36176 7293 36185 7327
rect 36185 7293 36219 7327
rect 36219 7293 36228 7327
rect 36176 7284 36228 7293
rect 36820 7259 36872 7268
rect 36820 7225 36829 7259
rect 36829 7225 36863 7259
rect 36863 7225 36872 7259
rect 36820 7216 36872 7225
rect 37924 7327 37976 7336
rect 37924 7293 37933 7327
rect 37933 7293 37967 7327
rect 37967 7293 37976 7327
rect 37924 7284 37976 7293
rect 42064 7420 42116 7472
rect 42248 7463 42300 7472
rect 42248 7429 42257 7463
rect 42257 7429 42291 7463
rect 42291 7429 42300 7463
rect 42248 7420 42300 7429
rect 42524 7420 42576 7472
rect 41788 7352 41840 7404
rect 41052 7284 41104 7336
rect 41696 7327 41748 7336
rect 41696 7293 41705 7327
rect 41705 7293 41739 7327
rect 41739 7293 41748 7327
rect 41696 7284 41748 7293
rect 42892 7352 42944 7404
rect 45928 7420 45980 7472
rect 47032 7420 47084 7472
rect 44272 7352 44324 7404
rect 45560 7352 45612 7404
rect 46388 7352 46440 7404
rect 46756 7352 46808 7404
rect 49884 7420 49936 7472
rect 54300 7488 54352 7540
rect 54668 7488 54720 7540
rect 55036 7488 55088 7540
rect 55128 7488 55180 7540
rect 43904 7327 43956 7336
rect 43904 7293 43913 7327
rect 43913 7293 43947 7327
rect 43947 7293 43956 7327
rect 43904 7284 43956 7293
rect 38844 7216 38896 7268
rect 39212 7148 39264 7200
rect 39304 7191 39356 7200
rect 39304 7157 39313 7191
rect 39313 7157 39347 7191
rect 39347 7157 39356 7191
rect 39304 7148 39356 7157
rect 41696 7148 41748 7200
rect 42064 7148 42116 7200
rect 43168 7148 43220 7200
rect 43260 7191 43312 7200
rect 43260 7157 43269 7191
rect 43269 7157 43303 7191
rect 43303 7157 43312 7191
rect 43260 7148 43312 7157
rect 46296 7327 46348 7336
rect 46296 7293 46305 7327
rect 46305 7293 46339 7327
rect 46339 7293 46348 7327
rect 46296 7284 46348 7293
rect 46480 7327 46532 7336
rect 46480 7293 46489 7327
rect 46489 7293 46523 7327
rect 46523 7293 46532 7327
rect 46480 7284 46532 7293
rect 48596 7352 48648 7404
rect 45560 7191 45612 7200
rect 45560 7157 45569 7191
rect 45569 7157 45603 7191
rect 45603 7157 45612 7191
rect 45560 7148 45612 7157
rect 51264 7284 51316 7336
rect 50160 7148 50212 7200
rect 50896 7191 50948 7200
rect 50896 7157 50905 7191
rect 50905 7157 50939 7191
rect 50939 7157 50948 7191
rect 50896 7148 50948 7157
rect 52000 7284 52052 7336
rect 54116 7395 54168 7404
rect 54116 7361 54125 7395
rect 54125 7361 54159 7395
rect 54159 7361 54168 7395
rect 54116 7352 54168 7361
rect 54852 7327 54904 7336
rect 54852 7293 54861 7327
rect 54861 7293 54895 7327
rect 54895 7293 54904 7327
rect 54852 7284 54904 7293
rect 56508 7488 56560 7540
rect 56692 7531 56744 7540
rect 56692 7497 56701 7531
rect 56701 7497 56735 7531
rect 56735 7497 56744 7531
rect 56692 7488 56744 7497
rect 56784 7531 56836 7540
rect 56784 7497 56793 7531
rect 56793 7497 56827 7531
rect 56827 7497 56836 7531
rect 56784 7488 56836 7497
rect 57888 7488 57940 7540
rect 58164 7488 58216 7540
rect 57796 7352 57848 7404
rect 57704 7284 57756 7336
rect 52276 7148 52328 7200
rect 53932 7148 53984 7200
rect 54300 7191 54352 7200
rect 54300 7157 54309 7191
rect 54309 7157 54343 7191
rect 54343 7157 54352 7191
rect 54300 7148 54352 7157
rect 56324 7191 56376 7200
rect 56324 7157 56333 7191
rect 56333 7157 56367 7191
rect 56367 7157 56376 7191
rect 56324 7148 56376 7157
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 22616 7046 22668 7098
rect 22680 7046 22732 7098
rect 22744 7046 22796 7098
rect 22808 7046 22860 7098
rect 22872 7046 22924 7098
rect 37060 7046 37112 7098
rect 37124 7046 37176 7098
rect 37188 7046 37240 7098
rect 37252 7046 37304 7098
rect 37316 7046 37368 7098
rect 51504 7046 51556 7098
rect 51568 7046 51620 7098
rect 51632 7046 51684 7098
rect 51696 7046 51748 7098
rect 51760 7046 51812 7098
rect 7380 6944 7432 6996
rect 10600 6944 10652 6996
rect 3056 6808 3108 6860
rect 5448 6808 5500 6860
rect 5816 6808 5868 6860
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6092 6851 6144 6860
rect 6092 6817 6126 6851
rect 6126 6817 6144 6851
rect 6092 6808 6144 6817
rect 7656 6808 7708 6860
rect 9772 6808 9824 6860
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3240 6740 3292 6792
rect 3516 6740 3568 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 4344 6740 4396 6792
rect 3424 6672 3476 6724
rect 3884 6672 3936 6724
rect 5632 6672 5684 6724
rect 6552 6672 6604 6724
rect 1952 6604 2004 6656
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 5540 6604 5592 6656
rect 7104 6740 7156 6792
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11244 6944 11296 6996
rect 12256 6944 12308 6996
rect 15200 6944 15252 6996
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 10968 6808 11020 6860
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12164 6808 12216 6860
rect 8024 6672 8076 6724
rect 10600 6672 10652 6724
rect 10968 6672 11020 6724
rect 11336 6715 11388 6724
rect 11336 6681 11345 6715
rect 11345 6681 11379 6715
rect 11379 6681 11388 6715
rect 11336 6672 11388 6681
rect 12164 6672 12216 6724
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 14372 6740 14424 6792
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15476 6808 15528 6860
rect 16120 6808 16172 6860
rect 18236 6944 18288 6996
rect 20720 6944 20772 6996
rect 20996 6944 21048 6996
rect 21640 6944 21692 6996
rect 22468 6944 22520 6996
rect 23020 6944 23072 6996
rect 24400 6944 24452 6996
rect 16304 6808 16356 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 17684 6808 17736 6860
rect 18328 6808 18380 6860
rect 19064 6808 19116 6860
rect 11796 6604 11848 6656
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 13912 6647 13964 6656
rect 13912 6613 13921 6647
rect 13921 6613 13955 6647
rect 13955 6613 13964 6647
rect 13912 6604 13964 6613
rect 14004 6604 14056 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 18052 6740 18104 6792
rect 17868 6715 17920 6724
rect 17868 6681 17877 6715
rect 17877 6681 17911 6715
rect 17911 6681 17920 6715
rect 17868 6672 17920 6681
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 19340 6740 19392 6792
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 21732 6740 21784 6792
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22560 6808 22612 6860
rect 23204 6808 23256 6860
rect 23480 6851 23532 6860
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23480 6808 23532 6817
rect 23940 6808 23992 6860
rect 26332 6808 26384 6860
rect 26608 6808 26660 6860
rect 26792 6808 26844 6860
rect 26976 6808 27028 6860
rect 27620 6808 27672 6860
rect 28540 6944 28592 6996
rect 32588 6944 32640 6996
rect 33600 6944 33652 6996
rect 27988 6808 28040 6860
rect 31944 6808 31996 6860
rect 33324 6876 33376 6928
rect 34152 6876 34204 6928
rect 35072 6876 35124 6928
rect 36728 6876 36780 6928
rect 37924 6944 37976 6996
rect 41052 6987 41104 6996
rect 41052 6953 41061 6987
rect 41061 6953 41095 6987
rect 41095 6953 41104 6987
rect 41052 6944 41104 6953
rect 33692 6808 33744 6860
rect 25780 6740 25832 6792
rect 25872 6783 25924 6792
rect 25872 6749 25881 6783
rect 25881 6749 25915 6783
rect 25915 6749 25924 6783
rect 25872 6740 25924 6749
rect 27160 6783 27212 6792
rect 27160 6749 27169 6783
rect 27169 6749 27203 6783
rect 27203 6749 27212 6783
rect 27160 6740 27212 6749
rect 28080 6740 28132 6792
rect 31300 6740 31352 6792
rect 31484 6740 31536 6792
rect 32312 6783 32364 6792
rect 32312 6749 32330 6783
rect 32330 6749 32364 6783
rect 32312 6740 32364 6749
rect 32404 6783 32456 6792
rect 32404 6749 32413 6783
rect 32413 6749 32447 6783
rect 32447 6749 32456 6783
rect 32404 6740 32456 6749
rect 33140 6783 33192 6792
rect 33140 6749 33149 6783
rect 33149 6749 33183 6783
rect 33183 6749 33192 6783
rect 33140 6740 33192 6749
rect 33324 6783 33376 6792
rect 33324 6749 33333 6783
rect 33333 6749 33367 6783
rect 33367 6749 33376 6783
rect 33324 6740 33376 6749
rect 23112 6672 23164 6724
rect 20996 6604 21048 6656
rect 22284 6604 22336 6656
rect 23204 6604 23256 6656
rect 24676 6672 24728 6724
rect 26792 6604 26844 6656
rect 27068 6604 27120 6656
rect 28908 6647 28960 6656
rect 28908 6613 28917 6647
rect 28917 6613 28951 6647
rect 28951 6613 28960 6647
rect 28908 6604 28960 6613
rect 30564 6604 30616 6656
rect 31668 6604 31720 6656
rect 32588 6604 32640 6656
rect 33968 6740 34020 6792
rect 36176 6808 36228 6860
rect 36360 6808 36412 6860
rect 36452 6851 36504 6860
rect 36452 6817 36461 6851
rect 36461 6817 36495 6851
rect 36495 6817 36504 6851
rect 36452 6808 36504 6817
rect 37004 6808 37056 6860
rect 37648 6808 37700 6860
rect 35256 6783 35308 6792
rect 35256 6749 35265 6783
rect 35265 6749 35299 6783
rect 35299 6749 35308 6783
rect 35256 6740 35308 6749
rect 34704 6672 34756 6724
rect 37188 6783 37240 6792
rect 37188 6749 37197 6783
rect 37197 6749 37231 6783
rect 37231 6749 37240 6783
rect 37188 6740 37240 6749
rect 35992 6715 36044 6724
rect 35992 6681 36001 6715
rect 36001 6681 36035 6715
rect 36035 6681 36044 6715
rect 35992 6672 36044 6681
rect 38614 6808 38666 6860
rect 38936 6808 38988 6860
rect 41972 6808 42024 6860
rect 42432 6851 42484 6860
rect 42432 6817 42441 6851
rect 42441 6817 42475 6851
rect 42475 6817 42484 6851
rect 42432 6808 42484 6817
rect 42984 6808 43036 6860
rect 46204 6987 46256 6996
rect 46204 6953 46213 6987
rect 46213 6953 46247 6987
rect 46247 6953 46256 6987
rect 46204 6944 46256 6953
rect 46388 6944 46440 6996
rect 47308 6944 47360 6996
rect 49792 6944 49844 6996
rect 47860 6876 47912 6928
rect 41880 6783 41932 6792
rect 41880 6749 41889 6783
rect 41889 6749 41923 6783
rect 41923 6749 41932 6783
rect 41880 6740 41932 6749
rect 42156 6783 42208 6792
rect 42156 6749 42165 6783
rect 42165 6749 42199 6783
rect 42199 6749 42208 6783
rect 42156 6740 42208 6749
rect 43260 6808 43312 6860
rect 45560 6851 45612 6860
rect 45560 6817 45569 6851
rect 45569 6817 45603 6851
rect 45603 6817 45612 6851
rect 45560 6808 45612 6817
rect 48044 6808 48096 6860
rect 51448 6808 51500 6860
rect 54208 6987 54260 6996
rect 54208 6953 54217 6987
rect 54217 6953 54251 6987
rect 54251 6953 54260 6987
rect 54208 6944 54260 6953
rect 57060 6944 57112 6996
rect 52828 6808 52880 6860
rect 53932 6851 53984 6860
rect 53932 6817 53941 6851
rect 53941 6817 53975 6851
rect 53975 6817 53984 6851
rect 53932 6808 53984 6817
rect 54300 6808 54352 6860
rect 56324 6808 56376 6860
rect 57428 6851 57480 6860
rect 57428 6817 57437 6851
rect 57437 6817 57471 6851
rect 57471 6817 57480 6851
rect 57428 6808 57480 6817
rect 58440 6808 58492 6860
rect 38936 6715 38988 6724
rect 38936 6681 38945 6715
rect 38945 6681 38979 6715
rect 38979 6681 38988 6715
rect 38936 6672 38988 6681
rect 40132 6672 40184 6724
rect 41328 6672 41380 6724
rect 40040 6647 40092 6656
rect 40040 6613 40049 6647
rect 40049 6613 40083 6647
rect 40083 6613 40092 6647
rect 40040 6604 40092 6613
rect 40408 6647 40460 6656
rect 40408 6613 40417 6647
rect 40417 6613 40451 6647
rect 40451 6613 40460 6647
rect 40408 6604 40460 6613
rect 42524 6604 42576 6656
rect 42616 6604 42668 6656
rect 44640 6740 44692 6792
rect 46848 6740 46900 6792
rect 48412 6783 48464 6792
rect 48412 6749 48421 6783
rect 48421 6749 48455 6783
rect 48455 6749 48464 6783
rect 48412 6740 48464 6749
rect 43260 6672 43312 6724
rect 46296 6672 46348 6724
rect 46388 6715 46440 6724
rect 46388 6681 46397 6715
rect 46397 6681 46431 6715
rect 46431 6681 46440 6715
rect 46388 6672 46440 6681
rect 47400 6672 47452 6724
rect 51632 6783 51684 6792
rect 51632 6749 51641 6783
rect 51641 6749 51675 6783
rect 51675 6749 51684 6783
rect 51632 6740 51684 6749
rect 43168 6647 43220 6656
rect 43168 6613 43177 6647
rect 43177 6613 43211 6647
rect 43211 6613 43220 6647
rect 43168 6604 43220 6613
rect 47032 6604 47084 6656
rect 47952 6604 48004 6656
rect 52000 6604 52052 6656
rect 52184 6604 52236 6656
rect 52644 6740 52696 6792
rect 55128 6740 55180 6792
rect 56600 6740 56652 6792
rect 56876 6715 56928 6724
rect 56876 6681 56885 6715
rect 56885 6681 56919 6715
rect 56919 6681 56928 6715
rect 56876 6672 56928 6681
rect 57612 6715 57664 6724
rect 57612 6681 57621 6715
rect 57621 6681 57655 6715
rect 57655 6681 57664 6715
rect 57612 6672 57664 6681
rect 57704 6672 57756 6724
rect 53380 6647 53432 6656
rect 53380 6613 53389 6647
rect 53389 6613 53423 6647
rect 53423 6613 53432 6647
rect 53380 6604 53432 6613
rect 55588 6647 55640 6656
rect 55588 6613 55597 6647
rect 55597 6613 55631 6647
rect 55631 6613 55640 6647
rect 55588 6604 55640 6613
rect 57244 6604 57296 6656
rect 58256 6672 58308 6724
rect 15394 6502 15446 6554
rect 15458 6502 15510 6554
rect 15522 6502 15574 6554
rect 15586 6502 15638 6554
rect 15650 6502 15702 6554
rect 29838 6502 29890 6554
rect 29902 6502 29954 6554
rect 29966 6502 30018 6554
rect 30030 6502 30082 6554
rect 30094 6502 30146 6554
rect 44282 6502 44334 6554
rect 44346 6502 44398 6554
rect 44410 6502 44462 6554
rect 44474 6502 44526 6554
rect 44538 6502 44590 6554
rect 58726 6502 58778 6554
rect 58790 6502 58842 6554
rect 58854 6502 58906 6554
rect 58918 6502 58970 6554
rect 58982 6502 59034 6554
rect 3424 6400 3476 6452
rect 4252 6400 4304 6452
rect 4988 6400 5040 6452
rect 6000 6400 6052 6452
rect 8944 6400 8996 6452
rect 11980 6400 12032 6452
rect 12072 6443 12124 6452
rect 12072 6409 12081 6443
rect 12081 6409 12115 6443
rect 12115 6409 12124 6443
rect 12072 6400 12124 6409
rect 12992 6400 13044 6452
rect 13360 6400 13412 6452
rect 14280 6400 14332 6452
rect 16488 6400 16540 6452
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3516 6264 3568 6316
rect 3884 6196 3936 6248
rect 11704 6332 11756 6384
rect 5908 6264 5960 6316
rect 8852 6264 8904 6316
rect 9772 6264 9824 6316
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 12440 6264 12492 6316
rect 12900 6264 12952 6316
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 10968 6196 11020 6248
rect 5264 6171 5316 6180
rect 5264 6137 5273 6171
rect 5273 6137 5307 6171
rect 5307 6137 5316 6171
rect 5264 6128 5316 6137
rect 5448 6128 5500 6180
rect 5632 6171 5684 6180
rect 5632 6137 5641 6171
rect 5641 6137 5675 6171
rect 5675 6137 5684 6171
rect 5632 6128 5684 6137
rect 5908 6128 5960 6180
rect 12348 6128 12400 6180
rect 16028 6332 16080 6384
rect 17776 6400 17828 6452
rect 17868 6400 17920 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 23112 6400 23164 6452
rect 23388 6400 23440 6452
rect 26332 6400 26384 6452
rect 27988 6443 28040 6452
rect 27988 6409 27997 6443
rect 27997 6409 28031 6443
rect 28031 6409 28040 6443
rect 27988 6400 28040 6409
rect 28632 6400 28684 6452
rect 30656 6400 30708 6452
rect 18328 6332 18380 6384
rect 15200 6307 15252 6316
rect 15200 6273 15234 6307
rect 15234 6273 15252 6307
rect 15200 6264 15252 6273
rect 17408 6264 17460 6316
rect 17592 6264 17644 6316
rect 18512 6264 18564 6316
rect 19064 6307 19116 6316
rect 19064 6273 19073 6307
rect 19073 6273 19107 6307
rect 19107 6273 19116 6307
rect 19064 6264 19116 6273
rect 19616 6264 19668 6316
rect 21732 6264 21784 6316
rect 22100 6375 22152 6384
rect 22100 6341 22134 6375
rect 22134 6341 22152 6375
rect 22100 6332 22152 6341
rect 29092 6332 29144 6384
rect 34888 6400 34940 6452
rect 36176 6400 36228 6452
rect 31852 6332 31904 6384
rect 32220 6332 32272 6384
rect 37832 6400 37884 6452
rect 38476 6400 38528 6452
rect 14188 6196 14240 6248
rect 14372 6196 14424 6248
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 4068 6060 4120 6112
rect 4344 6060 4396 6112
rect 18880 6196 18932 6248
rect 21180 6239 21232 6248
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6184 6060 6236 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 14004 6060 14056 6112
rect 14740 6060 14792 6112
rect 20720 6128 20772 6180
rect 17040 6060 17092 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 23296 6264 23348 6316
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 26516 6307 26568 6316
rect 26516 6273 26525 6307
rect 26525 6273 26559 6307
rect 26559 6273 26568 6307
rect 26516 6264 26568 6273
rect 27528 6264 27580 6316
rect 30472 6264 30524 6316
rect 31208 6264 31260 6316
rect 32312 6264 32364 6316
rect 32496 6264 32548 6316
rect 34612 6264 34664 6316
rect 36728 6264 36780 6316
rect 37188 6264 37240 6316
rect 38108 6264 38160 6316
rect 38844 6307 38896 6316
rect 38844 6273 38853 6307
rect 38853 6273 38887 6307
rect 38887 6273 38896 6307
rect 38844 6264 38896 6273
rect 39672 6307 39724 6316
rect 39672 6273 39706 6307
rect 39706 6273 39724 6307
rect 39672 6264 39724 6273
rect 39948 6264 40000 6316
rect 40408 6400 40460 6452
rect 41972 6400 42024 6452
rect 47400 6443 47452 6452
rect 47400 6409 47409 6443
rect 47409 6409 47443 6443
rect 47443 6409 47452 6443
rect 47400 6400 47452 6409
rect 48412 6400 48464 6452
rect 40132 6332 40184 6384
rect 42432 6332 42484 6384
rect 23204 6196 23256 6248
rect 24676 6196 24728 6248
rect 31760 6239 31812 6248
rect 31760 6205 31769 6239
rect 31769 6205 31803 6239
rect 31803 6205 31812 6239
rect 31760 6196 31812 6205
rect 22192 6060 22244 6112
rect 23296 6103 23348 6112
rect 23296 6069 23305 6103
rect 23305 6069 23339 6103
rect 23339 6069 23348 6103
rect 23296 6060 23348 6069
rect 34520 6128 34572 6180
rect 33876 6103 33928 6112
rect 33876 6069 33885 6103
rect 33885 6069 33919 6103
rect 33919 6069 33928 6103
rect 33876 6060 33928 6069
rect 37464 6060 37516 6112
rect 38292 6103 38344 6112
rect 38292 6069 38301 6103
rect 38301 6069 38335 6103
rect 38335 6069 38344 6103
rect 38292 6060 38344 6069
rect 41788 6264 41840 6316
rect 44548 6332 44600 6384
rect 42616 6196 42668 6248
rect 41052 6128 41104 6180
rect 41420 6128 41472 6180
rect 45928 6264 45980 6316
rect 46848 6264 46900 6316
rect 47308 6264 47360 6316
rect 48044 6307 48096 6316
rect 48044 6273 48053 6307
rect 48053 6273 48087 6307
rect 48087 6273 48096 6307
rect 48044 6264 48096 6273
rect 47400 6196 47452 6248
rect 50896 6332 50948 6384
rect 49332 6307 49384 6316
rect 49332 6273 49366 6307
rect 49366 6273 49384 6307
rect 49332 6264 49384 6273
rect 50160 6264 50212 6316
rect 52644 6400 52696 6452
rect 55404 6400 55456 6452
rect 56968 6400 57020 6452
rect 52276 6375 52328 6384
rect 52276 6341 52285 6375
rect 52285 6341 52319 6375
rect 52319 6341 52328 6375
rect 52276 6332 52328 6341
rect 52000 6264 52052 6316
rect 58256 6400 58308 6452
rect 54116 6196 54168 6248
rect 55496 6239 55548 6248
rect 55496 6205 55505 6239
rect 55505 6205 55539 6239
rect 55539 6205 55548 6239
rect 55496 6196 55548 6205
rect 43260 6103 43312 6112
rect 43260 6069 43269 6103
rect 43269 6069 43303 6103
rect 43303 6069 43312 6103
rect 43260 6060 43312 6069
rect 50436 6103 50488 6112
rect 50436 6069 50445 6103
rect 50445 6069 50479 6103
rect 50479 6069 50488 6103
rect 50436 6060 50488 6069
rect 50804 6060 50856 6112
rect 54852 6060 54904 6112
rect 54944 6103 54996 6112
rect 54944 6069 54953 6103
rect 54953 6069 54987 6103
rect 54987 6069 54996 6103
rect 54944 6060 54996 6069
rect 55404 6103 55456 6112
rect 55404 6069 55413 6103
rect 55413 6069 55447 6103
rect 55447 6069 55456 6103
rect 55404 6060 55456 6069
rect 56140 6103 56192 6112
rect 56140 6069 56149 6103
rect 56149 6069 56183 6103
rect 56183 6069 56192 6103
rect 56140 6060 56192 6069
rect 57060 6103 57112 6112
rect 57060 6069 57069 6103
rect 57069 6069 57103 6103
rect 57103 6069 57112 6103
rect 57060 6060 57112 6069
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 22616 5958 22668 6010
rect 22680 5958 22732 6010
rect 22744 5958 22796 6010
rect 22808 5958 22860 6010
rect 22872 5958 22924 6010
rect 37060 5958 37112 6010
rect 37124 5958 37176 6010
rect 37188 5958 37240 6010
rect 37252 5958 37304 6010
rect 37316 5958 37368 6010
rect 51504 5958 51556 6010
rect 51568 5958 51620 6010
rect 51632 5958 51684 6010
rect 51696 5958 51748 6010
rect 51760 5958 51812 6010
rect 1860 5856 1912 5908
rect 2964 5899 3016 5908
rect 1952 5788 2004 5840
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 3240 5788 3292 5840
rect 3148 5720 3200 5772
rect 5908 5856 5960 5908
rect 6092 5856 6144 5908
rect 7656 5856 7708 5908
rect 8760 5856 8812 5908
rect 12440 5856 12492 5908
rect 13544 5856 13596 5908
rect 15292 5856 15344 5908
rect 16120 5856 16172 5908
rect 17040 5856 17092 5908
rect 17684 5856 17736 5908
rect 19616 5856 19668 5908
rect 20536 5856 20588 5908
rect 20720 5856 20772 5908
rect 21732 5856 21784 5908
rect 28908 5856 28960 5908
rect 30564 5856 30616 5908
rect 31208 5899 31260 5908
rect 31208 5865 31217 5899
rect 31217 5865 31251 5899
rect 31251 5865 31260 5899
rect 31208 5856 31260 5865
rect 32588 5856 32640 5908
rect 35256 5856 35308 5908
rect 37464 5856 37516 5908
rect 38108 5899 38160 5908
rect 38108 5865 38117 5899
rect 38117 5865 38151 5899
rect 38151 5865 38160 5899
rect 38108 5856 38160 5865
rect 39304 5856 39356 5908
rect 39672 5856 39724 5908
rect 40132 5856 40184 5908
rect 42616 5856 42668 5908
rect 44548 5856 44600 5908
rect 47400 5899 47452 5908
rect 47400 5865 47409 5899
rect 47409 5865 47443 5899
rect 47443 5865 47452 5899
rect 47400 5856 47452 5865
rect 49332 5899 49384 5908
rect 49332 5865 49341 5899
rect 49341 5865 49375 5899
rect 49375 5865 49384 5899
rect 49332 5856 49384 5865
rect 9128 5720 9180 5772
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 14188 5763 14240 5772
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4344 5695 4396 5704
rect 4344 5661 4378 5695
rect 4378 5661 4396 5695
rect 4344 5652 4396 5661
rect 5448 5652 5500 5704
rect 5540 5652 5592 5704
rect 6184 5652 6236 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 12532 5652 12584 5704
rect 7196 5584 7248 5636
rect 9956 5584 10008 5636
rect 10140 5627 10192 5636
rect 10140 5593 10174 5627
rect 10174 5593 10192 5627
rect 10140 5584 10192 5593
rect 13912 5652 13964 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 14096 5584 14148 5636
rect 4528 5516 4580 5568
rect 5264 5516 5316 5568
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 14004 5516 14056 5568
rect 15936 5584 15988 5636
rect 17960 5652 18012 5704
rect 23480 5720 23532 5772
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 26608 5720 26660 5772
rect 26884 5720 26936 5772
rect 28632 5720 28684 5772
rect 31116 5788 31168 5840
rect 33232 5720 33284 5772
rect 33324 5720 33376 5772
rect 33784 5763 33836 5772
rect 33784 5729 33793 5763
rect 33793 5729 33827 5763
rect 33827 5729 33836 5763
rect 33784 5720 33836 5729
rect 35072 5788 35124 5840
rect 34704 5720 34756 5772
rect 34888 5720 34940 5772
rect 27160 5652 27212 5704
rect 15844 5516 15896 5568
rect 17684 5559 17736 5568
rect 17684 5525 17693 5559
rect 17693 5525 17727 5559
rect 17727 5525 17736 5559
rect 17684 5516 17736 5525
rect 19340 5516 19392 5568
rect 20352 5516 20404 5568
rect 25596 5584 25648 5636
rect 28816 5695 28868 5704
rect 28816 5661 28825 5695
rect 28825 5661 28859 5695
rect 28859 5661 28868 5695
rect 28816 5652 28868 5661
rect 33140 5652 33192 5704
rect 30656 5584 30708 5636
rect 33968 5652 34020 5704
rect 37648 5788 37700 5840
rect 41696 5788 41748 5840
rect 36820 5584 36872 5636
rect 41512 5720 41564 5772
rect 46296 5788 46348 5840
rect 49700 5788 49752 5840
rect 51264 5856 51316 5908
rect 55128 5899 55180 5908
rect 55128 5865 55137 5899
rect 55137 5865 55171 5899
rect 55171 5865 55180 5899
rect 55128 5856 55180 5865
rect 38660 5652 38712 5704
rect 40040 5652 40092 5704
rect 50620 5763 50672 5772
rect 43260 5652 43312 5704
rect 22192 5516 22244 5568
rect 26240 5516 26292 5568
rect 28264 5559 28316 5568
rect 28264 5525 28273 5559
rect 28273 5525 28307 5559
rect 28307 5525 28316 5559
rect 28264 5516 28316 5525
rect 29552 5559 29604 5568
rect 29552 5525 29561 5559
rect 29561 5525 29595 5559
rect 29595 5525 29604 5559
rect 29552 5516 29604 5525
rect 33324 5559 33376 5568
rect 33324 5525 33333 5559
rect 33333 5525 33367 5559
rect 33367 5525 33376 5559
rect 33324 5516 33376 5525
rect 33416 5516 33468 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 39120 5559 39172 5568
rect 39120 5525 39129 5559
rect 39129 5525 39163 5559
rect 39163 5525 39172 5559
rect 39120 5516 39172 5525
rect 41696 5559 41748 5568
rect 41696 5525 41705 5559
rect 41705 5525 41739 5559
rect 41739 5525 41748 5559
rect 41696 5516 41748 5525
rect 42708 5516 42760 5568
rect 42984 5516 43036 5568
rect 45468 5652 45520 5704
rect 46112 5695 46164 5704
rect 46112 5661 46121 5695
rect 46121 5661 46155 5695
rect 46155 5661 46164 5695
rect 46112 5652 46164 5661
rect 46204 5652 46256 5704
rect 44180 5584 44232 5636
rect 50620 5729 50629 5763
rect 50629 5729 50663 5763
rect 50663 5729 50672 5763
rect 50620 5720 50672 5729
rect 50804 5788 50856 5840
rect 52184 5788 52236 5840
rect 58348 5831 58400 5840
rect 58348 5797 58357 5831
rect 58357 5797 58391 5831
rect 58391 5797 58400 5831
rect 58348 5788 58400 5797
rect 51632 5763 51684 5772
rect 51632 5729 51641 5763
rect 51641 5729 51675 5763
rect 51675 5729 51684 5763
rect 51632 5720 51684 5729
rect 52000 5720 52052 5772
rect 51356 5652 51408 5704
rect 52736 5652 52788 5704
rect 56324 5652 56376 5704
rect 57060 5695 57112 5704
rect 57060 5661 57094 5695
rect 57094 5661 57112 5695
rect 57060 5652 57112 5661
rect 58532 5695 58584 5704
rect 58532 5661 58541 5695
rect 58541 5661 58575 5695
rect 58575 5661 58584 5695
rect 58532 5652 58584 5661
rect 44640 5559 44692 5568
rect 44640 5525 44649 5559
rect 44649 5525 44683 5559
rect 44683 5525 44692 5559
rect 44640 5516 44692 5525
rect 45560 5559 45612 5568
rect 45560 5525 45569 5559
rect 45569 5525 45603 5559
rect 45603 5525 45612 5559
rect 45560 5516 45612 5525
rect 46296 5516 46348 5568
rect 56140 5584 56192 5636
rect 52000 5516 52052 5568
rect 52644 5559 52696 5568
rect 52644 5525 52653 5559
rect 52653 5525 52687 5559
rect 52687 5525 52696 5559
rect 52644 5516 52696 5525
rect 52828 5516 52880 5568
rect 54668 5516 54720 5568
rect 56692 5559 56744 5568
rect 56692 5525 56701 5559
rect 56701 5525 56735 5559
rect 56735 5525 56744 5559
rect 56692 5516 56744 5525
rect 57244 5516 57296 5568
rect 15394 5414 15446 5466
rect 15458 5414 15510 5466
rect 15522 5414 15574 5466
rect 15586 5414 15638 5466
rect 15650 5414 15702 5466
rect 29838 5414 29890 5466
rect 29902 5414 29954 5466
rect 29966 5414 30018 5466
rect 30030 5414 30082 5466
rect 30094 5414 30146 5466
rect 44282 5414 44334 5466
rect 44346 5414 44398 5466
rect 44410 5414 44462 5466
rect 44474 5414 44526 5466
rect 44538 5414 44590 5466
rect 58726 5414 58778 5466
rect 58790 5414 58842 5466
rect 58854 5414 58906 5466
rect 58918 5414 58970 5466
rect 58982 5414 59034 5466
rect 3240 5312 3292 5364
rect 2964 5287 3016 5296
rect 2964 5253 2973 5287
rect 2973 5253 3007 5287
rect 3007 5253 3016 5287
rect 2964 5244 3016 5253
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 4436 5312 4488 5364
rect 5632 5312 5684 5364
rect 12256 5312 12308 5364
rect 3792 5287 3844 5296
rect 3792 5253 3801 5287
rect 3801 5253 3835 5287
rect 3835 5253 3844 5287
rect 3792 5244 3844 5253
rect 3516 5176 3568 5228
rect 5540 5244 5592 5296
rect 7656 5287 7708 5296
rect 7656 5253 7665 5287
rect 7665 5253 7699 5287
rect 7699 5253 7708 5287
rect 7656 5244 7708 5253
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 7288 5176 7340 5228
rect 9128 5176 9180 5228
rect 11152 5244 11204 5296
rect 22008 5312 22060 5364
rect 22836 5312 22888 5364
rect 23296 5312 23348 5364
rect 25596 5355 25648 5364
rect 25596 5321 25605 5355
rect 25605 5321 25639 5355
rect 25639 5321 25648 5355
rect 25596 5312 25648 5321
rect 26608 5355 26660 5364
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 32496 5355 32548 5364
rect 32496 5321 32505 5355
rect 32505 5321 32539 5355
rect 32539 5321 32548 5355
rect 32496 5312 32548 5321
rect 33140 5312 33192 5364
rect 33784 5312 33836 5364
rect 34704 5312 34756 5364
rect 36820 5312 36872 5364
rect 37556 5312 37608 5364
rect 9864 5176 9916 5228
rect 10048 5176 10100 5228
rect 11244 5176 11296 5228
rect 1860 5040 1912 5092
rect 3424 5040 3476 5092
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 3240 4972 3292 5024
rect 3976 5040 4028 5092
rect 5264 5040 5316 5092
rect 5356 5083 5408 5092
rect 5356 5049 5365 5083
rect 5365 5049 5399 5083
rect 5399 5049 5408 5083
rect 5356 5040 5408 5049
rect 5816 4972 5868 5024
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 9220 5083 9272 5092
rect 9220 5049 9229 5083
rect 9229 5049 9263 5083
rect 9263 5049 9272 5083
rect 9220 5040 9272 5049
rect 14740 5244 14792 5296
rect 15200 5244 15252 5296
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 15936 5244 15988 5296
rect 17684 5287 17736 5296
rect 17684 5253 17718 5287
rect 17718 5253 17736 5287
rect 17684 5244 17736 5253
rect 18420 5244 18472 5296
rect 18972 5244 19024 5296
rect 15844 5176 15896 5228
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 19340 5176 19392 5228
rect 21180 5176 21232 5228
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 16120 5040 16172 5092
rect 28264 5244 28316 5296
rect 35900 5244 35952 5296
rect 36728 5287 36780 5296
rect 36728 5253 36737 5287
rect 36737 5253 36771 5287
rect 36771 5253 36780 5287
rect 36728 5244 36780 5253
rect 41696 5244 41748 5296
rect 43168 5312 43220 5364
rect 45560 5312 45612 5364
rect 46112 5312 46164 5364
rect 43076 5244 43128 5296
rect 23388 5176 23440 5228
rect 25872 5176 25924 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 33324 5176 33376 5228
rect 33508 5176 33560 5228
rect 34520 5219 34572 5228
rect 34520 5185 34529 5219
rect 34529 5185 34563 5219
rect 34563 5185 34572 5219
rect 34520 5176 34572 5185
rect 34704 5219 34756 5228
rect 34704 5185 34713 5219
rect 34713 5185 34747 5219
rect 34747 5185 34756 5219
rect 34704 5176 34756 5185
rect 34888 5219 34940 5228
rect 34888 5185 34897 5219
rect 34897 5185 34931 5219
rect 34931 5185 34940 5219
rect 34888 5176 34940 5185
rect 37464 5176 37516 5228
rect 38200 5176 38252 5228
rect 39120 5176 39172 5228
rect 25320 5108 25372 5160
rect 39948 5108 40000 5160
rect 40868 5108 40920 5160
rect 41512 5108 41564 5160
rect 14924 4972 14976 5024
rect 17592 4972 17644 5024
rect 18144 4972 18196 5024
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 20996 5015 21048 5024
rect 19892 4972 19944 4981
rect 20996 4981 21005 5015
rect 21005 4981 21039 5015
rect 21039 4981 21048 5015
rect 20996 4972 21048 4981
rect 21732 4972 21784 5024
rect 23296 4972 23348 5024
rect 24032 4972 24084 5024
rect 30288 4972 30340 5024
rect 30656 4972 30708 5024
rect 36176 5040 36228 5092
rect 44180 5244 44232 5296
rect 47032 5312 47084 5364
rect 49700 5312 49752 5364
rect 51356 5312 51408 5364
rect 51632 5312 51684 5364
rect 45928 5176 45980 5228
rect 46480 5176 46532 5228
rect 52000 5244 52052 5296
rect 52368 5244 52420 5296
rect 52736 5355 52788 5364
rect 52736 5321 52745 5355
rect 52745 5321 52779 5355
rect 52779 5321 52788 5355
rect 52736 5312 52788 5321
rect 53380 5312 53432 5364
rect 55496 5312 55548 5364
rect 55588 5312 55640 5364
rect 57704 5355 57756 5364
rect 57704 5321 57713 5355
rect 57713 5321 57747 5355
rect 57747 5321 57756 5355
rect 57704 5312 57756 5321
rect 32404 5015 32456 5024
rect 32404 4981 32413 5015
rect 32413 4981 32447 5015
rect 32447 4981 32456 5015
rect 32404 4972 32456 4981
rect 34060 4972 34112 5024
rect 34796 4972 34848 5024
rect 38752 5015 38804 5024
rect 38752 4981 38761 5015
rect 38761 4981 38795 5015
rect 38795 4981 38804 5015
rect 38752 4972 38804 4981
rect 38844 4972 38896 5024
rect 40684 4972 40736 5024
rect 41512 4972 41564 5024
rect 41604 5015 41656 5024
rect 41604 4981 41613 5015
rect 41613 4981 41647 5015
rect 41647 4981 41656 5015
rect 41604 4972 41656 4981
rect 42248 4972 42300 5024
rect 45652 5108 45704 5160
rect 46296 5151 46348 5160
rect 46296 5117 46305 5151
rect 46305 5117 46339 5151
rect 46339 5117 46348 5151
rect 46296 5108 46348 5117
rect 47860 5108 47912 5160
rect 50436 5176 50488 5228
rect 51264 5176 51316 5228
rect 53564 5176 53616 5228
rect 53932 5176 53984 5228
rect 55128 5176 55180 5228
rect 55404 5176 55456 5228
rect 56324 5219 56376 5228
rect 56324 5185 56333 5219
rect 56333 5185 56367 5219
rect 56367 5185 56376 5219
rect 56324 5176 56376 5185
rect 56416 5176 56468 5228
rect 58440 5219 58492 5228
rect 58440 5185 58449 5219
rect 58449 5185 58483 5219
rect 58483 5185 58492 5219
rect 58440 5176 58492 5185
rect 43076 4972 43128 5024
rect 50252 5040 50304 5092
rect 46848 4972 46900 5024
rect 49332 4972 49384 5024
rect 49700 5015 49752 5024
rect 49700 4981 49709 5015
rect 49709 4981 49743 5015
rect 49743 4981 49752 5015
rect 49700 4972 49752 4981
rect 50988 4972 51040 5024
rect 51356 4972 51408 5024
rect 54668 4972 54720 5024
rect 54852 5015 54904 5024
rect 54852 4981 54861 5015
rect 54861 4981 54895 5015
rect 54895 4981 54904 5015
rect 54852 4972 54904 4981
rect 56324 5040 56376 5092
rect 56968 4972 57020 5024
rect 57888 5015 57940 5024
rect 57888 4981 57897 5015
rect 57897 4981 57931 5015
rect 57931 4981 57940 5015
rect 57888 4972 57940 4981
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 22616 4870 22668 4922
rect 22680 4870 22732 4922
rect 22744 4870 22796 4922
rect 22808 4870 22860 4922
rect 22872 4870 22924 4922
rect 37060 4870 37112 4922
rect 37124 4870 37176 4922
rect 37188 4870 37240 4922
rect 37252 4870 37304 4922
rect 37316 4870 37368 4922
rect 51504 4870 51556 4922
rect 51568 4870 51620 4922
rect 51632 4870 51684 4922
rect 51696 4870 51748 4922
rect 51760 4870 51812 4922
rect 2780 4768 2832 4820
rect 3240 4768 3292 4820
rect 7748 4768 7800 4820
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 4436 4675 4488 4684
rect 4436 4641 4445 4675
rect 4445 4641 4479 4675
rect 4479 4641 4488 4675
rect 4436 4632 4488 4641
rect 3424 4564 3476 4616
rect 4896 4607 4948 4616
rect 4896 4573 4913 4607
rect 4913 4573 4947 4607
rect 4947 4573 4948 4607
rect 4896 4564 4948 4573
rect 5264 4564 5316 4616
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 7012 4700 7064 4752
rect 10968 4700 11020 4752
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 11704 4768 11756 4820
rect 13452 4768 13504 4820
rect 15200 4768 15252 4820
rect 16488 4768 16540 4820
rect 16580 4768 16632 4820
rect 16764 4743 16816 4752
rect 16764 4709 16773 4743
rect 16773 4709 16807 4743
rect 16807 4709 16816 4743
rect 16764 4700 16816 4709
rect 17960 4768 18012 4820
rect 18328 4768 18380 4820
rect 20996 4768 21048 4820
rect 21456 4768 21508 4820
rect 24768 4768 24820 4820
rect 25044 4768 25096 4820
rect 25320 4768 25372 4820
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 1952 4428 2004 4480
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 5724 4496 5776 4548
rect 4988 4428 5040 4480
rect 5264 4428 5316 4480
rect 7380 4564 7432 4616
rect 8116 4564 8168 4616
rect 8392 4564 8444 4616
rect 10508 4564 10560 4616
rect 16580 4632 16632 4684
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18144 4632 18196 4641
rect 18420 4632 18472 4684
rect 9128 4496 9180 4548
rect 13728 4564 13780 4616
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 10968 4496 11020 4548
rect 14004 4496 14056 4548
rect 14096 4539 14148 4548
rect 14096 4505 14105 4539
rect 14105 4505 14139 4539
rect 14139 4505 14148 4539
rect 14096 4496 14148 4505
rect 14188 4496 14240 4548
rect 18236 4496 18288 4548
rect 18328 4496 18380 4548
rect 19340 4564 19392 4616
rect 19524 4607 19576 4616
rect 19524 4573 19533 4607
rect 19533 4573 19567 4607
rect 19567 4573 19576 4607
rect 19524 4564 19576 4573
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 24952 4632 25004 4684
rect 25044 4632 25096 4684
rect 27528 4632 27580 4684
rect 25228 4564 25280 4616
rect 25320 4607 25372 4616
rect 25320 4573 25329 4607
rect 25329 4573 25363 4607
rect 25363 4573 25372 4607
rect 25320 4564 25372 4573
rect 20076 4496 20128 4548
rect 20444 4496 20496 4548
rect 21732 4496 21784 4548
rect 24032 4496 24084 4548
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 7840 4428 7892 4480
rect 8300 4428 8352 4480
rect 10508 4471 10560 4480
rect 10508 4437 10517 4471
rect 10517 4437 10551 4471
rect 10551 4437 10560 4471
rect 10508 4428 10560 4437
rect 12440 4428 12492 4480
rect 14280 4428 14332 4480
rect 14924 4428 14976 4480
rect 15108 4428 15160 4480
rect 16120 4428 16172 4480
rect 18604 4471 18656 4480
rect 18604 4437 18613 4471
rect 18613 4437 18647 4471
rect 18647 4437 18656 4471
rect 18604 4428 18656 4437
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 20628 4428 20680 4480
rect 22284 4428 22336 4480
rect 23296 4428 23348 4480
rect 24216 4428 24268 4480
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 26240 4428 26292 4480
rect 27620 4428 27672 4480
rect 28816 4768 28868 4820
rect 28908 4768 28960 4820
rect 31392 4768 31444 4820
rect 28172 4700 28224 4752
rect 34152 4768 34204 4820
rect 34888 4768 34940 4820
rect 28172 4564 28224 4616
rect 29552 4564 29604 4616
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 32404 4632 32456 4684
rect 37556 4768 37608 4820
rect 38660 4768 38712 4820
rect 42616 4768 42668 4820
rect 42708 4768 42760 4820
rect 39120 4700 39172 4752
rect 30288 4496 30340 4548
rect 31392 4496 31444 4548
rect 33876 4564 33928 4616
rect 34060 4564 34112 4616
rect 34980 4564 35032 4616
rect 34152 4496 34204 4548
rect 28356 4428 28408 4480
rect 29184 4428 29236 4480
rect 29644 4428 29696 4480
rect 31116 4471 31168 4480
rect 31116 4437 31125 4471
rect 31125 4437 31159 4471
rect 31159 4437 31168 4471
rect 31116 4428 31168 4437
rect 32128 4428 32180 4480
rect 33508 4428 33560 4480
rect 33876 4471 33928 4480
rect 33876 4437 33885 4471
rect 33885 4437 33919 4471
rect 33919 4437 33928 4471
rect 33876 4428 33928 4437
rect 35900 4607 35952 4616
rect 38752 4675 38804 4684
rect 38752 4641 38761 4675
rect 38761 4641 38795 4675
rect 38795 4641 38804 4675
rect 38752 4632 38804 4641
rect 38844 4632 38896 4684
rect 39396 4632 39448 4684
rect 35900 4573 35914 4607
rect 35914 4573 35948 4607
rect 35948 4573 35952 4607
rect 35900 4564 35952 4573
rect 38292 4564 38344 4616
rect 36268 4496 36320 4548
rect 36452 4496 36504 4548
rect 39672 4564 39724 4616
rect 37648 4428 37700 4480
rect 40132 4496 40184 4548
rect 40868 4675 40920 4684
rect 40868 4641 40877 4675
rect 40877 4641 40911 4675
rect 40911 4641 40920 4675
rect 40868 4632 40920 4641
rect 45744 4700 45796 4752
rect 46480 4700 46532 4752
rect 41604 4564 41656 4616
rect 43076 4607 43128 4616
rect 43076 4573 43085 4607
rect 43085 4573 43119 4607
rect 43119 4573 43128 4607
rect 43076 4564 43128 4573
rect 44640 4632 44692 4684
rect 45928 4632 45980 4684
rect 49332 4768 49384 4820
rect 51356 4768 51408 4820
rect 51816 4768 51868 4820
rect 53840 4768 53892 4820
rect 54668 4811 54720 4820
rect 54668 4777 54677 4811
rect 54677 4777 54711 4811
rect 54711 4777 54720 4811
rect 54668 4768 54720 4777
rect 56416 4768 56468 4820
rect 57888 4768 57940 4820
rect 50160 4700 50212 4752
rect 42616 4496 42668 4548
rect 43812 4607 43864 4616
rect 43812 4573 43821 4607
rect 43821 4573 43855 4607
rect 43855 4573 43864 4607
rect 43812 4564 43864 4573
rect 44732 4607 44784 4616
rect 44732 4573 44741 4607
rect 44741 4573 44775 4607
rect 44775 4573 44784 4607
rect 44732 4564 44784 4573
rect 42248 4428 42300 4480
rect 43536 4428 43588 4480
rect 43628 4471 43680 4480
rect 43628 4437 43637 4471
rect 43637 4437 43671 4471
rect 43671 4437 43680 4471
rect 43628 4428 43680 4437
rect 43720 4428 43772 4480
rect 45284 4564 45336 4616
rect 46204 4564 46256 4616
rect 46848 4607 46900 4616
rect 46848 4573 46882 4607
rect 46882 4573 46900 4607
rect 46848 4564 46900 4573
rect 47768 4564 47820 4616
rect 49884 4607 49936 4616
rect 49884 4573 49893 4607
rect 49893 4573 49927 4607
rect 49927 4573 49936 4607
rect 49884 4564 49936 4573
rect 50160 4607 50212 4616
rect 50160 4573 50169 4607
rect 50169 4573 50203 4607
rect 50203 4573 50212 4607
rect 50160 4564 50212 4573
rect 53656 4700 53708 4752
rect 51816 4496 51868 4548
rect 45100 4428 45152 4480
rect 45468 4428 45520 4480
rect 46664 4428 46716 4480
rect 47124 4428 47176 4480
rect 47860 4428 47912 4480
rect 47952 4471 48004 4480
rect 47952 4437 47961 4471
rect 47961 4437 47995 4471
rect 47995 4437 48004 4471
rect 47952 4428 48004 4437
rect 48688 4471 48740 4480
rect 48688 4437 48697 4471
rect 48697 4437 48731 4471
rect 48731 4437 48740 4471
rect 48688 4428 48740 4437
rect 49700 4428 49752 4480
rect 50068 4428 50120 4480
rect 53012 4564 53064 4616
rect 53748 4607 53800 4616
rect 53748 4573 53757 4607
rect 53757 4573 53791 4607
rect 53791 4573 53800 4607
rect 53748 4564 53800 4573
rect 54852 4564 54904 4616
rect 56324 4675 56376 4684
rect 56324 4641 56333 4675
rect 56333 4641 56367 4675
rect 56367 4641 56376 4675
rect 56324 4632 56376 4641
rect 56692 4632 56744 4684
rect 52644 4496 52696 4548
rect 57152 4607 57204 4616
rect 57152 4573 57161 4607
rect 57161 4573 57195 4607
rect 57195 4573 57204 4607
rect 57152 4564 57204 4573
rect 57796 4496 57848 4548
rect 58624 4496 58676 4548
rect 53196 4428 53248 4480
rect 54116 4428 54168 4480
rect 54300 4471 54352 4480
rect 54300 4437 54309 4471
rect 54309 4437 54343 4471
rect 54343 4437 54352 4471
rect 54300 4428 54352 4437
rect 55220 4428 55272 4480
rect 15394 4326 15446 4378
rect 15458 4326 15510 4378
rect 15522 4326 15574 4378
rect 15586 4326 15638 4378
rect 15650 4326 15702 4378
rect 29838 4326 29890 4378
rect 29902 4326 29954 4378
rect 29966 4326 30018 4378
rect 30030 4326 30082 4378
rect 30094 4326 30146 4378
rect 44282 4326 44334 4378
rect 44346 4326 44398 4378
rect 44410 4326 44462 4378
rect 44474 4326 44526 4378
rect 44538 4326 44590 4378
rect 58726 4326 58778 4378
rect 58790 4326 58842 4378
rect 58854 4326 58906 4378
rect 58918 4326 58970 4378
rect 58982 4326 59034 4378
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2228 4088 2280 4140
rect 6000 4224 6052 4276
rect 2780 4156 2832 4208
rect 2872 4156 2924 4208
rect 3516 4088 3568 4140
rect 3976 4088 4028 4140
rect 4436 4156 4488 4208
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 2044 3884 2096 3936
rect 2228 3884 2280 3936
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 5356 4088 5408 4140
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 6460 4156 6512 4208
rect 5632 4088 5684 4140
rect 6184 4088 6236 4140
rect 7196 4088 7248 4140
rect 7840 4156 7892 4208
rect 9772 4156 9824 4208
rect 10508 4156 10560 4208
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 12440 4224 12492 4276
rect 4988 4020 5040 4029
rect 5724 4020 5776 4072
rect 6276 4020 6328 4072
rect 3792 3952 3844 3961
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 8116 3952 8168 4004
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8760 4088 8812 4140
rect 9220 4088 9272 4140
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 8668 3952 8720 4004
rect 9864 4020 9916 4072
rect 11060 4020 11112 4072
rect 3056 3884 3108 3936
rect 3332 3884 3384 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 7840 3884 7892 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 10600 3884 10652 3936
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 13544 4199 13596 4208
rect 13544 4165 13553 4199
rect 13553 4165 13587 4199
rect 13587 4165 13596 4199
rect 13544 4156 13596 4165
rect 13452 4131 13504 4140
rect 13452 4097 13456 4131
rect 13456 4097 13490 4131
rect 13490 4097 13504 4131
rect 14648 4224 14700 4276
rect 14740 4224 14792 4276
rect 13452 4088 13504 4097
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 14280 4156 14332 4208
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 15200 4156 15252 4208
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 20904 4224 20956 4276
rect 16396 4156 16448 4208
rect 16120 4088 16172 4140
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 17868 4199 17920 4208
rect 17868 4165 17877 4199
rect 17877 4165 17911 4199
rect 17911 4165 17920 4199
rect 17868 4156 17920 4165
rect 18144 4199 18196 4208
rect 18144 4165 18153 4199
rect 18153 4165 18187 4199
rect 18187 4165 18196 4199
rect 18144 4156 18196 4165
rect 18880 4156 18932 4208
rect 16028 4020 16080 4072
rect 16304 4063 16356 4072
rect 16304 4029 16313 4063
rect 16313 4029 16347 4063
rect 16347 4029 16356 4063
rect 16304 4020 16356 4029
rect 16396 4020 16448 4072
rect 18052 4020 18104 4072
rect 13360 3952 13412 4004
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14740 3952 14792 4004
rect 18236 3952 18288 4004
rect 15936 3884 15988 3936
rect 17316 3884 17368 3936
rect 18512 4131 18564 4140
rect 18512 4097 18526 4131
rect 18526 4097 18560 4131
rect 18560 4097 18564 4131
rect 18512 4088 18564 4097
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 19432 4088 19484 4140
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20076 4131 20128 4140
rect 21732 4156 21784 4208
rect 20076 4097 20090 4131
rect 20090 4097 20124 4131
rect 20124 4097 20128 4131
rect 20076 4088 20128 4097
rect 22284 4156 22336 4208
rect 23388 4267 23440 4276
rect 23388 4233 23397 4267
rect 23397 4233 23431 4267
rect 23431 4233 23440 4267
rect 23388 4224 23440 4233
rect 27896 4224 27948 4276
rect 24216 4156 24268 4208
rect 22192 4131 22244 4140
rect 22192 4097 22226 4131
rect 22226 4097 22244 4131
rect 19064 4020 19116 4072
rect 19248 4063 19300 4072
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 21548 4020 21600 4072
rect 22192 4088 22244 4097
rect 23480 4088 23532 4140
rect 28080 4224 28132 4276
rect 30288 4224 30340 4276
rect 30380 4224 30432 4276
rect 32128 4224 32180 4276
rect 33416 4224 33468 4276
rect 33508 4224 33560 4276
rect 33968 4224 34020 4276
rect 35072 4224 35124 4276
rect 35900 4224 35952 4276
rect 24952 4131 25004 4140
rect 24952 4097 24959 4131
rect 24959 4097 25004 4131
rect 24952 4088 25004 4097
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25044 4088 25096 4097
rect 21732 4020 21784 4072
rect 18696 3952 18748 4004
rect 24124 4020 24176 4072
rect 24768 4020 24820 4072
rect 25412 4088 25464 4140
rect 26792 4131 26844 4140
rect 26792 4097 26801 4131
rect 26801 4097 26835 4131
rect 26835 4097 26844 4131
rect 26792 4088 26844 4097
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 27528 4088 27580 4140
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 28356 4131 28408 4140
rect 28356 4097 28360 4131
rect 28360 4097 28394 4131
rect 28394 4097 28408 4131
rect 28356 4088 28408 4097
rect 28448 4131 28500 4140
rect 28448 4097 28457 4131
rect 28457 4097 28491 4131
rect 28491 4097 28500 4131
rect 28448 4088 28500 4097
rect 19892 3884 19944 3936
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 21640 3927 21692 3936
rect 21640 3893 21649 3927
rect 21649 3893 21683 3927
rect 21683 3893 21692 3927
rect 21640 3884 21692 3893
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 25044 3952 25096 4004
rect 27252 4020 27304 4072
rect 28724 4131 28776 4140
rect 28724 4097 28733 4131
rect 28733 4097 28767 4131
rect 28767 4097 28776 4131
rect 28724 4088 28776 4097
rect 29184 4156 29236 4208
rect 29644 4156 29696 4208
rect 27160 3995 27212 4004
rect 27160 3961 27169 3995
rect 27169 3961 27203 3995
rect 27203 3961 27212 3995
rect 27160 3952 27212 3961
rect 28080 3952 28132 4004
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 28816 3995 28868 4004
rect 28816 3961 28825 3995
rect 28825 3961 28859 3995
rect 28859 3961 28868 3995
rect 28816 3952 28868 3961
rect 30012 4088 30064 4140
rect 30656 4131 30708 4140
rect 30656 4097 30665 4131
rect 30665 4097 30699 4131
rect 30699 4097 30708 4131
rect 30656 4088 30708 4097
rect 33876 4156 33928 4208
rect 34796 4199 34848 4208
rect 34796 4165 34830 4199
rect 34830 4165 34848 4199
rect 34796 4156 34848 4165
rect 30472 4063 30524 4072
rect 30472 4029 30481 4063
rect 30481 4029 30515 4063
rect 30515 4029 30524 4063
rect 30472 4020 30524 4029
rect 29644 3952 29696 4004
rect 29736 3952 29788 4004
rect 30380 3952 30432 4004
rect 33508 4131 33560 4140
rect 33508 4097 33517 4131
rect 33517 4097 33551 4131
rect 33551 4097 33560 4131
rect 33508 4088 33560 4097
rect 36360 4131 36412 4140
rect 36360 4097 36369 4131
rect 36369 4097 36403 4131
rect 36403 4097 36412 4131
rect 36360 4088 36412 4097
rect 36544 4088 36596 4140
rect 37648 4156 37700 4208
rect 39304 4224 39356 4276
rect 38384 4156 38436 4208
rect 38108 4131 38160 4140
rect 38108 4097 38115 4131
rect 38115 4097 38160 4131
rect 38108 4088 38160 4097
rect 38200 4131 38252 4140
rect 38200 4097 38209 4131
rect 38209 4097 38243 4131
rect 38243 4097 38252 4131
rect 38200 4088 38252 4097
rect 38660 4088 38712 4140
rect 36268 4020 36320 4072
rect 36912 4020 36964 4072
rect 39764 4131 39816 4140
rect 39764 4097 39773 4131
rect 39773 4097 39807 4131
rect 39807 4097 39816 4131
rect 39764 4088 39816 4097
rect 44640 4224 44692 4276
rect 44824 4224 44876 4276
rect 40132 4199 40184 4208
rect 40132 4165 40141 4199
rect 40141 4165 40175 4199
rect 40175 4165 40184 4199
rect 40132 4156 40184 4165
rect 39948 4020 40000 4072
rect 40684 4020 40736 4072
rect 41512 4156 41564 4208
rect 41420 4131 41472 4140
rect 41420 4097 41429 4131
rect 41429 4097 41463 4131
rect 41463 4097 41472 4131
rect 41420 4088 41472 4097
rect 41972 4131 42024 4140
rect 41972 4097 41981 4131
rect 41981 4097 42015 4131
rect 42015 4097 42024 4131
rect 41972 4088 42024 4097
rect 42248 4199 42300 4208
rect 42248 4165 42257 4199
rect 42257 4165 42291 4199
rect 42291 4165 42300 4199
rect 42248 4156 42300 4165
rect 43720 4199 43772 4208
rect 43720 4165 43729 4199
rect 43729 4165 43763 4199
rect 43763 4165 43772 4199
rect 43720 4156 43772 4165
rect 45100 4156 45152 4208
rect 45652 4224 45704 4276
rect 45468 4199 45520 4208
rect 45468 4165 45477 4199
rect 45477 4165 45511 4199
rect 45511 4165 45520 4199
rect 45468 4156 45520 4165
rect 30656 3927 30708 3936
rect 30656 3893 30665 3927
rect 30665 3893 30699 3927
rect 30699 3893 30708 3927
rect 30656 3884 30708 3893
rect 30748 3927 30800 3936
rect 30748 3893 30757 3927
rect 30757 3893 30791 3927
rect 30791 3893 30800 3927
rect 30748 3884 30800 3893
rect 31668 3927 31720 3936
rect 31668 3893 31677 3927
rect 31677 3893 31711 3927
rect 31711 3893 31720 3927
rect 31668 3884 31720 3893
rect 32864 3884 32916 3936
rect 35624 3884 35676 3936
rect 36452 3884 36504 3936
rect 36820 3927 36872 3936
rect 36820 3893 36829 3927
rect 36829 3893 36863 3927
rect 36863 3893 36872 3927
rect 36820 3884 36872 3893
rect 38752 3927 38804 3936
rect 38752 3893 38761 3927
rect 38761 3893 38795 3927
rect 38795 3893 38804 3927
rect 38752 3884 38804 3893
rect 39580 3927 39632 3936
rect 39580 3893 39589 3927
rect 39589 3893 39623 3927
rect 39623 3893 39632 3927
rect 39580 3884 39632 3893
rect 41512 3952 41564 4004
rect 43076 4063 43128 4072
rect 43076 4029 43085 4063
rect 43085 4029 43119 4063
rect 43119 4029 43128 4063
rect 43076 4020 43128 4029
rect 42984 3952 43036 4004
rect 45284 4121 45336 4140
rect 45284 4088 45288 4121
rect 45288 4088 45322 4121
rect 45322 4088 45336 4121
rect 46296 4156 46348 4208
rect 45744 4131 45796 4140
rect 45744 4097 45753 4131
rect 45753 4097 45787 4131
rect 45787 4097 45796 4131
rect 45744 4088 45796 4097
rect 46664 4156 46716 4208
rect 47032 4224 47084 4276
rect 47768 4224 47820 4276
rect 47952 4088 48004 4140
rect 48688 4224 48740 4276
rect 49884 4224 49936 4276
rect 50988 4156 51040 4208
rect 53564 4267 53616 4276
rect 53564 4233 53573 4267
rect 53573 4233 53607 4267
rect 53607 4233 53616 4267
rect 53564 4224 53616 4233
rect 49240 4088 49292 4140
rect 49424 4131 49476 4140
rect 49424 4097 49433 4131
rect 49433 4097 49467 4131
rect 49467 4097 49476 4131
rect 49424 4088 49476 4097
rect 50436 4088 50488 4140
rect 50712 4088 50764 4140
rect 51172 4131 51224 4140
rect 51172 4097 51181 4131
rect 51181 4097 51215 4131
rect 51215 4097 51224 4131
rect 51172 4088 51224 4097
rect 44088 3952 44140 4004
rect 44732 4020 44784 4072
rect 45008 4063 45060 4072
rect 45008 4029 45017 4063
rect 45017 4029 45051 4063
rect 45051 4029 45060 4063
rect 45008 4020 45060 4029
rect 47124 4020 47176 4072
rect 47492 4020 47544 4072
rect 48964 4063 49016 4072
rect 48964 4029 48973 4063
rect 48973 4029 49007 4063
rect 49007 4029 49016 4063
rect 48964 4020 49016 4029
rect 40684 3884 40736 3936
rect 41788 3884 41840 3936
rect 43444 3927 43496 3936
rect 43444 3893 43453 3927
rect 43453 3893 43487 3927
rect 43487 3893 43496 3927
rect 43444 3884 43496 3893
rect 43904 3927 43956 3936
rect 43904 3893 43913 3927
rect 43913 3893 43947 3927
rect 43947 3893 43956 3927
rect 43904 3884 43956 3893
rect 44180 3927 44232 3936
rect 44180 3893 44189 3927
rect 44189 3893 44223 3927
rect 44223 3893 44232 3927
rect 44180 3884 44232 3893
rect 49792 4020 49844 4072
rect 52000 4088 52052 4140
rect 53932 4224 53984 4276
rect 56324 4224 56376 4276
rect 56600 4224 56652 4276
rect 52460 4088 52512 4140
rect 52828 4088 52880 4140
rect 53380 4131 53432 4140
rect 53380 4097 53389 4131
rect 53389 4097 53423 4131
rect 53423 4097 53432 4131
rect 53380 4088 53432 4097
rect 54116 4131 54168 4140
rect 54116 4097 54125 4131
rect 54125 4097 54159 4131
rect 54159 4097 54168 4131
rect 54116 4088 54168 4097
rect 54300 4131 54352 4140
rect 54300 4097 54309 4131
rect 54309 4097 54343 4131
rect 54343 4097 54352 4131
rect 54300 4088 54352 4097
rect 54576 4088 54628 4140
rect 57152 4224 57204 4276
rect 56968 4131 57020 4140
rect 56968 4097 56972 4131
rect 56972 4097 57006 4131
rect 57006 4097 57020 4131
rect 51356 3952 51408 4004
rect 54852 4020 54904 4072
rect 56968 4088 57020 4097
rect 57244 4156 57296 4208
rect 57336 4199 57388 4208
rect 57336 4165 57345 4199
rect 57345 4165 57379 4199
rect 57379 4165 57388 4199
rect 57336 4156 57388 4165
rect 56876 4020 56928 4072
rect 57428 4131 57480 4140
rect 57428 4097 57437 4131
rect 57437 4097 57471 4131
rect 57471 4097 57480 4131
rect 57428 4088 57480 4097
rect 45836 3884 45888 3936
rect 46480 3884 46532 3936
rect 47768 3927 47820 3936
rect 47768 3893 47777 3927
rect 47777 3893 47811 3927
rect 47811 3893 47820 3927
rect 47768 3884 47820 3893
rect 48044 3884 48096 3936
rect 50252 3884 50304 3936
rect 52368 3927 52420 3936
rect 52368 3893 52377 3927
rect 52377 3893 52411 3927
rect 52411 3893 52420 3927
rect 52368 3884 52420 3893
rect 54300 3927 54352 3936
rect 54300 3893 54309 3927
rect 54309 3893 54343 3927
rect 54343 3893 54352 3927
rect 54300 3884 54352 3893
rect 54576 3927 54628 3936
rect 54576 3893 54585 3927
rect 54585 3893 54619 3927
rect 54619 3893 54628 3927
rect 54576 3884 54628 3893
rect 55404 3927 55456 3936
rect 55404 3893 55413 3927
rect 55413 3893 55447 3927
rect 55447 3893 55456 3927
rect 55404 3884 55456 3893
rect 57612 3927 57664 3936
rect 57612 3893 57621 3927
rect 57621 3893 57655 3927
rect 57655 3893 57664 3927
rect 57612 3884 57664 3893
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 22616 3782 22668 3834
rect 22680 3782 22732 3834
rect 22744 3782 22796 3834
rect 22808 3782 22860 3834
rect 22872 3782 22924 3834
rect 37060 3782 37112 3834
rect 37124 3782 37176 3834
rect 37188 3782 37240 3834
rect 37252 3782 37304 3834
rect 37316 3782 37368 3834
rect 51504 3782 51556 3834
rect 51568 3782 51620 3834
rect 51632 3782 51684 3834
rect 51696 3782 51748 3834
rect 51760 3782 51812 3834
rect 2964 3680 3016 3732
rect 6184 3723 6236 3732
rect 6184 3689 6193 3723
rect 6193 3689 6227 3723
rect 6227 3689 6236 3723
rect 6184 3680 6236 3689
rect 6276 3723 6328 3732
rect 6276 3689 6285 3723
rect 6285 3689 6319 3723
rect 6319 3689 6328 3723
rect 6276 3680 6328 3689
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 11060 3680 11112 3732
rect 9956 3612 10008 3664
rect 13452 3680 13504 3732
rect 13544 3680 13596 3732
rect 14372 3680 14424 3732
rect 16488 3680 16540 3732
rect 17592 3723 17644 3732
rect 17592 3689 17601 3723
rect 17601 3689 17635 3723
rect 17635 3689 17644 3723
rect 17592 3680 17644 3689
rect 18052 3680 18104 3732
rect 18696 3680 18748 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 20812 3680 20864 3732
rect 3056 3544 3108 3596
rect 4068 3544 4120 3596
rect 3332 3519 3384 3528
rect 3332 3485 3341 3519
rect 3341 3485 3375 3519
rect 3375 3485 3384 3519
rect 3332 3476 3384 3485
rect 3516 3476 3568 3528
rect 3700 3476 3752 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 6368 3544 6420 3596
rect 1768 3408 1820 3460
rect 2136 3340 2188 3392
rect 3976 3408 4028 3460
rect 5356 3408 5408 3460
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 8852 3476 8904 3528
rect 14832 3612 14884 3664
rect 15292 3612 15344 3664
rect 24124 3680 24176 3732
rect 25136 3680 25188 3732
rect 25504 3680 25556 3732
rect 14280 3544 14332 3596
rect 10048 3476 10100 3528
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 7564 3408 7616 3460
rect 8760 3408 8812 3460
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 8668 3340 8720 3392
rect 9496 3408 9548 3460
rect 10508 3451 10560 3460
rect 10508 3417 10517 3451
rect 10517 3417 10551 3451
rect 10551 3417 10560 3451
rect 10508 3408 10560 3417
rect 10600 3408 10652 3460
rect 9404 3340 9456 3392
rect 10232 3340 10284 3392
rect 12072 3340 12124 3392
rect 13360 3408 13412 3460
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14740 3476 14792 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 17408 3544 17460 3596
rect 14556 3408 14608 3460
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 18604 3408 18656 3460
rect 12256 3340 12308 3392
rect 15200 3340 15252 3392
rect 15936 3340 15988 3392
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 17592 3340 17644 3392
rect 19984 3340 20036 3392
rect 20444 3408 20496 3460
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 22468 3544 22520 3596
rect 22284 3476 22336 3528
rect 21364 3451 21416 3460
rect 21364 3417 21398 3451
rect 21398 3417 21416 3451
rect 21364 3408 21416 3417
rect 21640 3408 21692 3460
rect 22744 3476 22796 3528
rect 24124 3408 24176 3460
rect 26240 3451 26292 3460
rect 26240 3417 26274 3451
rect 26274 3417 26292 3451
rect 26240 3408 26292 3417
rect 27712 3476 27764 3528
rect 28816 3680 28868 3732
rect 30748 3680 30800 3732
rect 31668 3680 31720 3732
rect 31484 3587 31536 3596
rect 31484 3553 31493 3587
rect 31493 3553 31527 3587
rect 31527 3553 31536 3587
rect 31484 3544 31536 3553
rect 33508 3680 33560 3732
rect 31392 3519 31444 3528
rect 31392 3485 31401 3519
rect 31401 3485 31435 3519
rect 31435 3485 31444 3519
rect 31392 3476 31444 3485
rect 34612 3612 34664 3664
rect 35808 3519 35860 3528
rect 38200 3680 38252 3732
rect 38568 3680 38620 3732
rect 39764 3680 39816 3732
rect 40040 3680 40092 3732
rect 44824 3723 44876 3732
rect 44824 3689 44833 3723
rect 44833 3689 44867 3723
rect 44867 3689 44876 3723
rect 44824 3680 44876 3689
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 27344 3383 27396 3392
rect 27344 3349 27353 3383
rect 27353 3349 27387 3383
rect 27387 3349 27396 3383
rect 27344 3340 27396 3349
rect 28448 3408 28500 3460
rect 30380 3408 30432 3460
rect 30840 3408 30892 3460
rect 34888 3408 34940 3460
rect 35164 3408 35216 3460
rect 29276 3383 29328 3392
rect 29276 3349 29285 3383
rect 29285 3349 29319 3383
rect 29319 3349 29328 3383
rect 29276 3340 29328 3349
rect 33692 3340 33744 3392
rect 35348 3383 35400 3392
rect 35348 3349 35357 3383
rect 35357 3349 35391 3383
rect 35391 3349 35400 3383
rect 35348 3340 35400 3349
rect 35808 3485 35822 3519
rect 35822 3485 35856 3519
rect 35856 3485 35860 3519
rect 35808 3476 35860 3485
rect 37464 3476 37516 3528
rect 40868 3544 40920 3596
rect 45928 3680 45980 3732
rect 46940 3655 46992 3664
rect 46940 3621 46949 3655
rect 46949 3621 46983 3655
rect 46983 3621 46992 3655
rect 46940 3612 46992 3621
rect 50160 3680 50212 3732
rect 53840 3680 53892 3732
rect 56600 3680 56652 3732
rect 57152 3680 57204 3732
rect 58256 3680 58308 3732
rect 49240 3655 49292 3664
rect 49240 3621 49249 3655
rect 49249 3621 49283 3655
rect 49283 3621 49292 3655
rect 49240 3612 49292 3621
rect 35624 3451 35676 3460
rect 35624 3417 35633 3451
rect 35633 3417 35667 3451
rect 35667 3417 35676 3451
rect 35624 3408 35676 3417
rect 36820 3408 36872 3460
rect 38752 3408 38804 3460
rect 35900 3340 35952 3392
rect 36176 3340 36228 3392
rect 38108 3340 38160 3392
rect 39396 3340 39448 3392
rect 39488 3383 39540 3392
rect 39488 3349 39497 3383
rect 39497 3349 39531 3383
rect 39531 3349 39540 3383
rect 39488 3340 39540 3349
rect 40132 3451 40184 3460
rect 40132 3417 40166 3451
rect 40166 3417 40184 3451
rect 40132 3408 40184 3417
rect 42616 3408 42668 3460
rect 43168 3519 43220 3528
rect 43168 3485 43177 3519
rect 43177 3485 43211 3519
rect 43211 3485 43220 3519
rect 43168 3476 43220 3485
rect 43536 3476 43588 3528
rect 44640 3476 44692 3528
rect 45836 3476 45888 3528
rect 47124 3519 47176 3528
rect 47124 3485 47133 3519
rect 47133 3485 47167 3519
rect 47167 3485 47176 3519
rect 47124 3476 47176 3485
rect 48044 3519 48096 3528
rect 48044 3485 48078 3519
rect 48078 3485 48096 3519
rect 48044 3476 48096 3485
rect 49056 3476 49108 3528
rect 50068 3476 50120 3528
rect 52368 3476 52420 3528
rect 53012 3519 53064 3528
rect 53012 3485 53021 3519
rect 53021 3485 53055 3519
rect 53055 3485 53064 3519
rect 53012 3476 53064 3485
rect 43352 3451 43404 3460
rect 43352 3417 43361 3451
rect 43361 3417 43395 3451
rect 43395 3417 43404 3451
rect 43352 3408 43404 3417
rect 46204 3408 46256 3460
rect 47492 3408 47544 3460
rect 48964 3408 49016 3460
rect 51172 3408 51224 3460
rect 40500 3340 40552 3392
rect 41236 3383 41288 3392
rect 41236 3349 41245 3383
rect 41245 3349 41279 3383
rect 41279 3349 41288 3383
rect 41236 3340 41288 3349
rect 41972 3340 42024 3392
rect 42340 3340 42392 3392
rect 42708 3340 42760 3392
rect 45008 3340 45060 3392
rect 46572 3340 46624 3392
rect 48596 3340 48648 3392
rect 49148 3383 49200 3392
rect 49148 3349 49157 3383
rect 49157 3349 49191 3383
rect 49191 3349 49200 3383
rect 49148 3340 49200 3349
rect 52184 3408 52236 3460
rect 52552 3340 52604 3392
rect 53104 3383 53156 3392
rect 53104 3349 53113 3383
rect 53113 3349 53147 3383
rect 53147 3349 53156 3383
rect 53104 3340 53156 3349
rect 54300 3408 54352 3460
rect 55128 3519 55180 3528
rect 55128 3485 55137 3519
rect 55137 3485 55171 3519
rect 55171 3485 55180 3519
rect 55128 3476 55180 3485
rect 55220 3476 55272 3528
rect 55404 3408 55456 3460
rect 54944 3340 54996 3392
rect 56876 3340 56928 3392
rect 58164 3408 58216 3460
rect 15394 3238 15446 3290
rect 15458 3238 15510 3290
rect 15522 3238 15574 3290
rect 15586 3238 15638 3290
rect 15650 3238 15702 3290
rect 29838 3238 29890 3290
rect 29902 3238 29954 3290
rect 29966 3238 30018 3290
rect 30030 3238 30082 3290
rect 30094 3238 30146 3290
rect 44282 3238 44334 3290
rect 44346 3238 44398 3290
rect 44410 3238 44462 3290
rect 44474 3238 44526 3290
rect 44538 3238 44590 3290
rect 58726 3238 58778 3290
rect 58790 3238 58842 3290
rect 58854 3238 58906 3290
rect 58918 3238 58970 3290
rect 58982 3238 59034 3290
rect 1768 3136 1820 3188
rect 2228 3136 2280 3188
rect 3700 3136 3752 3188
rect 4528 3136 4580 3188
rect 4712 3136 4764 3188
rect 7748 3136 7800 3188
rect 8024 3136 8076 3188
rect 8116 3136 8168 3188
rect 8576 3136 8628 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 9220 3136 9272 3188
rect 9404 3136 9456 3188
rect 3516 3068 3568 3120
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 2044 2932 2096 2984
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 4160 2932 4212 2984
rect 3700 2864 3752 2916
rect 3976 2864 4028 2916
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 9680 3068 9732 3120
rect 10600 3136 10652 3188
rect 10876 3136 10928 3188
rect 10232 3068 10284 3120
rect 14372 3136 14424 3188
rect 15384 3136 15436 3188
rect 15752 3136 15804 3188
rect 13084 3068 13136 3120
rect 14188 3068 14240 3120
rect 14648 3068 14700 3120
rect 16212 3136 16264 3188
rect 16304 3136 16356 3188
rect 16488 3136 16540 3188
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 6736 2864 6788 2916
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 9956 3043 10008 3052
rect 9956 3009 9970 3043
rect 9970 3009 10004 3043
rect 10004 3009 10008 3043
rect 9956 3000 10008 3009
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10692 3000 10744 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 14464 3000 14516 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 10232 2932 10284 2984
rect 11980 2932 12032 2984
rect 13636 2932 13688 2984
rect 16580 3068 16632 3120
rect 16672 3068 16724 3120
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17040 3136 17092 3188
rect 19524 3136 19576 3188
rect 20076 3136 20128 3188
rect 20996 3136 21048 3188
rect 21548 3136 21600 3188
rect 23388 3136 23440 3188
rect 24124 3136 24176 3188
rect 25044 3136 25096 3188
rect 25228 3136 25280 3188
rect 26516 3136 26568 3188
rect 29276 3136 29328 3188
rect 30656 3136 30708 3188
rect 31392 3136 31444 3188
rect 32864 3136 32916 3188
rect 34336 3136 34388 3188
rect 34796 3136 34848 3188
rect 34888 3136 34940 3188
rect 35348 3136 35400 3188
rect 35716 3136 35768 3188
rect 37004 3179 37056 3188
rect 37004 3145 37013 3179
rect 37013 3145 37047 3179
rect 37047 3145 37056 3179
rect 37004 3136 37056 3145
rect 38200 3136 38252 3188
rect 38936 3136 38988 3188
rect 39396 3136 39448 3188
rect 40684 3136 40736 3188
rect 41236 3136 41288 3188
rect 41420 3136 41472 3188
rect 43168 3136 43220 3188
rect 46204 3136 46256 3188
rect 46940 3179 46992 3188
rect 46940 3145 46949 3179
rect 46949 3145 46983 3179
rect 46983 3145 46992 3179
rect 46940 3136 46992 3145
rect 47124 3136 47176 3188
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17316 3000 17368 3052
rect 10324 2907 10376 2916
rect 10324 2873 10333 2907
rect 10333 2873 10367 2907
rect 10367 2873 10376 2907
rect 10324 2864 10376 2873
rect 3516 2796 3568 2848
rect 7104 2796 7156 2848
rect 7840 2796 7892 2848
rect 16028 2864 16080 2916
rect 19064 3000 19116 3052
rect 21088 3043 21140 3052
rect 21088 3009 21097 3043
rect 21097 3009 21131 3043
rect 21131 3009 21140 3043
rect 21088 3000 21140 3009
rect 22744 3068 22796 3120
rect 24308 3068 24360 3120
rect 24676 3068 24728 3120
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 19156 2932 19208 2984
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 21640 3043 21692 3052
rect 21640 3009 21649 3043
rect 21649 3009 21683 3043
rect 21683 3009 21692 3043
rect 21640 3000 21692 3009
rect 21824 3000 21876 3052
rect 23296 3000 23348 3052
rect 24032 3000 24084 3052
rect 20628 2864 20680 2916
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 24216 3000 24268 3009
rect 30932 3043 30984 3052
rect 30932 3009 30941 3043
rect 30941 3009 30975 3043
rect 30975 3009 30984 3043
rect 30932 3000 30984 3009
rect 31208 3043 31260 3052
rect 31208 3009 31217 3043
rect 31217 3009 31251 3043
rect 31251 3009 31260 3043
rect 31208 3000 31260 3009
rect 33416 3043 33468 3052
rect 24676 2975 24728 2984
rect 24676 2941 24685 2975
rect 24685 2941 24719 2975
rect 24719 2941 24728 2975
rect 24676 2932 24728 2941
rect 23572 2864 23624 2916
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 26700 2864 26752 2916
rect 26884 2864 26936 2916
rect 28540 2975 28592 2984
rect 28540 2941 28549 2975
rect 28549 2941 28583 2975
rect 28583 2941 28592 2975
rect 28540 2932 28592 2941
rect 29368 2932 29420 2984
rect 30564 2932 30616 2984
rect 31852 2932 31904 2984
rect 18788 2796 18840 2848
rect 21732 2796 21784 2848
rect 29092 2839 29144 2848
rect 29092 2805 29101 2839
rect 29101 2805 29135 2839
rect 29135 2805 29144 2839
rect 29092 2796 29144 2805
rect 31944 2839 31996 2848
rect 31944 2805 31953 2839
rect 31953 2805 31987 2839
rect 31987 2805 31996 2839
rect 31944 2796 31996 2805
rect 33416 3009 33449 3043
rect 33449 3009 33468 3043
rect 33416 3000 33468 3009
rect 33140 2932 33192 2984
rect 33600 2932 33652 2984
rect 35072 2932 35124 2984
rect 35256 2975 35308 2984
rect 35256 2941 35265 2975
rect 35265 2941 35299 2975
rect 35299 2941 35308 2975
rect 35256 2932 35308 2941
rect 36544 3043 36596 3052
rect 36544 3009 36553 3043
rect 36553 3009 36587 3043
rect 36587 3009 36596 3043
rect 36544 3000 36596 3009
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 39304 3068 39356 3120
rect 39212 3043 39264 3052
rect 39212 3009 39221 3043
rect 39221 3009 39255 3043
rect 39255 3009 39264 3043
rect 39212 3000 39264 3009
rect 32956 2864 33008 2916
rect 36176 2864 36228 2916
rect 34704 2796 34756 2848
rect 37648 2932 37700 2984
rect 40224 3000 40276 3052
rect 43628 3000 43680 3052
rect 44824 3000 44876 3052
rect 46664 3068 46716 3120
rect 46756 3111 46808 3120
rect 46756 3077 46765 3111
rect 46765 3077 46799 3111
rect 46799 3077 46808 3111
rect 46756 3068 46808 3077
rect 46848 3068 46900 3120
rect 48320 3111 48372 3120
rect 48320 3077 48329 3111
rect 48329 3077 48363 3111
rect 48363 3077 48372 3111
rect 48320 3068 48372 3077
rect 48688 3136 48740 3188
rect 40684 2932 40736 2984
rect 41788 2932 41840 2984
rect 43996 2932 44048 2984
rect 45100 2932 45152 2984
rect 46572 2932 46624 2984
rect 48596 3111 48648 3120
rect 48596 3077 48605 3111
rect 48605 3077 48639 3111
rect 48639 3077 48648 3111
rect 48596 3068 48648 3077
rect 48964 3136 49016 3188
rect 51908 3136 51960 3188
rect 51080 3068 51132 3120
rect 52552 3068 52604 3120
rect 53104 3068 53156 3120
rect 53564 3068 53616 3120
rect 53656 3111 53708 3120
rect 53656 3077 53665 3111
rect 53665 3077 53699 3111
rect 53699 3077 53708 3111
rect 53656 3068 53708 3077
rect 46756 2932 46808 2984
rect 49056 3000 49108 3052
rect 49148 3043 49200 3052
rect 49148 3009 49157 3043
rect 49157 3009 49191 3043
rect 49191 3009 49200 3043
rect 49148 3000 49200 3009
rect 51356 3000 51408 3052
rect 46940 2864 46992 2916
rect 48964 2932 49016 2984
rect 50068 2932 50120 2984
rect 49424 2864 49476 2916
rect 50988 2864 51040 2916
rect 52000 3000 52052 3052
rect 51724 2932 51776 2984
rect 53840 3033 53892 3052
rect 58532 3179 58584 3188
rect 58532 3145 58541 3179
rect 58541 3145 58575 3179
rect 58575 3145 58584 3179
rect 58532 3136 58584 3145
rect 53840 3000 53885 3033
rect 53885 3000 53892 3033
rect 57704 3043 57756 3052
rect 57704 3009 57713 3043
rect 57713 3009 57747 3043
rect 57747 3009 57756 3043
rect 57704 3000 57756 3009
rect 53748 2975 53800 2984
rect 53748 2941 53757 2975
rect 53757 2941 53791 2975
rect 53791 2941 53800 2975
rect 53748 2932 53800 2941
rect 54208 2932 54260 2984
rect 55036 2932 55088 2984
rect 57244 2975 57296 2984
rect 57244 2941 57253 2975
rect 57253 2941 57287 2975
rect 57287 2941 57296 2975
rect 57244 2932 57296 2941
rect 58348 2932 58400 2984
rect 38660 2796 38712 2848
rect 39764 2796 39816 2848
rect 43444 2796 43496 2848
rect 45560 2796 45612 2848
rect 46296 2796 46348 2848
rect 51172 2839 51224 2848
rect 51172 2805 51181 2839
rect 51181 2805 51215 2839
rect 51215 2805 51224 2839
rect 51172 2796 51224 2805
rect 56968 2796 57020 2848
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 22616 2694 22668 2746
rect 22680 2694 22732 2746
rect 22744 2694 22796 2746
rect 22808 2694 22860 2746
rect 22872 2694 22924 2746
rect 37060 2694 37112 2746
rect 37124 2694 37176 2746
rect 37188 2694 37240 2746
rect 37252 2694 37304 2746
rect 37316 2694 37368 2746
rect 51504 2694 51556 2746
rect 51568 2694 51620 2746
rect 51632 2694 51684 2746
rect 51696 2694 51748 2746
rect 51760 2694 51812 2746
rect 4896 2592 4948 2644
rect 7656 2592 7708 2644
rect 10140 2592 10192 2644
rect 10232 2592 10284 2644
rect 11796 2592 11848 2644
rect 12348 2592 12400 2644
rect 14832 2592 14884 2644
rect 16028 2592 16080 2644
rect 17132 2592 17184 2644
rect 20720 2592 20772 2644
rect 21088 2592 21140 2644
rect 24400 2635 24452 2644
rect 24400 2601 24409 2635
rect 24409 2601 24443 2635
rect 24443 2601 24452 2635
rect 24400 2592 24452 2601
rect 25412 2592 25464 2644
rect 27620 2592 27672 2644
rect 29368 2592 29420 2644
rect 30380 2592 30432 2644
rect 30932 2592 30984 2644
rect 33140 2592 33192 2644
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 2412 2456 2464 2508
rect 1952 2388 2004 2440
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 4804 2388 4856 2440
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 5264 2363 5316 2372
rect 5264 2329 5273 2363
rect 5273 2329 5307 2363
rect 5307 2329 5316 2363
rect 5264 2320 5316 2329
rect 6000 2252 6052 2304
rect 23480 2524 23532 2576
rect 27528 2524 27580 2576
rect 36084 2592 36136 2644
rect 36820 2592 36872 2644
rect 38568 2592 38620 2644
rect 39212 2592 39264 2644
rect 40132 2592 40184 2644
rect 40500 2592 40552 2644
rect 41512 2592 41564 2644
rect 43812 2592 43864 2644
rect 44180 2592 44232 2644
rect 47216 2635 47268 2644
rect 47216 2601 47225 2635
rect 47225 2601 47259 2635
rect 47259 2601 47268 2635
rect 47216 2592 47268 2601
rect 49792 2635 49844 2644
rect 49792 2601 49801 2635
rect 49801 2601 49835 2635
rect 49835 2601 49844 2635
rect 49792 2592 49844 2601
rect 50160 2635 50212 2644
rect 50160 2601 50169 2635
rect 50169 2601 50203 2635
rect 50203 2601 50212 2635
rect 50160 2592 50212 2601
rect 51172 2592 51224 2644
rect 52000 2592 52052 2644
rect 53380 2592 53432 2644
rect 55128 2635 55180 2644
rect 55128 2601 55137 2635
rect 55137 2601 55171 2635
rect 55171 2601 55180 2635
rect 55128 2592 55180 2601
rect 56600 2592 56652 2644
rect 56784 2592 56836 2644
rect 57428 2592 57480 2644
rect 8392 2456 8444 2508
rect 9772 2456 9824 2508
rect 14188 2456 14240 2508
rect 15292 2456 15344 2508
rect 15844 2499 15896 2508
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 17868 2456 17920 2508
rect 19984 2456 20036 2508
rect 7012 2388 7064 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 12164 2388 12216 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 13544 2388 13596 2440
rect 7564 2363 7616 2372
rect 7564 2329 7573 2363
rect 7573 2329 7607 2363
rect 7607 2329 7616 2363
rect 7564 2320 7616 2329
rect 11060 2252 11112 2304
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 19432 2388 19484 2440
rect 20076 2388 20128 2440
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 21824 2456 21876 2508
rect 22468 2456 22520 2508
rect 22192 2388 22244 2440
rect 22744 2456 22796 2508
rect 25872 2499 25924 2508
rect 25872 2465 25881 2499
rect 25881 2465 25915 2499
rect 25915 2465 25924 2499
rect 25872 2456 25924 2465
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2388 25280 2440
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 27712 2456 27764 2508
rect 31024 2499 31076 2508
rect 31024 2465 31033 2499
rect 31033 2465 31067 2499
rect 31067 2465 31076 2499
rect 31024 2456 31076 2465
rect 31116 2456 31168 2508
rect 35624 2524 35676 2576
rect 44732 2524 44784 2576
rect 27252 2431 27304 2440
rect 27252 2397 27261 2431
rect 27261 2397 27295 2431
rect 27295 2397 27304 2431
rect 27252 2388 27304 2397
rect 27344 2388 27396 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 15292 2320 15344 2372
rect 29092 2388 29144 2440
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 30196 2388 30248 2440
rect 30840 2388 30892 2440
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 33692 2431 33744 2440
rect 33692 2397 33701 2431
rect 33701 2397 33735 2431
rect 33735 2397 33744 2431
rect 33692 2388 33744 2397
rect 32404 2320 32456 2372
rect 33968 2363 34020 2372
rect 33968 2329 33977 2363
rect 33977 2329 34011 2363
rect 34011 2329 34020 2363
rect 33968 2320 34020 2329
rect 35072 2456 35124 2508
rect 35808 2456 35860 2508
rect 38660 2456 38712 2508
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 35900 2388 35952 2397
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 36820 2388 36872 2440
rect 36912 2388 36964 2440
rect 38752 2431 38804 2440
rect 38752 2397 38761 2431
rect 38761 2397 38795 2431
rect 38795 2397 38804 2431
rect 38752 2388 38804 2397
rect 39028 2456 39080 2508
rect 42616 2456 42668 2508
rect 45560 2499 45612 2508
rect 45560 2465 45569 2499
rect 45569 2465 45603 2499
rect 45603 2465 45612 2499
rect 45560 2456 45612 2465
rect 47676 2456 47728 2508
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 39948 2431 40000 2440
rect 39948 2397 39957 2431
rect 39957 2397 39991 2431
rect 39991 2397 40000 2431
rect 39948 2388 40000 2397
rect 40132 2388 40184 2440
rect 42248 2431 42300 2440
rect 42248 2397 42257 2431
rect 42257 2397 42291 2431
rect 42291 2397 42300 2431
rect 42248 2388 42300 2397
rect 42340 2388 42392 2440
rect 43168 2388 43220 2440
rect 44824 2431 44876 2440
rect 44824 2397 44833 2431
rect 44833 2397 44867 2431
rect 44867 2397 44876 2431
rect 44824 2388 44876 2397
rect 46572 2388 46624 2440
rect 34520 2320 34572 2372
rect 45652 2320 45704 2372
rect 47952 2388 48004 2440
rect 48412 2388 48464 2440
rect 49700 2388 49752 2440
rect 52092 2431 52144 2440
rect 52092 2397 52101 2431
rect 52101 2397 52135 2431
rect 52135 2397 52144 2431
rect 52092 2388 52144 2397
rect 52460 2456 52512 2508
rect 52552 2388 52604 2440
rect 53380 2388 53432 2440
rect 56784 2456 56836 2508
rect 47860 2320 47912 2372
rect 50804 2320 50856 2372
rect 52920 2320 52972 2372
rect 56876 2431 56928 2440
rect 56876 2397 56885 2431
rect 56885 2397 56919 2431
rect 56919 2397 56928 2431
rect 56876 2388 56928 2397
rect 56968 2388 57020 2440
rect 55680 2320 55732 2372
rect 56324 2320 56376 2372
rect 15200 2252 15252 2304
rect 15394 2150 15446 2202
rect 15458 2150 15510 2202
rect 15522 2150 15574 2202
rect 15586 2150 15638 2202
rect 15650 2150 15702 2202
rect 29838 2150 29890 2202
rect 29902 2150 29954 2202
rect 29966 2150 30018 2202
rect 30030 2150 30082 2202
rect 30094 2150 30146 2202
rect 44282 2150 44334 2202
rect 44346 2150 44398 2202
rect 44410 2150 44462 2202
rect 44474 2150 44526 2202
rect 44538 2150 44590 2202
rect 58726 2150 58778 2202
rect 58790 2150 58842 2202
rect 58854 2150 58906 2202
rect 58918 2150 58970 2202
rect 58982 2150 59034 2202
rect 26332 2048 26384 2100
rect 26976 2048 27028 2100
<< metal2 >>
rect 8172 27772 8480 27781
rect 8172 27770 8178 27772
rect 8234 27770 8258 27772
rect 8314 27770 8338 27772
rect 8394 27770 8418 27772
rect 8474 27770 8480 27772
rect 8234 27718 8236 27770
rect 8416 27718 8418 27770
rect 8172 27716 8178 27718
rect 8234 27716 8258 27718
rect 8314 27716 8338 27718
rect 8394 27716 8418 27718
rect 8474 27716 8480 27718
rect 8172 27707 8480 27716
rect 22616 27772 22924 27781
rect 22616 27770 22622 27772
rect 22678 27770 22702 27772
rect 22758 27770 22782 27772
rect 22838 27770 22862 27772
rect 22918 27770 22924 27772
rect 22678 27718 22680 27770
rect 22860 27718 22862 27770
rect 22616 27716 22622 27718
rect 22678 27716 22702 27718
rect 22758 27716 22782 27718
rect 22838 27716 22862 27718
rect 22918 27716 22924 27718
rect 22616 27707 22924 27716
rect 37060 27772 37368 27781
rect 37060 27770 37066 27772
rect 37122 27770 37146 27772
rect 37202 27770 37226 27772
rect 37282 27770 37306 27772
rect 37362 27770 37368 27772
rect 37122 27718 37124 27770
rect 37304 27718 37306 27770
rect 37060 27716 37066 27718
rect 37122 27716 37146 27718
rect 37202 27716 37226 27718
rect 37282 27716 37306 27718
rect 37362 27716 37368 27718
rect 37060 27707 37368 27716
rect 51504 27772 51812 27781
rect 51504 27770 51510 27772
rect 51566 27770 51590 27772
rect 51646 27770 51670 27772
rect 51726 27770 51750 27772
rect 51806 27770 51812 27772
rect 51566 27718 51568 27770
rect 51748 27718 51750 27770
rect 51504 27716 51510 27718
rect 51566 27716 51590 27718
rect 51646 27716 51670 27718
rect 51726 27716 51750 27718
rect 51806 27716 51812 27718
rect 51504 27707 51812 27716
rect 51356 27464 51408 27470
rect 51356 27406 51408 27412
rect 15394 27228 15702 27237
rect 15394 27226 15400 27228
rect 15456 27226 15480 27228
rect 15536 27226 15560 27228
rect 15616 27226 15640 27228
rect 15696 27226 15702 27228
rect 15456 27174 15458 27226
rect 15638 27174 15640 27226
rect 15394 27172 15400 27174
rect 15456 27172 15480 27174
rect 15536 27172 15560 27174
rect 15616 27172 15640 27174
rect 15696 27172 15702 27174
rect 15394 27163 15702 27172
rect 29838 27228 30146 27237
rect 29838 27226 29844 27228
rect 29900 27226 29924 27228
rect 29980 27226 30004 27228
rect 30060 27226 30084 27228
rect 30140 27226 30146 27228
rect 29900 27174 29902 27226
rect 30082 27174 30084 27226
rect 29838 27172 29844 27174
rect 29900 27172 29924 27174
rect 29980 27172 30004 27174
rect 30060 27172 30084 27174
rect 30140 27172 30146 27174
rect 29838 27163 30146 27172
rect 44282 27228 44590 27237
rect 44282 27226 44288 27228
rect 44344 27226 44368 27228
rect 44424 27226 44448 27228
rect 44504 27226 44528 27228
rect 44584 27226 44590 27228
rect 44344 27174 44346 27226
rect 44526 27174 44528 27226
rect 44282 27172 44288 27174
rect 44344 27172 44368 27174
rect 44424 27172 44448 27174
rect 44504 27172 44528 27174
rect 44584 27172 44590 27174
rect 44282 27163 44590 27172
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28724 26920 28776 26926
rect 28724 26862 28776 26868
rect 30196 26920 30248 26926
rect 30196 26862 30248 26868
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 8172 26684 8480 26693
rect 8172 26682 8178 26684
rect 8234 26682 8258 26684
rect 8314 26682 8338 26684
rect 8394 26682 8418 26684
rect 8474 26682 8480 26684
rect 8234 26630 8236 26682
rect 8416 26630 8418 26682
rect 8172 26628 8178 26630
rect 8234 26628 8258 26630
rect 8314 26628 8338 26630
rect 8394 26628 8418 26630
rect 8474 26628 8480 26630
rect 8172 26619 8480 26628
rect 17328 26586 17356 26862
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 27804 26784 27856 26790
rect 27804 26726 27856 26732
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 25906 15148 26182
rect 15394 26140 15702 26149
rect 15394 26138 15400 26140
rect 15456 26138 15480 26140
rect 15536 26138 15560 26140
rect 15616 26138 15640 26140
rect 15696 26138 15702 26140
rect 15456 26086 15458 26138
rect 15638 26086 15640 26138
rect 15394 26084 15400 26086
rect 15456 26084 15480 26086
rect 15536 26084 15560 26086
rect 15616 26084 15640 26086
rect 15696 26084 15702 26086
rect 15394 26075 15702 26084
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25294 6500 25638
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4908 24886 4936 25094
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24274 4016 24550
rect 5552 24410 5580 25230
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5920 24274 5948 24754
rect 6380 24682 6408 25230
rect 7024 24954 7052 25774
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 24954 7144 25094
rect 7208 24954 7236 25638
rect 7760 25498 7788 25774
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 6368 24676 6420 24682
rect 6368 24618 6420 24624
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6196 24410 6224 24550
rect 7208 24410 7236 24890
rect 7944 24886 7972 25638
rect 8036 25498 8064 25774
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 8172 25596 8480 25605
rect 8172 25594 8178 25596
rect 8234 25594 8258 25596
rect 8314 25594 8338 25596
rect 8394 25594 8418 25596
rect 8474 25594 8480 25596
rect 8234 25542 8236 25594
rect 8416 25542 8418 25594
rect 8172 25540 8178 25542
rect 8234 25540 8258 25542
rect 8314 25540 8338 25542
rect 8394 25540 8418 25542
rect 8474 25540 8480 25542
rect 8172 25531 8480 25540
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 8864 25362 8892 25638
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 7932 24880 7984 24886
rect 7932 24822 7984 24828
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4540 23322 4568 24074
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5368 23798 5396 24006
rect 5920 23866 5948 24210
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4528 23316 4580 23322
rect 4528 23258 4580 23264
rect 4724 23186 4752 23462
rect 5368 23322 5396 23598
rect 5356 23316 5408 23322
rect 5356 23258 5408 23264
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 5368 22522 5396 23258
rect 5276 22494 5396 22522
rect 5448 22500 5500 22506
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4172 21146 4200 21422
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4816 20466 4844 21830
rect 5184 21690 5212 21898
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2148 19514 2176 19790
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18766 2084 19110
rect 2240 18970 2268 20334
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1872 18086 1900 18566
rect 2056 18290 2084 18702
rect 2792 18358 2820 19790
rect 2884 19514 2912 20198
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2976 18766 3004 19654
rect 3436 19514 3464 19790
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18970 3372 19110
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 3528 18426 3556 19790
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3712 18426 3740 18566
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 2056 16046 2084 18226
rect 3804 17882 3832 18634
rect 3896 18426 3924 19382
rect 3988 18766 4016 19654
rect 4540 19514 4568 19654
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 18834 4108 19314
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18902 4200 19246
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 4540 18834 4568 19450
rect 5276 19174 5304 22494
rect 5448 22442 5500 22448
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5368 21622 5396 22374
rect 5460 22234 5488 22442
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5552 21894 5580 23802
rect 6104 23526 6132 24210
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7484 24154 7512 24210
rect 8036 24154 8064 25298
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 8576 25220 8628 25226
rect 8576 25162 8628 25168
rect 8172 24508 8480 24517
rect 8172 24506 8178 24508
rect 8234 24506 8258 24508
rect 8314 24506 8338 24508
rect 8394 24506 8418 24508
rect 8474 24506 8480 24508
rect 8234 24454 8236 24506
rect 8416 24454 8418 24506
rect 8172 24452 8178 24454
rect 8234 24452 8258 24454
rect 8314 24452 8338 24454
rect 8394 24452 8418 24454
rect 8474 24452 8480 24454
rect 8172 24443 8480 24452
rect 8588 24274 8616 25162
rect 9508 24954 9536 25230
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 10428 24886 10456 25638
rect 10980 25498 11008 25774
rect 12440 25764 12492 25770
rect 12440 25706 12492 25712
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 12452 25650 12480 25706
rect 12900 25696 12952 25702
rect 12452 25622 12572 25650
rect 12900 25638 12952 25644
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 11440 24954 11468 25230
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 6092 23520 6144 23526
rect 6932 23508 6960 24142
rect 7024 23866 7052 24142
rect 7484 24126 7696 24154
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7012 23520 7064 23526
rect 6932 23480 7012 23508
rect 6092 23462 6144 23468
rect 7012 23462 7064 23468
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 5920 22234 5948 22510
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 6932 22166 6960 22374
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 20942 5948 21286
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5552 20602 5580 20810
rect 6012 20806 6040 21830
rect 6472 21690 6500 21966
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 7024 21486 7052 23462
rect 7484 22094 7512 24126
rect 7668 24070 7696 24126
rect 7944 24126 8064 24154
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7576 22778 7604 24006
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7392 22066 7512 22094
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7208 21554 7236 21898
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7300 21554 7328 21830
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 21146 7328 21286
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7196 20868 7248 20874
rect 7196 20810 7248 20816
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 7208 20602 7236 20810
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6288 19514 6316 19722
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 4080 18426 4108 18770
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4448 18290 4476 18770
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4724 18630 4752 18702
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 16250 3004 16390
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2056 15502 2084 15982
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15162 2176 15370
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2700 15094 2728 15438
rect 3436 15094 3464 16934
rect 3988 16250 4016 17070
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16250 4200 16594
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15570 4108 15846
rect 4172 15706 4200 16050
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2792 14618 2820 14894
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 4264 14482 4292 18090
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4356 17746 4384 18022
rect 4724 17882 4752 18022
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4724 17338 4752 17818
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4356 16046 4384 17274
rect 5276 17066 5304 19110
rect 5368 18834 5396 19110
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4724 16658 4752 17002
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4448 15366 4476 16186
rect 4632 16046 4660 16526
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4908 15570 4936 16458
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4356 15026 4384 15302
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2976 12918 3004 13126
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 12306 3004 12582
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 11898 1624 12038
rect 2976 11898 3004 12106
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 11898 3096 12038
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 2872 11280 2924 11286
rect 2502 11248 2558 11257
rect 2872 11222 2924 11228
rect 2502 11183 2558 11192
rect 2516 11150 2544 11183
rect 2884 11150 2912 11222
rect 3160 11150 3188 11562
rect 2504 11144 2556 11150
rect 2780 11144 2832 11150
rect 2504 11086 2556 11092
rect 2778 11112 2780 11121
rect 2872 11144 2924 11150
rect 2832 11112 2834 11121
rect 2872 11086 2924 11092
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2778 11047 2834 11056
rect 2792 10810 2820 11047
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10810 2912 10950
rect 3252 10826 3280 12174
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3344 11132 3372 12038
rect 3436 11558 3464 12038
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3424 11144 3476 11150
rect 3344 11104 3424 11132
rect 3424 11086 3476 11092
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2872 10804 2924 10810
rect 3252 10798 3372 10826
rect 2872 10746 2924 10752
rect 3344 10674 3372 10798
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10198 3096 10474
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 3068 6866 3096 9930
rect 3160 9178 3188 10542
rect 3252 10470 3280 10610
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3344 10266 3372 10610
rect 3436 10266 3464 11086
rect 3528 11014 3556 13262
rect 3896 12238 3924 13262
rect 4264 12434 4292 14418
rect 4448 14346 4476 15302
rect 4816 14822 4844 15438
rect 5092 15162 5120 15982
rect 5368 15586 5396 18770
rect 5552 18222 5580 18906
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5552 17746 5580 18158
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5276 15570 5396 15586
rect 6104 15570 6132 18022
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6288 16794 6316 17546
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6472 15638 6500 19246
rect 6932 18970 6960 19790
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7024 18766 7052 19654
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7116 18290 7144 19110
rect 7208 18358 7236 19110
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17338 6960 17478
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 16794 6776 16934
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 5264 15564 5396 15570
rect 5316 15558 5396 15564
rect 5264 15506 5316 15512
rect 5368 15162 5396 15558
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6104 15366 6132 15506
rect 6564 15502 6592 15846
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6748 15162 6776 15574
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14414 5028 14758
rect 5368 14618 5396 15098
rect 6932 14822 6960 15302
rect 7024 14958 7052 15506
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5552 14346 5580 14758
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 6012 13326 6040 14350
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14074 6960 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6840 13326 6868 13670
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12434 4844 12582
rect 6472 12442 6500 13194
rect 6840 12714 6868 13262
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 4264 12406 4384 12434
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11898 3924 12174
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11898 4292 12106
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 11150 4108 11562
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3804 11014 3832 11086
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3528 10798 3924 10826
rect 3988 10810 4016 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10810 4292 10950
rect 3528 10674 3556 10798
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3896 10690 3924 10798
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3804 10606 3832 10678
rect 3896 10674 4200 10690
rect 3896 10668 4212 10674
rect 3896 10662 4160 10668
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3804 10062 3832 10542
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9722 3372 9862
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3160 8430 3188 8978
rect 3252 8974 3280 9318
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8498 3832 8910
rect 3896 8566 3924 10662
rect 4160 10610 4212 10616
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4172 10418 4200 10610
rect 4080 10062 4108 10406
rect 4172 10390 4292 10418
rect 4264 10130 4292 10390
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4080 9178 4108 9998
rect 4172 9926 4200 9998
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8634 4292 8978
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5914 1900 6190
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1964 5846 1992 6598
rect 2976 5914 3004 6734
rect 3160 6118 3188 8366
rect 3528 8090 3556 8434
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3804 8022 3832 8434
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3712 7546 3740 7822
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3804 7274 3832 7686
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 3160 5778 3188 6054
rect 3252 5846 3280 6734
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 6458 3464 6666
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 6322 3556 6734
rect 3516 6316 3568 6322
rect 3436 6276 3516 6304
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3252 5370 3280 5782
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 1860 5092 1912 5098
rect 1860 5034 1912 5040
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 800 980 3431
rect 1412 2774 1440 4082
rect 1582 4040 1638 4049
rect 1582 3975 1584 3984
rect 1636 3975 1638 3984
rect 1584 3946 1636 3952
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 3194 1808 3402
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1872 2990 1900 5034
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4826 2820 4966
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1412 2746 1532 2774
rect 1504 800 1532 2746
rect 1872 2514 1900 2926
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1964 2446 1992 4422
rect 2792 4214 2820 4422
rect 2780 4208 2832 4214
rect 2240 4146 2360 4162
rect 2780 4150 2832 4156
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2228 4140 2360 4146
rect 2280 4134 2360 4140
rect 2228 4082 2280 4088
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2056 2990 2084 3878
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2148 2446 2176 3334
rect 2240 3194 2268 3878
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2228 2984 2280 2990
rect 2226 2952 2228 2961
rect 2280 2952 2282 2961
rect 2226 2887 2282 2896
rect 2332 2774 2360 4134
rect 2884 2774 2912 4150
rect 2976 3738 3004 5238
rect 3436 5098 3464 6276
rect 3516 6258 3568 6264
rect 3804 5302 3832 7210
rect 4356 6798 4384 12406
rect 4724 12406 4844 12434
rect 6460 12436 6512 12442
rect 4724 11762 4752 12406
rect 6460 12378 6512 12384
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 5092 11694 5120 12038
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4816 11354 4844 11630
rect 6656 11558 6684 12174
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4436 11280 4488 11286
rect 4434 11248 4436 11257
rect 4488 11248 4490 11257
rect 4490 11206 4568 11234
rect 4434 11183 4490 11192
rect 4436 11144 4488 11150
rect 4434 11112 4436 11121
rect 4488 11112 4490 11121
rect 4434 11047 4490 11056
rect 4540 10266 4568 11206
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5276 8498 5304 8842
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 7886 5304 8434
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3896 6254 3924 6666
rect 4264 6458 4292 6734
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 6458 5028 6598
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5370 3924 6190
rect 5276 6186 5304 7822
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6866 5488 7346
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5460 6186 5488 6802
rect 5552 6662 5580 7278
rect 5828 6866 5856 7278
rect 6012 6866 6040 11494
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6380 9926 6408 10134
rect 6472 10062 6500 10406
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6196 9110 6224 9522
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6196 8430 6224 9046
rect 6380 8838 6408 9522
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8498 6408 8774
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7886 6224 8366
rect 6380 7886 6408 8434
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 6866 6132 7686
rect 6380 7546 6408 7822
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4080 5710 4108 6054
rect 4356 5710 4384 6054
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4826 3280 4966
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3436 4622 3464 5034
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3528 4146 3556 5170
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3068 3602 3096 3878
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3344 3534 3372 3878
rect 3528 3534 3556 4082
rect 3804 4010 3832 5238
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4146 4016 5034
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3528 3126 3556 3470
rect 3712 3194 3740 3470
rect 3988 3466 4016 4082
rect 4080 3602 4108 5646
rect 5276 5574 5304 6122
rect 5460 5710 5488 6122
rect 5552 5710 5580 6598
rect 5644 6186 5672 6666
rect 5828 6338 5856 6802
rect 6012 6458 6040 6802
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5828 6322 5948 6338
rect 5828 6316 5960 6322
rect 5828 6310 5908 6316
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4448 4690 4476 5306
rect 4540 5234 4568 5510
rect 5552 5302 5580 5646
rect 5644 5370 5672 6122
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4448 4214 4476 4626
rect 5276 4622 5304 5034
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 4049 4844 4082
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3528 2854 3556 3062
rect 3988 2922 4016 3402
rect 4540 3194 4568 3470
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3194 4752 3334
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2332 2746 2636 2774
rect 2884 2746 3004 2774
rect 2332 2514 2452 2530
rect 2332 2508 2464 2514
rect 2332 2502 2412 2508
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2056 870 2176 898
rect 2056 800 2084 870
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2148 762 2176 870
rect 2332 762 2360 2502
rect 2412 2450 2464 2456
rect 2608 800 2636 2746
rect 2976 2122 3004 2746
rect 2976 2094 3188 2122
rect 3160 800 3188 2094
rect 3712 800 3740 2858
rect 4172 1578 4200 2926
rect 4908 2650 4936 4558
rect 5276 4486 5304 4558
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5000 4078 5028 4422
rect 5368 4146 5396 5034
rect 5828 5030 5856 6310
rect 5908 6258 5960 6264
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5920 5914 5948 6122
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6104 5914 6132 6054
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 5710 6224 6054
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5644 4146 5672 4558
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5736 4078 5764 4490
rect 6012 4282 6040 4558
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6472 4214 6500 9998
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9178 6592 9930
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6564 6730 6592 9114
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3466 5396 3878
rect 6196 3738 6224 4082
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6288 3738 6316 4014
rect 6656 3738 6684 11494
rect 6932 11150 6960 13670
rect 7024 12918 7052 14894
rect 7116 14006 7144 15370
rect 7208 15026 7236 15370
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12306 7052 12582
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10674 6868 10950
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9586 6776 10066
rect 7024 9654 7052 10134
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9042 6776 9522
rect 7116 9450 7144 13806
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6748 8566 6776 8978
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6932 7886 6960 8978
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7116 6798 7144 9386
rect 7208 9110 7236 14418
rect 7300 13870 7328 21082
rect 7392 19922 7420 22066
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7484 20806 7512 21898
rect 7576 21146 7604 22442
rect 7668 21690 7696 22578
rect 7760 22166 7788 22646
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 20398 7512 20742
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7392 19310 7420 19654
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16794 7420 17070
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7392 12782 7420 16730
rect 7484 15450 7512 20334
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7576 19514 7604 19790
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7564 19304 7616 19310
rect 7760 19258 7788 22102
rect 7944 22094 7972 24126
rect 8172 23420 8480 23429
rect 8172 23418 8178 23420
rect 8234 23418 8258 23420
rect 8314 23418 8338 23420
rect 8394 23418 8418 23420
rect 8474 23418 8480 23420
rect 8234 23366 8236 23418
rect 8416 23366 8418 23418
rect 8172 23364 8178 23366
rect 8234 23364 8258 23366
rect 8314 23364 8338 23366
rect 8394 23364 8418 23366
rect 8474 23364 8480 23366
rect 8172 23355 8480 23364
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8588 22574 8616 22918
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8172 22332 8480 22341
rect 8172 22330 8178 22332
rect 8234 22330 8258 22332
rect 8314 22330 8338 22332
rect 8394 22330 8418 22332
rect 8474 22330 8480 22332
rect 8234 22278 8236 22330
rect 8416 22278 8418 22330
rect 8172 22276 8178 22278
rect 8234 22276 8258 22278
rect 8314 22276 8338 22278
rect 8394 22276 8418 22278
rect 8474 22276 8480 22278
rect 8172 22267 8480 22276
rect 8588 22094 8616 22510
rect 7852 22066 7972 22094
rect 8496 22066 8616 22094
rect 7852 20346 7880 22066
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8312 21554 8340 21830
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 20806 7972 21422
rect 8496 21350 8524 22066
rect 8680 22012 8708 24686
rect 9876 24206 9904 24686
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11256 24274 11284 24550
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10704 23866 10732 24074
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 11256 23798 11284 24210
rect 11716 24070 11744 25094
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 11900 24410 11928 24550
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 12360 24138 12388 24550
rect 12452 24206 12480 25230
rect 12544 24750 12572 25622
rect 12912 25294 12940 25638
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24750 12664 25094
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12544 24290 12572 24686
rect 13188 24682 13216 25706
rect 13832 24954 13860 25774
rect 14384 25498 14412 25774
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13820 24948 13872 24954
rect 13820 24890 13872 24896
rect 13924 24834 13952 25094
rect 13740 24806 13952 24834
rect 14292 24818 14320 25434
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14752 24954 14780 25094
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14280 24812 14332 24818
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 12544 24262 12756 24290
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11244 23792 11296 23798
rect 11244 23734 11296 23740
rect 11348 23186 11376 24006
rect 11440 23866 11468 24006
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 12360 23322 12388 24074
rect 12636 23526 12664 24074
rect 12624 23520 12676 23526
rect 12452 23468 12624 23474
rect 12452 23462 12676 23468
rect 12452 23446 12664 23462
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 10600 22568 10652 22574
rect 10600 22510 10652 22516
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8864 22098 8892 22374
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8588 21984 8708 22012
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8036 20874 8064 21286
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7944 20534 7972 20742
rect 7932 20528 7984 20534
rect 7932 20470 7984 20476
rect 7852 20318 7972 20346
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7852 19530 7880 19858
rect 7944 19718 7972 20318
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7852 19502 7972 19530
rect 7564 19246 7616 19252
rect 7576 18766 7604 19246
rect 7668 19230 7788 19258
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7668 19174 7696 19230
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7668 18834 7696 19110
rect 7852 18970 7880 19246
rect 7944 19174 7972 19502
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 17814 7604 18702
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7576 17066 7604 17750
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7668 15570 7696 18770
rect 7944 18086 7972 19110
rect 8036 18850 8064 20810
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 8036 18822 8156 18850
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 8036 18426 8064 18702
rect 8128 18426 8156 18822
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 8588 17882 8616 21984
rect 9140 21554 9168 22442
rect 9416 22234 9444 22510
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9416 21690 9444 21830
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8772 18086 8800 21286
rect 9692 21010 9720 21966
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 18766 9076 20334
rect 9692 20058 9720 20402
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9784 19854 9812 21286
rect 10336 21010 10364 21966
rect 10612 21894 10640 22510
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10704 21962 10732 22374
rect 11348 22234 11376 22510
rect 11900 22234 11928 22510
rect 12268 22234 12296 22646
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12452 22030 12480 23446
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 12544 21894 12572 22374
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10520 20942 10548 21286
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19417 10088 19654
rect 10046 19408 10102 19417
rect 9864 19372 9916 19378
rect 10046 19343 10102 19352
rect 9864 19314 9916 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8760 18080 8812 18086
rect 8680 18040 8760 18068
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 16114 7788 17682
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15706 7880 15982
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7484 15422 7696 15450
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15162 7512 15302
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7380 12776 7432 12782
rect 7300 12724 7380 12730
rect 7300 12718 7432 12724
rect 7300 12702 7420 12718
rect 7300 11830 7328 12702
rect 7484 12434 7512 14962
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7576 14618 7604 14894
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7668 14498 7696 15422
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7576 14470 7696 14498
rect 7576 12442 7604 14470
rect 7852 14414 7880 15098
rect 8128 15094 8156 15302
rect 8496 15094 8524 15642
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8128 14822 8156 15030
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8036 14618 8064 14758
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7760 12986 7788 14350
rect 8036 14090 8064 14418
rect 8036 14062 8156 14090
rect 8680 14074 8708 18040
rect 8760 18022 8812 18028
rect 9048 17746 9076 18702
rect 9416 18698 9444 19110
rect 9692 18970 9720 19246
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9232 18290 9260 18634
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9416 18222 9444 18634
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8772 17338 8800 17478
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 9140 17270 9168 18158
rect 9876 17882 9904 19314
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10152 18290 10180 18906
rect 10244 18766 10272 19110
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9968 17882 9996 18158
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9508 17270 9536 17546
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9876 17082 9904 17818
rect 9968 17270 9996 17818
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9956 17128 10008 17134
rect 9876 17076 9956 17082
rect 9876 17070 10008 17076
rect 9876 17054 9996 17070
rect 9770 16688 9826 16697
rect 9770 16623 9772 16632
rect 9824 16623 9826 16632
rect 9772 16594 9824 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16250 9352 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 15162 9168 15302
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8128 14006 8156 14062
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7392 12406 7512 12434
rect 7564 12436 7616 12442
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7300 11082 7328 11766
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7392 9178 7420 12406
rect 7564 12378 7616 12384
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7484 10810 7512 11698
rect 7576 11354 7604 12038
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7668 9178 7696 12854
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11218 7788 12310
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10810 7788 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7852 9926 7880 13806
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 8772 13258 8800 14486
rect 9140 14482 9168 15098
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9232 14550 9260 14826
rect 9692 14618 9720 15438
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8864 13734 8892 14350
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8864 13394 8892 13670
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12986 8156 13126
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12238 8064 12582
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 9508 12306 9536 13942
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11694 8064 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 9772 12096 9824 12102
rect 9876 12084 9904 14758
rect 9968 12434 9996 17054
rect 10152 13274 10180 17274
rect 10244 17202 10272 18022
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10428 17134 10456 20402
rect 10612 19718 10640 21830
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 12728 21554 12756 24262
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 13004 22094 13032 22918
rect 12820 22066 13032 22094
rect 12820 22030 12848 22066
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21554 13032 21830
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 10704 21146 10732 21286
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 11992 21078 12020 21286
rect 12360 21146 12388 21422
rect 12728 21350 12756 21490
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10612 19310 10640 19654
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10336 16590 10364 16934
rect 10428 16794 10456 17070
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10428 15638 10456 16730
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10428 14958 10456 15574
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10336 14414 10364 14758
rect 10520 14618 10548 14758
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10612 14482 10640 19246
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18426 10732 18566
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10796 16658 10824 20198
rect 10888 19718 10916 20334
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10704 16538 10732 16594
rect 10888 16538 10916 19654
rect 11716 18698 11744 20198
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19378 12572 19790
rect 12820 19446 12848 20742
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 12544 17746 12572 19314
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12544 17270 12572 17682
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12544 16794 12572 17206
rect 12636 17202 12664 18022
rect 13004 17882 13032 18158
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13096 17814 13124 24142
rect 13188 21418 13216 24618
rect 13556 24410 13584 24686
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13556 23866 13584 24346
rect 13648 24070 13676 24686
rect 13740 24206 13768 24806
rect 14280 24754 14332 24760
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13648 23730 13676 24006
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13280 22982 13308 23598
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 13188 20262 13216 21354
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 13280 16538 13308 22918
rect 13556 22778 13584 23054
rect 13648 22778 13676 23666
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13740 23118 13768 23462
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13636 22772 13688 22778
rect 13688 22732 13768 22760
rect 13636 22714 13688 22720
rect 13544 22500 13596 22506
rect 13544 22442 13596 22448
rect 13556 22094 13584 22442
rect 13636 22094 13688 22098
rect 13556 22092 13688 22094
rect 13556 22066 13636 22092
rect 13636 22034 13688 22040
rect 13740 21962 13768 22732
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13464 20602 13492 20878
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13372 19514 13400 19722
rect 13740 19718 13768 21898
rect 13832 21622 13860 24142
rect 14108 23866 14136 24142
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 22234 13952 22510
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13924 21554 13952 22170
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13924 20806 13952 21286
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13372 17066 13400 18158
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 10704 16510 10916 16538
rect 12808 16516 12860 16522
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10336 13870 10364 14350
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 13870 10456 14214
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10152 13246 10272 13274
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9968 12406 10088 12434
rect 9824 12056 9904 12084
rect 9772 12038 9824 12044
rect 8680 11762 8708 12038
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7944 11354 7972 11630
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8036 10606 8064 11630
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8588 10742 8616 11494
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8024 10600 8076 10606
rect 8680 10554 8708 11698
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8024 10542 8076 10548
rect 8036 10266 8064 10542
rect 8588 10526 8708 10554
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7208 8498 7236 9046
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7410 7328 7822
rect 7392 7410 7420 8434
rect 7668 8294 7696 8774
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7576 7546 7604 8026
rect 7668 7750 7696 8230
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 7002 7420 7346
rect 7668 7274 7696 7686
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4758 7052 4966
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7024 3890 7052 4694
rect 7208 4185 7236 5578
rect 7300 5234 7328 6190
rect 7668 5914 7696 6802
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7668 5302 7696 5850
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4622 7420 4966
rect 7760 4826 7788 8842
rect 7852 8634 7880 9522
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 7954 7880 8366
rect 7840 7948 7892 7954
rect 8036 7936 8064 9454
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 8588 9110 8616 10526
rect 8956 10198 8984 11086
rect 9784 10606 9812 12038
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 11354 9996 11630
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9968 10810 9996 11018
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10198 9444 10406
rect 9876 10266 9904 10474
rect 10060 10266 10088 12406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9382 8800 9862
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9678 9480 9734 9489
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8772 8906 8800 9318
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8220 8566 8248 8774
rect 8496 8634 8524 8774
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 8588 8090 8616 8230
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8036 7908 8156 7936
rect 7840 7890 7892 7896
rect 7852 7410 7880 7890
rect 8128 7818 8156 7908
rect 8680 7886 8708 8842
rect 8956 8498 8984 9318
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7410 8156 7754
rect 9232 7410 9260 9046
rect 9416 7546 9444 9454
rect 9678 9415 9734 9424
rect 9692 9382 9720 9415
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9508 7410 9536 8570
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 8772 6798 8800 7278
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4214 7880 4422
rect 7840 4208 7892 4214
rect 7194 4176 7250 4185
rect 7840 4150 7892 4156
rect 7194 4111 7196 4120
rect 7248 4111 7250 4120
rect 7932 4140 7984 4146
rect 7196 4082 7248 4088
rect 7932 4082 7984 4088
rect 7564 3936 7616 3942
rect 7024 3862 7144 3890
rect 7564 3878 7616 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 6196 2446 6224 3674
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 2990 6408 3538
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6368 2984 6420 2990
rect 6366 2952 6368 2961
rect 6420 2952 6422 2961
rect 6748 2922 6776 3470
rect 7116 3058 7144 3862
rect 7576 3466 7604 3878
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7760 3194 7788 3878
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 6366 2887 6422 2896
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 7116 2854 7144 2994
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7668 2650 7696 2994
rect 7852 2854 7880 3878
rect 7944 3074 7972 4082
rect 8036 3194 8064 6666
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 8772 5914 8800 6734
rect 8864 6322 8892 7142
rect 8956 6458 8984 7346
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 9140 5778 9168 6054
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 9140 4826 9168 5170
rect 9232 5098 9260 5646
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8128 4010 8156 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8404 4078 8432 4558
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8116 4004 8168 4010
rect 8107 3952 8116 3992
rect 8107 3946 8168 3952
rect 8107 3720 8135 3946
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 8107 3692 8156 3720
rect 8128 3194 8156 3692
rect 8588 3194 8616 4014
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8680 3398 8708 3946
rect 8772 3466 8800 4082
rect 8852 3528 8904 3534
rect 9140 3482 9168 4490
rect 9218 4176 9274 4185
rect 9218 4111 9220 4120
rect 9272 4111 9274 4120
rect 9220 4082 9272 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 8904 3476 9168 3482
rect 8852 3470 9168 3476
rect 8760 3460 8812 3466
rect 8864 3454 9168 3470
rect 8760 3402 8812 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 7944 3046 8156 3074
rect 8128 2990 8156 3046
rect 8116 2984 8168 2990
rect 8114 2952 8116 2961
rect 8168 2952 8170 2961
rect 8114 2887 8170 2896
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 4172 1550 4292 1578
rect 4264 800 4292 1550
rect 4816 800 4844 2382
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5276 1170 5304 2314
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5276 1142 5396 1170
rect 5368 800 5396 1142
rect 2148 734 2360 762
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6012 762 6040 2246
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 7024 800 7052 2382
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7576 800 7604 2314
rect 8404 1306 8432 2450
rect 8680 2446 8708 3334
rect 9140 3194 9168 3454
rect 9232 3194 9260 3878
rect 9508 3466 9536 3878
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3194 9444 3334
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9692 3126 9720 9318
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 6866 9812 7482
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6322 9812 6802
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9876 5778 9904 8502
rect 9968 7546 9996 10066
rect 10152 9586 10180 13126
rect 10244 12850 10272 13246
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10244 12238 10272 12786
rect 10336 12646 10364 13806
rect 10704 13394 10732 15846
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10336 11694 10364 12582
rect 10796 12442 10824 16510
rect 12808 16458 12860 16464
rect 13188 16510 13308 16538
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10980 14278 11008 14894
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10888 13530 10916 14214
rect 11072 14006 11100 14418
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 12322 10824 12378
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10704 12294 10824 12322
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11150 10364 11630
rect 10520 11218 10548 12242
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10266 10272 11018
rect 10336 10538 10364 11086
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10060 9178 10088 9386
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8634 10088 8910
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10244 8430 10272 9386
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9954 6352 10010 6361
rect 9954 6287 9956 6296
rect 10008 6287 10010 6296
rect 9956 6258 10008 6264
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 4214 9812 5510
rect 9876 5234 9904 5714
rect 9968 5642 9996 6258
rect 10152 5642 10180 6734
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9876 2990 9904 4014
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 3058 9996 3606
rect 10060 3534 10088 5170
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10244 3210 10272 3334
rect 10060 3182 10272 3210
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 8404 1278 8708 1306
rect 8680 800 8708 1278
rect 9232 800 9260 2382
rect 9784 800 9812 2450
rect 10060 2446 10088 3182
rect 10244 3126 10272 3182
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10152 2650 10180 2994
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10244 2650 10272 2926
rect 10336 2922 10364 9998
rect 10428 7886 10456 11018
rect 10612 10810 10640 11494
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10612 10674 10640 10746
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10704 10554 10732 12294
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10612 10526 10732 10554
rect 10612 9674 10640 10526
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10266 10732 10406
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10612 9646 10732 9674
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10520 8430 10548 8842
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 8022 10548 8366
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10520 7834 10548 7958
rect 10520 7806 10640 7834
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7478 10548 7686
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 4622 10548 7142
rect 10612 7002 10640 7806
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10598 6760 10654 6769
rect 10598 6695 10600 6704
rect 10652 6695 10654 6704
rect 10600 6666 10652 6672
rect 10600 6248 10652 6254
rect 10704 6236 10732 9646
rect 10652 6208 10732 6236
rect 10600 6190 10652 6196
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4214 10548 4422
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10506 4040 10562 4049
rect 10506 3975 10562 3984
rect 10520 3466 10548 3975
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3466 10640 3878
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 3194 10640 3402
rect 10796 3210 10824 12174
rect 10888 11558 10916 13126
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11694 11008 12038
rect 11256 11898 11284 14758
rect 11440 12434 11468 16390
rect 12820 16250 12848 16458
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 13188 16114 13216 16510
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16250 13308 16390
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13464 16114 13492 16934
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13188 15638 13216 16050
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 14006 12020 15302
rect 12544 15162 12572 15438
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14890 12480 15030
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 14618 12480 14826
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12268 12986 12296 13670
rect 12360 13326 12388 13874
rect 12452 13530 12480 14282
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 11348 12406 11468 12434
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11348 11762 11376 12406
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10888 10062 10916 11494
rect 10980 11014 11008 11494
rect 11072 11121 11100 11494
rect 11336 11144 11388 11150
rect 11058 11112 11114 11121
rect 11336 11086 11388 11092
rect 11058 11047 11114 11056
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10980 10606 11008 10746
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10888 8430 10916 9658
rect 10980 8634 11008 10406
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7342 10916 8230
rect 10980 7954 11008 8570
rect 11072 8566 11100 9318
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11072 7818 11100 8502
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6730 11008 6802
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 4758 11008 6190
rect 11164 5302 11192 10542
rect 11256 9654 11284 10950
rect 11348 10674 11376 11086
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11440 10606 11468 12106
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11440 9586 11468 9862
rect 11624 9654 11652 11698
rect 12084 11642 12112 11698
rect 11992 11614 12112 11642
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11716 11218 11744 11290
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11716 10062 11744 10678
rect 11900 10130 11928 11086
rect 11992 10130 12020 11614
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10266 12112 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9722 11744 9998
rect 11992 9722 12020 10066
rect 11704 9716 11756 9722
rect 11980 9716 12032 9722
rect 11756 9664 11836 9674
rect 11704 9658 11836 9664
rect 11980 9658 12032 9664
rect 11612 9648 11664 9654
rect 11716 9646 11836 9658
rect 11612 9590 11664 9596
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 7546 11284 8774
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11256 6798 11284 6938
rect 11702 6896 11758 6905
rect 11702 6831 11758 6840
rect 11716 6798 11744 6831
rect 11244 6792 11296 6798
rect 11704 6792 11756 6798
rect 11244 6734 11296 6740
rect 11334 6760 11390 6769
rect 11704 6734 11756 6740
rect 11334 6695 11336 6704
rect 11388 6695 11390 6704
rect 11336 6666 11388 6672
rect 11716 6390 11744 6734
rect 11808 6662 11836 9646
rect 12176 9602 12204 12242
rect 12268 12238 12296 12922
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 9994 12296 12174
rect 12360 11762 12388 13262
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12544 11150 12572 14214
rect 12912 14074 12940 15438
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 15026 13492 15302
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13188 14618 13216 14894
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13464 14278 13492 14962
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13004 13394 13032 14214
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13530 13308 13670
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12728 12102 12756 12922
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 13372 11286 13400 13806
rect 13556 12374 13584 17682
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13648 13190 13676 13942
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12986 13676 13126
rect 13740 12986 13768 19654
rect 13924 18154 13952 20742
rect 14016 20602 14044 21286
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19378 14136 19654
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17678 13860 18022
rect 13924 17882 13952 18090
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 17202 13952 17478
rect 14200 17338 14228 23734
rect 14292 17338 14320 24754
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14844 23050 14872 23462
rect 15120 23118 15148 25842
rect 15752 25356 15804 25362
rect 15752 25298 15804 25304
rect 15394 25052 15702 25061
rect 15394 25050 15400 25052
rect 15456 25050 15480 25052
rect 15536 25050 15560 25052
rect 15616 25050 15640 25052
rect 15696 25050 15702 25052
rect 15456 24998 15458 25050
rect 15638 24998 15640 25050
rect 15394 24996 15400 24998
rect 15456 24996 15480 24998
rect 15536 24996 15560 24998
rect 15616 24996 15640 24998
rect 15696 24996 15702 24998
rect 15394 24987 15702 24996
rect 15764 24818 15792 25298
rect 15856 24818 15884 26250
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 17316 26240 17368 26246
rect 17316 26182 17368 26188
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16500 25362 16528 25978
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 16040 24818 16068 25094
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15394 23964 15702 23973
rect 15394 23962 15400 23964
rect 15456 23962 15480 23964
rect 15536 23962 15560 23964
rect 15616 23962 15640 23964
rect 15696 23962 15702 23964
rect 15456 23910 15458 23962
rect 15638 23910 15640 23962
rect 15394 23908 15400 23910
rect 15456 23908 15480 23910
rect 15536 23908 15560 23910
rect 15616 23908 15640 23910
rect 15696 23908 15702 23910
rect 15394 23899 15702 23908
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14752 22234 14780 22510
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14752 22098 14780 22170
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 19854 14504 21422
rect 15120 20466 15148 23054
rect 15212 22778 15240 23598
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15394 22876 15702 22885
rect 15394 22874 15400 22876
rect 15456 22874 15480 22876
rect 15536 22874 15560 22876
rect 15616 22874 15640 22876
rect 15696 22874 15702 22876
rect 15456 22822 15458 22874
rect 15638 22822 15640 22874
rect 15394 22820 15400 22822
rect 15456 22820 15480 22822
rect 15536 22820 15560 22822
rect 15616 22820 15640 22822
rect 15696 22820 15702 22822
rect 15394 22811 15702 22820
rect 15856 22778 15884 23462
rect 16132 22778 16160 25230
rect 16592 24818 16620 25638
rect 16776 25362 16804 26182
rect 17328 25838 17356 26182
rect 17316 25832 17368 25838
rect 17316 25774 17368 25780
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17592 25832 17644 25838
rect 17592 25774 17644 25780
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16224 23526 16252 24618
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15580 22030 15608 22510
rect 15856 22098 15884 22714
rect 16132 22642 16160 22714
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 15844 22092 15896 22098
rect 16132 22094 16160 22578
rect 15844 22034 15896 22040
rect 15948 22066 16160 22094
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15394 21788 15702 21797
rect 15394 21786 15400 21788
rect 15456 21786 15480 21788
rect 15536 21786 15560 21788
rect 15616 21786 15640 21788
rect 15696 21786 15702 21788
rect 15456 21734 15458 21786
rect 15638 21734 15640 21786
rect 15394 21732 15400 21734
rect 15456 21732 15480 21734
rect 15536 21732 15560 21734
rect 15616 21732 15640 21734
rect 15696 21732 15702 21734
rect 15394 21723 15702 21732
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15304 20602 15332 21286
rect 15844 20800 15896 20806
rect 15948 20788 15976 22066
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 21146 16160 21422
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15896 20760 15976 20788
rect 15844 20742 15896 20748
rect 15394 20700 15702 20709
rect 15394 20698 15400 20700
rect 15456 20698 15480 20700
rect 15536 20698 15560 20700
rect 15616 20698 15640 20700
rect 15696 20698 15702 20700
rect 15456 20646 15458 20698
rect 15638 20646 15640 20698
rect 15394 20644 15400 20646
rect 15456 20644 15480 20646
rect 15536 20644 15560 20646
rect 15616 20644 15640 20646
rect 15696 20644 15702 20646
rect 15394 20635 15702 20644
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14568 19174 14596 20334
rect 14660 19922 14688 20402
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13832 16250 13860 17138
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13924 15162 13952 17138
rect 14292 17134 14320 17274
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 15162 14136 16594
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14482 13860 14758
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13924 14414 13952 15098
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 12986 13860 13874
rect 13924 13258 13952 14350
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13648 12434 13676 12922
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13924 12442 13952 12650
rect 13912 12436 13964 12442
rect 13648 12406 13860 12434
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13832 12322 13860 12406
rect 13912 12378 13964 12384
rect 13832 12294 13952 12322
rect 14108 12306 14136 15098
rect 14292 12434 14320 17070
rect 14464 16040 14516 16046
rect 14384 16000 14464 16028
rect 14384 14770 14412 16000
rect 14464 15982 14516 15988
rect 14384 14742 14504 14770
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12918 14412 13126
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14200 12406 14320 12434
rect 13924 12238 13952 12294
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12544 10470 12572 11086
rect 13556 10674 13584 11154
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 11992 9574 12204 9602
rect 12912 9586 12940 10406
rect 13188 10266 13216 10406
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13556 9722 13584 10610
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13740 9654 13768 11698
rect 13924 11558 13952 12038
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13832 10130 13860 11494
rect 13924 11354 13952 11494
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 12900 9580 12952 9586
rect 11992 7886 12020 9574
rect 12900 9522 12952 9528
rect 13832 9382 13860 9862
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9042 13860 9318
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 12360 8634 12388 8978
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11992 6458 12020 7822
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12084 6458 12112 7278
rect 12176 6866 12204 7278
rect 12268 7002 12296 7822
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 6730 12204 6802
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11164 4826 11192 5238
rect 11256 5234 11284 5510
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11716 4826 11744 6326
rect 12268 5370 12296 6938
rect 12360 6186 12388 8570
rect 12452 7342 12480 8842
rect 14200 8566 14228 12406
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14292 11540 14320 12174
rect 14372 11552 14424 11558
rect 14292 11512 14372 11540
rect 14372 11494 14424 11500
rect 14384 11014 14412 11494
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10742 14412 10950
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14384 9178 14412 9522
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14292 8634 14320 8978
rect 14476 8906 14504 14742
rect 14568 14634 14596 19110
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14648 15156 14700 15162
rect 14700 15116 14780 15144
rect 14648 15098 14700 15104
rect 14568 14606 14688 14634
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14568 11558 14596 12650
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 9994 14596 10950
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12544 7478 12572 7890
rect 12820 7478 12848 8434
rect 13280 8090 13308 8434
rect 14200 8430 14228 8502
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14476 8362 14504 8842
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13832 7954 13860 8298
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7546 13032 7686
rect 14016 7546 14044 7822
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6458 13032 6598
rect 13372 6458 13400 6734
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12452 5914 12480 6258
rect 12912 6225 12940 6258
rect 12898 6216 12954 6225
rect 12898 6151 12954 6160
rect 13556 5914 13584 7278
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12452 5234 12480 5850
rect 13924 5710 13952 6598
rect 14016 6118 14044 6598
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10980 4554 11008 4694
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 4282 11008 4490
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11072 3738 11100 4014
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 10796 3194 10916 3210
rect 10600 3188 10652 3194
rect 10796 3188 10928 3194
rect 10796 3182 10876 3188
rect 10600 3130 10652 3136
rect 10876 3130 10928 3136
rect 10704 3058 10916 3074
rect 12084 3058 12112 3334
rect 10692 3052 10916 3058
rect 10744 3046 10916 3052
rect 10692 2994 10744 3000
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10888 800 10916 3046
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11072 2310 11100 2994
rect 11808 2650 11836 2994
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11520 2440 11572 2446
rect 11440 2400 11520 2428
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11440 800 11468 2400
rect 11520 2382 11572 2388
rect 11992 800 12020 2926
rect 12176 2446 12204 3878
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 2774 12296 3334
rect 12268 2746 12388 2774
rect 12360 2650 12388 2746
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12452 2446 12480 4218
rect 12544 3534 12572 5646
rect 14016 5574 14044 6054
rect 14108 5642 14136 6598
rect 14200 6254 14228 7822
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6458 14320 7142
rect 14568 6866 14596 7482
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14384 6254 14412 6734
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14200 5778 14228 6190
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13464 4146 13492 4762
rect 14016 4644 14228 4672
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 13372 3466 13400 3946
rect 13464 3738 13492 4082
rect 13556 3738 13584 4150
rect 13740 4078 13768 4558
rect 14016 4554 14044 4644
rect 14200 4554 14228 4644
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14108 4146 14136 4490
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4214 14320 4422
rect 14660 4282 14688 14606
rect 14752 14414 14780 15116
rect 14844 15026 14872 17818
rect 14936 17082 14964 18022
rect 15028 17270 15056 18022
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 14936 17054 15056 17082
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14936 16250 14964 16594
rect 15028 16590 15056 17054
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15120 16250 15148 18158
rect 15212 17882 15240 19314
rect 15304 18834 15332 20198
rect 15394 19612 15702 19621
rect 15394 19610 15400 19612
rect 15456 19610 15480 19612
rect 15536 19610 15560 19612
rect 15616 19610 15640 19612
rect 15696 19610 15702 19612
rect 15456 19558 15458 19610
rect 15638 19558 15640 19610
rect 15394 19556 15400 19558
rect 15456 19556 15480 19558
rect 15536 19556 15560 19558
rect 15616 19556 15640 19558
rect 15696 19556 15702 19558
rect 15394 19547 15702 19556
rect 15856 19378 15884 20742
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15672 18970 15700 19314
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15394 18524 15702 18533
rect 15394 18522 15400 18524
rect 15456 18522 15480 18524
rect 15536 18522 15560 18524
rect 15616 18522 15640 18524
rect 15696 18522 15702 18524
rect 15456 18470 15458 18522
rect 15638 18470 15640 18522
rect 15394 18468 15400 18470
rect 15456 18468 15480 18470
rect 15536 18468 15560 18470
rect 15616 18468 15640 18470
rect 15696 18468 15702 18470
rect 15394 18459 15702 18468
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15764 17678 15792 18158
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15394 17436 15702 17445
rect 15394 17434 15400 17436
rect 15456 17434 15480 17436
rect 15536 17434 15560 17436
rect 15616 17434 15640 17436
rect 15696 17434 15702 17436
rect 15456 17382 15458 17434
rect 15638 17382 15640 17434
rect 15394 17380 15400 17382
rect 15456 17380 15480 17382
rect 15536 17380 15560 17382
rect 15616 17380 15640 17382
rect 15696 17380 15702 17382
rect 15394 17371 15702 17380
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14936 14890 14964 15846
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14844 14278 14872 14350
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14832 14068 14884 14074
rect 14936 14056 14964 14826
rect 14884 14028 14964 14056
rect 14832 14010 14884 14016
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14752 12238 14780 12582
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 10470 14780 11494
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14752 5302 14780 6054
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13096 800 13124 3062
rect 13556 2446 13584 3674
rect 14200 3126 14228 4082
rect 14292 3602 14320 4150
rect 14752 4128 14780 4218
rect 14660 4100 14780 4128
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3738 14412 3878
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3194 14412 3470
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14568 3058 14596 3402
rect 14660 3126 14688 4100
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14752 3534 14780 3946
rect 14844 3670 14872 12718
rect 14936 11626 14964 13330
rect 15028 12918 15056 15302
rect 15212 15026 15240 16390
rect 15304 15910 15332 16594
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15856 16538 15884 19314
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 16658 15976 17070
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16794 16068 16934
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15394 16348 15702 16357
rect 15394 16346 15400 16348
rect 15456 16346 15480 16348
rect 15536 16346 15560 16348
rect 15616 16346 15640 16348
rect 15696 16346 15702 16348
rect 15456 16294 15458 16346
rect 15638 16294 15640 16346
rect 15394 16292 15400 16294
rect 15456 16292 15480 16294
rect 15536 16292 15560 16294
rect 15616 16292 15640 16294
rect 15696 16292 15702 16294
rect 15394 16283 15702 16292
rect 15764 16250 15792 16526
rect 15856 16510 15976 16538
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15394 15260 15702 15269
rect 15394 15258 15400 15260
rect 15456 15258 15480 15260
rect 15536 15258 15560 15260
rect 15616 15258 15640 15260
rect 15696 15258 15702 15260
rect 15456 15206 15458 15258
rect 15638 15206 15640 15258
rect 15394 15204 15400 15206
rect 15456 15204 15480 15206
rect 15536 15204 15560 15206
rect 15616 15204 15640 15206
rect 15696 15204 15702 15206
rect 15394 15195 15702 15204
rect 15764 15042 15792 15438
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15672 15014 15792 15042
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15212 14550 15240 14826
rect 15304 14618 15332 14962
rect 15672 14890 15700 15014
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15394 14172 15702 14181
rect 15394 14170 15400 14172
rect 15456 14170 15480 14172
rect 15536 14170 15560 14172
rect 15616 14170 15640 14172
rect 15696 14170 15702 14172
rect 15456 14118 15458 14170
rect 15638 14118 15640 14170
rect 15394 14116 15400 14118
rect 15456 14116 15480 14118
rect 15536 14116 15560 14118
rect 15616 14116 15640 14118
rect 15696 14116 15702 14118
rect 15394 14107 15702 14116
rect 15764 14074 15792 14894
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15856 14414 15884 14758
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15120 13258 15148 13874
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15212 12918 15240 13874
rect 15856 13326 15884 14350
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15394 13084 15702 13093
rect 15394 13082 15400 13084
rect 15456 13082 15480 13084
rect 15536 13082 15560 13084
rect 15616 13082 15640 13084
rect 15696 13082 15702 13084
rect 15456 13030 15458 13082
rect 15638 13030 15640 13082
rect 15394 13028 15400 13030
rect 15456 13028 15480 13030
rect 15536 13028 15560 13030
rect 15616 13028 15640 13030
rect 15696 13028 15702 13030
rect 15394 13019 15702 13028
rect 15764 12918 15792 13126
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 15212 11286 15240 12718
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15394 11996 15702 12005
rect 15394 11994 15400 11996
rect 15456 11994 15480 11996
rect 15536 11994 15560 11996
rect 15616 11994 15640 11996
rect 15696 11994 15702 11996
rect 15456 11942 15458 11994
rect 15638 11942 15640 11994
rect 15394 11940 15400 11942
rect 15456 11940 15480 11942
rect 15536 11940 15560 11942
rect 15616 11940 15640 11942
rect 15696 11940 15702 11942
rect 15394 11931 15702 11940
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10810 15240 11086
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15016 10668 15068 10674
rect 15304 10656 15332 10950
rect 15394 10908 15702 10917
rect 15394 10906 15400 10908
rect 15456 10906 15480 10908
rect 15536 10906 15560 10908
rect 15616 10906 15640 10908
rect 15696 10906 15702 10908
rect 15456 10854 15458 10906
rect 15638 10854 15640 10906
rect 15394 10852 15400 10854
rect 15456 10852 15480 10854
rect 15536 10852 15560 10854
rect 15616 10852 15640 10854
rect 15696 10852 15702 10854
rect 15394 10843 15702 10852
rect 15764 10690 15792 12106
rect 15068 10628 15332 10656
rect 15580 10662 15792 10690
rect 15856 10690 15884 13126
rect 15948 12442 15976 16510
rect 16132 16250 16160 17138
rect 16224 16998 16252 23462
rect 16408 23322 16436 23598
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16868 23050 16896 23462
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 17132 22500 17184 22506
rect 17052 22460 17132 22488
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16120 16244 16172 16250
rect 16040 16204 16120 16232
rect 16040 13394 16068 16204
rect 16120 16186 16172 16192
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 13190 16068 13330
rect 16132 13326 16160 14418
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 16316 12186 16344 21830
rect 16408 20534 16436 22170
rect 16580 22024 16632 22030
rect 16632 21984 16712 22012
rect 16580 21966 16632 21972
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 20602 16620 20878
rect 16684 20602 16712 21984
rect 17052 21418 17080 22460
rect 17132 22442 17184 22448
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17144 22098 17172 22170
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 17236 21146 17264 21966
rect 17328 21894 17356 25774
rect 17420 25226 17448 25774
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17420 24954 17448 25162
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 22778 17448 23598
rect 17512 22778 17540 25638
rect 17604 25430 17632 25774
rect 17880 25770 17908 26250
rect 18708 25838 18736 26726
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17592 25424 17644 25430
rect 17592 25366 17644 25372
rect 17880 24886 17908 25706
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 17972 23866 18000 25434
rect 18236 25220 18288 25226
rect 18236 25162 18288 25168
rect 18248 24954 18276 25162
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18616 24818 18644 25638
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18708 23730 18736 25774
rect 18984 25770 19012 26726
rect 22616 26684 22924 26693
rect 22616 26682 22622 26684
rect 22678 26682 22702 26684
rect 22758 26682 22782 26684
rect 22838 26682 22862 26684
rect 22918 26682 22924 26684
rect 22678 26630 22680 26682
rect 22860 26630 22862 26682
rect 22616 26628 22622 26630
rect 22678 26628 22702 26630
rect 22758 26628 22782 26630
rect 22838 26628 22862 26630
rect 22918 26628 22924 26630
rect 22616 26619 22924 26628
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19812 26042 19840 26318
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 19800 26036 19852 26042
rect 19800 25978 19852 25984
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 19260 25498 19288 25774
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18800 23662 18828 25230
rect 19800 24880 19852 24886
rect 19800 24822 19852 24828
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 23866 19380 24754
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23866 19472 24006
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18800 23186 18828 23598
rect 19352 23322 19380 23802
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17500 22636 17552 22642
rect 17604 22624 17632 22918
rect 18800 22642 18828 23122
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19076 22710 19104 22918
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 17552 22596 17632 22624
rect 17500 22578 17552 22584
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16960 20058 16988 20334
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17134 16436 18022
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16500 12434 16528 18566
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16040 12158 16344 12186
rect 16408 12406 16528 12434
rect 15856 10662 15976 10690
rect 15016 10610 15068 10616
rect 15212 9722 15240 10628
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15304 9602 15332 10134
rect 15580 9908 15608 10662
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15764 10146 15792 10542
rect 15856 10266 15884 10542
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15764 10118 15884 10146
rect 15580 9880 15792 9908
rect 15394 9820 15702 9829
rect 15394 9818 15400 9820
rect 15456 9818 15480 9820
rect 15536 9818 15560 9820
rect 15616 9818 15640 9820
rect 15696 9818 15702 9820
rect 15456 9766 15458 9818
rect 15638 9766 15640 9818
rect 15394 9764 15400 9766
rect 15456 9764 15480 9766
rect 15536 9764 15560 9766
rect 15616 9764 15640 9766
rect 15696 9764 15702 9766
rect 15394 9755 15702 9764
rect 15764 9674 15792 9880
rect 15212 9574 15332 9602
rect 15580 9646 15792 9674
rect 15212 7886 15240 9574
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9178 15332 9318
rect 15488 9178 15516 9386
rect 15580 9382 15608 9646
rect 15856 9602 15884 10118
rect 15672 9574 15884 9602
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15672 8956 15700 9574
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15304 8928 15700 8956
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 7546 15056 7754
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15212 7002 15240 7822
rect 15304 7528 15332 8928
rect 15394 8732 15702 8741
rect 15394 8730 15400 8732
rect 15456 8730 15480 8732
rect 15536 8730 15560 8732
rect 15616 8730 15640 8732
rect 15696 8730 15702 8732
rect 15456 8678 15458 8730
rect 15638 8678 15640 8730
rect 15394 8676 15400 8678
rect 15456 8676 15480 8678
rect 15536 8676 15560 8678
rect 15616 8676 15640 8678
rect 15696 8676 15702 8678
rect 15394 8667 15702 8676
rect 15764 8514 15792 9318
rect 15856 8634 15884 9454
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15764 8486 15884 8514
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15488 7954 15516 8366
rect 15764 8090 15792 8366
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15394 7644 15702 7653
rect 15394 7642 15400 7644
rect 15456 7642 15480 7644
rect 15536 7642 15560 7644
rect 15616 7642 15640 7644
rect 15696 7642 15702 7644
rect 15456 7590 15458 7642
rect 15638 7590 15640 7642
rect 15394 7588 15400 7590
rect 15456 7588 15480 7590
rect 15536 7588 15560 7590
rect 15616 7588 15640 7590
rect 15696 7588 15702 7590
rect 15394 7579 15702 7588
rect 15764 7546 15792 7686
rect 15752 7540 15804 7546
rect 15304 7500 15516 7528
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15212 5302 15240 6258
rect 15304 5914 15332 7278
rect 15396 7002 15424 7346
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15488 6866 15516 7500
rect 15752 7482 15804 7488
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15394 6556 15702 6565
rect 15394 6554 15400 6556
rect 15456 6554 15480 6556
rect 15536 6554 15560 6556
rect 15616 6554 15640 6556
rect 15696 6554 15702 6556
rect 15456 6502 15458 6554
rect 15638 6502 15640 6554
rect 15394 6500 15400 6502
rect 15456 6500 15480 6502
rect 15536 6500 15560 6502
rect 15616 6500 15640 6502
rect 15696 6500 15702 6502
rect 15394 6491 15702 6500
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15856 5658 15884 8486
rect 15948 7546 15976 10662
rect 16040 10198 16068 12158
rect 16408 12102 16436 12406
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16040 7954 16068 9658
rect 16132 8498 16160 12038
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16224 8634 16252 11222
rect 16316 8906 16344 11698
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16040 6390 16068 7890
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16040 5710 16068 6326
rect 16132 5914 16160 6802
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15304 5630 15884 5658
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 5636 15988 5642
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4486 14964 4966
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14936 4146 14964 4422
rect 15120 4146 15148 4422
rect 15212 4214 15240 4762
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15304 3670 15332 5630
rect 15936 5578 15988 5584
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15394 5468 15702 5477
rect 15394 5466 15400 5468
rect 15456 5466 15480 5468
rect 15536 5466 15560 5468
rect 15616 5466 15640 5468
rect 15696 5466 15702 5468
rect 15456 5414 15458 5466
rect 15638 5414 15640 5466
rect 15394 5412 15400 5414
rect 15456 5412 15480 5414
rect 15536 5412 15560 5414
rect 15616 5412 15640 5414
rect 15696 5412 15702 5414
rect 15394 5403 15702 5412
rect 15856 5234 15884 5510
rect 15948 5302 15976 5578
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15394 4380 15702 4389
rect 15394 4378 15400 4380
rect 15456 4378 15480 4380
rect 15536 4378 15560 4380
rect 15616 4378 15640 4380
rect 15696 4378 15702 4380
rect 15456 4326 15458 4378
rect 15638 4326 15640 4378
rect 15394 4324 15400 4326
rect 15456 4324 15480 4326
rect 15536 4324 15560 4326
rect 15616 4324 15640 4326
rect 15696 4324 15702 4326
rect 15394 4315 15702 4324
rect 15384 4140 15436 4146
rect 15436 4100 15792 4128
rect 15384 4082 15436 4088
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13648 800 13676 2926
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14200 800 14228 2450
rect 14476 1578 14504 2994
rect 14844 2650 14872 3470
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15212 2310 15240 3334
rect 15394 3292 15702 3301
rect 15394 3290 15400 3292
rect 15456 3290 15480 3292
rect 15536 3290 15560 3292
rect 15616 3290 15640 3292
rect 15696 3290 15702 3292
rect 15456 3238 15458 3290
rect 15638 3238 15640 3290
rect 15394 3236 15400 3238
rect 15456 3236 15480 3238
rect 15536 3236 15560 3238
rect 15616 3236 15640 3238
rect 15696 3236 15702 3238
rect 15394 3227 15702 3236
rect 15764 3194 15792 4100
rect 16040 4078 16068 4558
rect 16132 4486 16160 5034
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16132 4146 16160 4422
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3398 15976 3878
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15396 2774 15424 3130
rect 16132 3040 16160 4082
rect 16224 3194 16252 8570
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7750 16344 8230
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 6866 16344 7686
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16408 4214 16436 12038
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 9518 16528 11834
rect 16592 10538 16620 16934
rect 16684 15570 16712 19450
rect 17052 19310 17080 19790
rect 17328 19514 17356 20538
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 18970 17080 19246
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17052 18426 17080 18906
rect 17420 18766 17448 22374
rect 17604 22234 17632 22596
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18616 22234 18644 22510
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 19812 22094 19840 24822
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20180 23866 20208 24142
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20272 23866 20300 24074
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19904 23186 19932 23530
rect 20456 23526 20484 25638
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20824 24206 20852 24686
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 20824 23662 20852 24142
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20180 22642 20208 23054
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20180 22234 20208 22578
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20732 22094 20760 22646
rect 20824 22574 20852 23462
rect 20916 22778 20944 24142
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 21284 23730 21312 24006
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21284 23186 21312 23666
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 21192 22234 21220 23122
rect 21272 22636 21324 22642
rect 21376 22624 21404 23462
rect 21468 23118 21496 24006
rect 22112 23798 22140 24006
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21468 22982 21496 23054
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21744 22710 21772 23054
rect 22020 22710 22048 23530
rect 22112 23322 22140 23734
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22204 22778 22232 24142
rect 22480 23186 22508 26250
rect 27620 26240 27672 26246
rect 27620 26182 27672 26188
rect 27632 25906 27660 26182
rect 27816 25974 27844 26726
rect 27804 25968 27856 25974
rect 27804 25910 27856 25916
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 22616 25596 22924 25605
rect 22616 25594 22622 25596
rect 22678 25594 22702 25596
rect 22758 25594 22782 25596
rect 22838 25594 22862 25596
rect 22918 25594 22924 25596
rect 22678 25542 22680 25594
rect 22860 25542 22862 25594
rect 22616 25540 22622 25542
rect 22678 25540 22702 25542
rect 22758 25540 22782 25542
rect 22838 25540 22862 25542
rect 22918 25540 22924 25542
rect 22616 25531 22924 25540
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 22616 24508 22924 24517
rect 22616 24506 22622 24508
rect 22678 24506 22702 24508
rect 22758 24506 22782 24508
rect 22838 24506 22862 24508
rect 22918 24506 22924 24508
rect 22678 24454 22680 24506
rect 22860 24454 22862 24506
rect 22616 24452 22622 24454
rect 22678 24452 22702 24454
rect 22758 24452 22782 24454
rect 22838 24452 22862 24454
rect 22918 24452 22924 24454
rect 22616 24443 22924 24452
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23308 23866 23336 24074
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22616 23420 22924 23429
rect 22616 23418 22622 23420
rect 22678 23418 22702 23420
rect 22758 23418 22782 23420
rect 22838 23418 22862 23420
rect 22918 23418 22924 23420
rect 22678 23366 22680 23418
rect 22860 23366 22862 23418
rect 22616 23364 22622 23366
rect 22678 23364 22702 23366
rect 22758 23364 22782 23366
rect 22838 23364 22862 23366
rect 22918 23364 22924 23366
rect 22616 23355 22924 23364
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 21324 22596 21404 22624
rect 21272 22578 21324 22584
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 19812 22066 19932 22094
rect 19904 21894 19932 22066
rect 20640 22066 20760 22094
rect 20640 21962 20668 22066
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17604 19854 17632 20198
rect 17880 19922 17908 20198
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 18064 19718 18092 20470
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17338 16804 17614
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 14074 16988 14350
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17052 13462 17080 18362
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17328 17270 17356 17682
rect 18064 17610 18092 19654
rect 18248 19514 18276 20334
rect 18616 19922 18644 20946
rect 19076 20058 19104 21422
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20602 19380 20878
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19536 19990 19564 20742
rect 19628 20534 19656 21286
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18616 19174 18644 19858
rect 19536 19854 19564 19926
rect 19720 19922 19748 20198
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19812 19802 19840 21830
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 18788 19780 18840 19786
rect 18972 19780 19024 19786
rect 18840 19740 18972 19768
rect 18788 19722 18840 19728
rect 19812 19774 19932 19802
rect 18972 19722 19024 19728
rect 19904 19718 19932 19774
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17328 16658 17356 17206
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 16250 17356 16594
rect 17696 16590 17724 17478
rect 18064 16998 18092 17546
rect 18248 17338 18276 17614
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 17338 18552 17478
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18616 17218 18644 19110
rect 19260 18970 19288 19314
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19536 18834 19564 19654
rect 19904 19514 19932 19654
rect 19996 19514 20024 20334
rect 20456 20330 20484 21830
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18524 17190 18644 17218
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17052 13258 17080 13398
rect 17236 13274 17264 15302
rect 17328 13394 17356 16186
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17604 15162 17632 16050
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17972 15026 18000 15302
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17420 13326 17448 13670
rect 17408 13320 17460 13326
rect 17040 13252 17092 13258
rect 17236 13246 17356 13274
rect 17408 13262 17460 13268
rect 17040 13194 17092 13200
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 16776 12850 16804 13126
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16776 12442 16804 12786
rect 16764 12436 16816 12442
rect 17236 12434 17264 13126
rect 16764 12378 16816 12384
rect 17052 12406 17264 12434
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 11286 16896 11562
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16960 11082 16988 11494
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16776 10130 16804 10610
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16948 10124 17000 10130
rect 17052 10112 17080 12406
rect 17328 12238 17356 13246
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17604 12442 17632 12786
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10130 17172 10950
rect 17512 10810 17540 11630
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17696 10130 17724 10950
rect 17000 10084 17080 10112
rect 17132 10124 17184 10130
rect 16948 10066 17000 10072
rect 17132 10066 17184 10072
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9722 16620 9998
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16500 8906 16528 9454
rect 16592 9178 16620 9658
rect 16960 9586 16988 10066
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 16684 9178 16712 9318
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 16946 7848 17002 7857
rect 16672 7812 16724 7818
rect 16946 7783 16948 7792
rect 16672 7754 16724 7760
rect 17000 7783 17002 7792
rect 16948 7754 17000 7760
rect 16684 7206 16712 7754
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16500 6458 16528 6734
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16500 4826 16528 5170
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16316 3194 16344 4014
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16212 3052 16264 3058
rect 16132 3012 16212 3040
rect 16212 2994 16264 3000
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15304 2746 15424 2774
rect 15304 2514 15332 2746
rect 16040 2650 16068 2858
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14476 1550 14780 1578
rect 14752 800 14780 1550
rect 15304 800 15332 2314
rect 15394 2204 15702 2213
rect 15394 2202 15400 2204
rect 15456 2202 15480 2204
rect 15536 2202 15560 2204
rect 15616 2202 15640 2204
rect 15696 2202 15702 2204
rect 15456 2150 15458 2202
rect 15638 2150 15640 2202
rect 15394 2148 15400 2150
rect 15456 2148 15480 2150
rect 15536 2148 15560 2150
rect 15616 2148 15640 2150
rect 15696 2148 15702 2150
rect 15394 2139 15702 2148
rect 15856 800 15884 2450
rect 16408 800 16436 4014
rect 16500 3890 16528 4762
rect 16592 4690 16620 4762
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16776 4049 16804 4694
rect 16762 4040 16818 4049
rect 16762 3975 16818 3984
rect 16500 3862 16620 3890
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16500 3194 16528 3674
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 3126 16620 3862
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3126 16712 3334
rect 16960 3194 16988 7346
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6322 17448 7142
rect 17604 6866 17632 8230
rect 17696 7954 17724 9318
rect 17788 8634 17816 14894
rect 18064 14890 18092 16934
rect 18432 16182 18460 17138
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18432 15994 18460 16118
rect 18340 15966 18460 15994
rect 18340 15434 18368 15966
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 18340 14074 18368 15370
rect 18432 15026 18460 15846
rect 18524 15570 18552 17190
rect 18984 16794 19012 17614
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18524 15026 18552 15506
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17880 13190 17908 13670
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17972 12434 18000 13670
rect 18524 13530 18552 14350
rect 18708 14090 18736 14486
rect 18708 14062 18920 14090
rect 18708 13870 18736 14062
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 17972 12406 18092 12434
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10674 18000 10950
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17868 10260 17920 10266
rect 18064 10248 18092 12406
rect 18156 11762 18184 12582
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18340 11558 18368 12038
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 17920 10220 18092 10248
rect 17868 10202 17920 10208
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7206 17724 7890
rect 17972 7886 18000 9862
rect 18064 9382 18092 10220
rect 18156 9654 18184 10406
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18248 9178 18276 9862
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18064 7954 18092 8570
rect 18340 8430 18368 11494
rect 18432 11354 18460 13194
rect 18800 12170 18828 13942
rect 18892 12442 18920 14062
rect 18984 13716 19012 15846
rect 19076 15502 19104 16662
rect 19168 16250 19196 18158
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19536 16114 19564 17206
rect 19628 16454 19656 17478
rect 19812 17202 19840 18022
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16250 19656 16390
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 15162 19104 15438
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19168 13802 19196 15302
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19064 13728 19116 13734
rect 18984 13688 19064 13716
rect 19064 13670 19116 13676
rect 19076 13326 19104 13670
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12850 19104 13126
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18432 10130 18460 11290
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18708 10266 18736 10542
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18432 9178 18460 9318
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18524 7954 18552 9318
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17696 6866 17724 7142
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17604 6322 17632 6802
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5914 17080 6054
rect 17696 5914 17724 6802
rect 18064 6798 18092 7686
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 7002 18276 7346
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18340 6866 18368 7278
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17880 6458 17908 6666
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17696 5302 17724 5510
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 3194 17080 3470
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 17328 3058 17356 3878
rect 17420 3602 17448 5102
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4622 17632 4966
rect 17972 4826 18000 5646
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 18156 4690 18184 4966
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17866 4312 17922 4321
rect 17866 4247 17922 4256
rect 17880 4214 17908 4247
rect 18156 4214 18184 4626
rect 18248 4554 18276 6054
rect 18340 4826 18368 6326
rect 18524 6322 18552 7686
rect 18892 7546 18920 12378
rect 19260 11014 19288 14826
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 14074 19380 14282
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19536 13938 19564 16050
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19628 15366 19656 15982
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19720 14414 19748 16730
rect 19904 16590 19932 19450
rect 20456 19174 20484 20266
rect 20548 19922 20576 20402
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20628 19712 20680 19718
rect 20680 19660 20760 19666
rect 20628 19654 20760 19660
rect 20640 19638 20760 19654
rect 20732 19378 20760 19638
rect 21008 19514 21036 20334
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17338 20300 17614
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20180 16658 20208 17274
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19904 15910 19932 16526
rect 20364 16182 20392 17478
rect 20456 16658 20484 19110
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20732 18154 20760 18362
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 17218 20760 18090
rect 20916 18086 20944 19110
rect 21100 18970 21128 19994
rect 21192 19854 21220 20470
rect 21284 20466 21312 22578
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22204 22030 22232 22442
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21192 19446 21220 19790
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21284 19378 21312 20402
rect 22020 20398 22048 20742
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21468 20058 21496 20266
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21456 19916 21508 19922
rect 21560 19904 21588 20198
rect 21508 19876 21588 19904
rect 21456 19858 21508 19864
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21744 19446 21772 19654
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21836 19394 21864 20198
rect 21836 19378 21956 19394
rect 21272 19372 21324 19378
rect 21836 19372 21968 19378
rect 21836 19366 21916 19372
rect 21272 19314 21324 19320
rect 21916 19314 21968 19320
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20824 17338 20852 17478
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20640 17202 20760 17218
rect 20628 17196 20760 17202
rect 20680 17190 20760 17196
rect 20628 17138 20680 17144
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 20456 15434 20484 16594
rect 20628 16244 20680 16250
rect 20732 16232 20760 17070
rect 20824 16794 20852 17274
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20680 16204 20760 16232
rect 20628 16186 20680 16192
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20916 15366 20944 18022
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17338 21036 17614
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16522 21036 16934
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19720 11898 19748 13874
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19812 11762 19840 14418
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20088 13410 20116 14214
rect 20180 13530 20208 14214
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20088 13382 20208 13410
rect 20180 13326 20208 13382
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19904 13190 19932 13262
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19996 12442 20024 12854
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20088 12238 20116 13262
rect 20364 12434 20392 15302
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14074 20852 14350
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20456 13394 20484 13670
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20364 12406 20484 12434
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19904 11762 19932 12038
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 20088 11694 20116 12174
rect 20180 11694 20208 12242
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20456 11626 20484 12406
rect 20732 12102 20760 13330
rect 20916 12850 20944 13670
rect 21008 12986 21036 16458
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 21100 12730 21128 13262
rect 20824 12702 21128 12730
rect 20824 12306 20852 12702
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12442 21128 12582
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19536 10810 19564 11494
rect 20456 11150 20484 11562
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 18984 9926 19012 10542
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18892 6254 18920 7482
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18984 5302 19012 9862
rect 19444 8090 19472 10542
rect 19812 9654 19840 11018
rect 20364 10810 20392 11086
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20548 10674 20576 10950
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20272 10062 20300 10610
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19904 9110 19932 9930
rect 20272 9178 20300 9998
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 9178 20484 9318
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 20272 8634 20300 9114
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19076 6322 19104 6802
rect 19352 6798 19380 7142
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18432 4690 18460 5238
rect 19352 5234 19380 5510
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 19352 4622 19380 5170
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3738 17632 4082
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18064 3738 18092 4014
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18248 3913 18276 3946
rect 18234 3904 18290 3913
rect 18234 3839 18290 3848
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17144 2650 17172 2994
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17604 2446 17632 3334
rect 17788 2514 17908 2530
rect 17788 2508 17920 2514
rect 17788 2502 17868 2508
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 16960 800 16988 2382
rect 17512 870 17632 898
rect 17512 800 17540 870
rect 6012 734 6408 762
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 17604 762 17632 870
rect 17788 762 17816 2502
rect 17868 2450 17920 2456
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 17604 734 17816 762
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 4490
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 4049 18552 4082
rect 18510 4040 18566 4049
rect 18510 3975 18566 3984
rect 18616 3466 18644 4422
rect 18708 4146 18736 4558
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 3738 18736 3946
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18616 800 18644 2926
rect 18800 2854 18828 4422
rect 18878 4312 18934 4321
rect 18878 4247 18934 4256
rect 18892 4214 18920 4247
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 19444 4146 19472 8026
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7546 20208 7686
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20548 7478 20576 9454
rect 20640 8906 20668 9454
rect 20824 9042 20852 9862
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19628 5914 19656 6258
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 20364 5574 20392 7278
rect 20732 7002 20760 7822
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5914 20576 6054
rect 20732 5914 20760 6122
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19076 3738 19104 4014
rect 19260 3913 19288 4014
rect 19246 3904 19302 3913
rect 19246 3839 19302 3848
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19076 3058 19104 3674
rect 19536 3194 19564 4558
rect 19904 4146 19932 4966
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20088 4146 20116 4490
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19904 3942 19932 4082
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19996 3398 20024 4082
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 19168 800 19196 2926
rect 19996 2514 20024 3334
rect 20088 3194 20116 4082
rect 20456 3466 20484 4490
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20640 2922 20668 4422
rect 20824 3738 20852 7754
rect 20916 4706 20944 12106
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 8090 21036 12038
rect 21192 11762 21220 14214
rect 21284 12646 21312 19314
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 14958 21496 18566
rect 22020 18154 22048 20334
rect 22296 18834 22324 22918
rect 22480 22642 22508 23122
rect 23124 22642 23152 23462
rect 23400 23118 23428 24006
rect 23952 23866 23980 24142
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 24228 23322 24256 24686
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24872 23798 24900 24210
rect 25148 24206 25176 25094
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25228 24676 25280 24682
rect 25228 24618 25280 24624
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 24860 23656 24912 23662
rect 24780 23604 24860 23610
rect 24780 23598 24912 23604
rect 24780 23582 24900 23598
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 24780 23066 24808 23582
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23186 24900 23462
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24780 23038 24900 23066
rect 24400 22976 24452 22982
rect 24400 22918 24452 22924
rect 24412 22642 24440 22918
rect 24872 22778 24900 23038
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 22480 22098 22508 22578
rect 24964 22438 24992 24142
rect 25044 24064 25096 24070
rect 25044 24006 25096 24012
rect 25056 23662 25084 24006
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 25056 22710 25084 23598
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 22616 22332 22924 22341
rect 22616 22330 22622 22332
rect 22678 22330 22702 22332
rect 22758 22330 22782 22332
rect 22838 22330 22862 22332
rect 22918 22330 22924 22332
rect 22678 22278 22680 22330
rect 22860 22278 22862 22330
rect 22616 22276 22622 22278
rect 22678 22276 22702 22278
rect 22758 22276 22782 22278
rect 22838 22276 22862 22278
rect 22918 22276 22924 22278
rect 22616 22267 22924 22276
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24872 21690 24900 21830
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 22616 21244 22924 21253
rect 22616 21242 22622 21244
rect 22678 21242 22702 21244
rect 22758 21242 22782 21244
rect 22838 21242 22862 21244
rect 22918 21242 22924 21244
rect 22678 21190 22680 21242
rect 22860 21190 22862 21242
rect 22616 21188 22622 21190
rect 22678 21188 22702 21190
rect 22758 21188 22782 21190
rect 22838 21188 22862 21190
rect 22918 21188 22924 21190
rect 22616 21179 22924 21188
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22388 19922 22416 20742
rect 22480 20602 22508 20742
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22480 20058 22508 20538
rect 22616 20156 22924 20165
rect 22616 20154 22622 20156
rect 22678 20154 22702 20156
rect 22758 20154 22782 20156
rect 22838 20154 22862 20156
rect 22918 20154 22924 20156
rect 22678 20102 22680 20154
rect 22860 20102 22862 20154
rect 22616 20100 22622 20102
rect 22678 20100 22702 20102
rect 22758 20100 22782 20102
rect 22838 20100 22862 20102
rect 22918 20100 22924 20102
rect 22616 20091 22924 20100
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22388 19514 22416 19858
rect 23032 19514 23060 20878
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23216 19854 23244 20198
rect 23676 20058 23704 20878
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24596 20534 24624 20742
rect 24872 20602 24900 21626
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24584 20528 24636 20534
rect 24584 20470 24636 20476
rect 24872 20262 24900 20538
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23952 19446 23980 20198
rect 24872 20058 24900 20198
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 25056 19786 25084 21830
rect 25148 19802 25176 24142
rect 25240 23866 25268 24618
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25332 23798 25360 24754
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25608 22778 25636 25094
rect 26252 24614 26280 25230
rect 27252 25152 27304 25158
rect 27252 25094 27304 25100
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26528 24410 26556 24754
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 25884 23118 25912 23734
rect 26068 23186 26096 24142
rect 26528 24070 26556 24346
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 27080 23866 27108 24142
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 27264 23526 27292 25094
rect 27632 24818 27660 25842
rect 28368 25498 28396 26862
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28356 25492 28408 25498
rect 28356 25434 28408 25440
rect 27712 25424 27764 25430
rect 27712 25366 27764 25372
rect 27724 24886 27752 25366
rect 27712 24880 27764 24886
rect 27712 24822 27764 24828
rect 28460 24818 28488 26250
rect 28736 25838 28764 26862
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30116 26382 30144 26726
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 30104 26376 30156 26382
rect 30104 26318 30156 26324
rect 29276 26240 29328 26246
rect 29276 26182 29328 26188
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 28724 25832 28776 25838
rect 28724 25774 28776 25780
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27540 23866 27568 24074
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 26792 23316 26844 23322
rect 26792 23258 26844 23264
rect 26056 23180 26108 23186
rect 26056 23122 26108 23128
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25792 22658 25820 23054
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 25976 22778 26004 22918
rect 25964 22772 26016 22778
rect 25964 22714 26016 22720
rect 25700 22630 25820 22658
rect 25700 21690 25728 22630
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22234 25820 22510
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 26344 22166 26372 23122
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26332 22160 26384 22166
rect 26332 22102 26384 22108
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25240 20398 25268 20878
rect 25332 20602 25360 20878
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25412 20528 25464 20534
rect 25412 20470 25464 20476
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25424 19922 25452 20470
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25044 19780 25096 19786
rect 25148 19774 25268 19802
rect 25044 19722 25096 19728
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 22616 19068 22924 19077
rect 22616 19066 22622 19068
rect 22678 19066 22702 19068
rect 22758 19066 22782 19068
rect 22838 19066 22862 19068
rect 22918 19066 22924 19068
rect 22678 19014 22680 19066
rect 22860 19014 22862 19066
rect 22616 19012 22622 19014
rect 22678 19012 22702 19014
rect 22758 19012 22782 19014
rect 22838 19012 22862 19014
rect 22918 19012 22924 19014
rect 22616 19003 22924 19012
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21560 16998 21588 17206
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21652 16250 21680 17614
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 21836 16794 21864 17138
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 22112 16250 22140 17138
rect 22204 16250 22232 18566
rect 22616 17980 22924 17989
rect 22616 17978 22622 17980
rect 22678 17978 22702 17980
rect 22758 17978 22782 17980
rect 22838 17978 22862 17980
rect 22918 17978 22924 17980
rect 22678 17926 22680 17978
rect 22860 17926 22862 17978
rect 22616 17924 22622 17926
rect 22678 17924 22702 17926
rect 22758 17924 22782 17926
rect 22838 17924 22862 17926
rect 22918 17924 22924 17926
rect 22616 17915 22924 17924
rect 23400 17610 23428 19110
rect 24412 18970 24440 19314
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24964 18834 24992 19654
rect 25148 19378 25176 19654
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 25240 18698 25268 19774
rect 25424 19174 25452 19858
rect 25792 19514 25820 20878
rect 25976 20398 26004 21286
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 26068 20466 26096 20742
rect 26436 20618 26464 22578
rect 26804 22094 26832 23258
rect 27540 23186 27568 23802
rect 27528 23180 27580 23186
rect 27448 23140 27528 23168
rect 27448 22778 27476 23140
rect 27528 23122 27580 23128
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27540 22642 27568 22918
rect 27632 22642 27660 24754
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 23322 27752 23598
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27816 23118 27844 24006
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 27908 22778 27936 22918
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26712 22066 26832 22094
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26344 20602 26464 20618
rect 26332 20596 26464 20602
rect 26384 20590 26464 20596
rect 26332 20538 26384 20544
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 26068 19922 26096 20402
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26160 19802 26188 20198
rect 26240 19848 26292 19854
rect 26160 19796 26240 19802
rect 26160 19790 26292 19796
rect 26160 19774 26280 19790
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 26344 19378 26372 20538
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26436 20058 26464 20402
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26528 19922 26556 20742
rect 26712 20602 26740 22066
rect 26988 21026 27016 22102
rect 27632 22094 27660 22578
rect 28000 22438 28028 24686
rect 28080 23520 28132 23526
rect 28080 23462 28132 23468
rect 28092 23186 28120 23462
rect 28080 23180 28132 23186
rect 28080 23122 28132 23128
rect 27988 22432 28040 22438
rect 27988 22374 28040 22380
rect 27804 22094 27856 22098
rect 27632 22092 27856 22094
rect 27632 22066 27804 22092
rect 27804 22034 27856 22040
rect 26804 20998 27016 21026
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26528 19718 26556 19858
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25976 18086 26004 18634
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25240 17882 25268 18022
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 23400 17134 23428 17546
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 22616 16892 22924 16901
rect 22616 16890 22622 16892
rect 22678 16890 22702 16892
rect 22758 16890 22782 16892
rect 22838 16890 22862 16892
rect 22918 16890 22924 16892
rect 22678 16838 22680 16890
rect 22860 16838 22862 16890
rect 22616 16836 22622 16838
rect 22678 16836 22702 16838
rect 22758 16836 22782 16838
rect 22838 16836 22862 16838
rect 22918 16836 22924 16838
rect 22616 16827 22924 16836
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22572 16046 22600 16730
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23400 16250 23428 16390
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 22284 16040 22336 16046
rect 22560 16040 22612 16046
rect 22284 15982 22336 15988
rect 22480 16000 22560 16028
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21468 14414 21496 14894
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13326 21404 14214
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21468 13530 21496 13806
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21468 12986 21496 13194
rect 21928 13190 21956 13738
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21560 12442 21588 13126
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21192 9382 21220 11086
rect 21284 10470 21312 11494
rect 21468 11286 21496 12310
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 10810 21496 11086
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21468 10266 21496 10542
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21560 9518 21588 10950
rect 21928 9674 21956 13126
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22112 12306 22140 12922
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22296 11234 22324 15982
rect 22480 15570 22508 16000
rect 22560 15982 22612 15988
rect 22616 15804 22924 15813
rect 22616 15802 22622 15804
rect 22678 15802 22702 15804
rect 22758 15802 22782 15804
rect 22838 15802 22862 15804
rect 22918 15802 22924 15804
rect 22678 15750 22680 15802
rect 22860 15750 22862 15802
rect 22616 15748 22622 15750
rect 22678 15748 22702 15750
rect 22758 15748 22782 15750
rect 22838 15748 22862 15750
rect 22918 15748 22924 15750
rect 22616 15739 22924 15748
rect 22468 15564 22520 15570
rect 22388 15524 22468 15552
rect 22388 13394 22416 15524
rect 22468 15506 22520 15512
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 22616 14716 22924 14725
rect 22616 14714 22622 14716
rect 22678 14714 22702 14716
rect 22758 14714 22782 14716
rect 22838 14714 22862 14716
rect 22918 14714 22924 14716
rect 22678 14662 22680 14714
rect 22860 14662 22862 14714
rect 22616 14660 22622 14662
rect 22678 14660 22702 14662
rect 22758 14660 22782 14662
rect 22838 14660 22862 14662
rect 22918 14660 22924 14662
rect 22616 14651 22924 14660
rect 23216 14618 23244 15370
rect 23860 15094 23888 17274
rect 24780 17134 24808 17274
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 16590 23980 16934
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 24412 16250 24440 17070
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24780 16046 24808 16390
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23400 14618 23428 14758
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 22928 14544 22980 14550
rect 22928 14486 22980 14492
rect 22940 14278 22968 14486
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 23584 14006 23612 14554
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22480 13462 22508 13670
rect 22616 13628 22924 13637
rect 22616 13626 22622 13628
rect 22678 13626 22702 13628
rect 22758 13626 22782 13628
rect 22838 13626 22862 13628
rect 22918 13626 22924 13628
rect 22678 13574 22680 13626
rect 22860 13574 22862 13626
rect 22616 13572 22622 13574
rect 22678 13572 22702 13574
rect 22758 13572 22782 13574
rect 22838 13572 22862 13574
rect 22918 13572 22924 13574
rect 22616 13563 22924 13572
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 12850 22416 13330
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22616 12540 22924 12549
rect 22616 12538 22622 12540
rect 22678 12538 22702 12540
rect 22758 12538 22782 12540
rect 22838 12538 22862 12540
rect 22918 12538 22924 12540
rect 22678 12486 22680 12538
rect 22860 12486 22862 12538
rect 22616 12484 22622 12486
rect 22678 12484 22702 12486
rect 22758 12484 22782 12486
rect 22838 12484 22862 12486
rect 22918 12484 22924 12486
rect 22616 12475 22924 12484
rect 23032 12442 23060 12786
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23400 12102 23428 12378
rect 23478 12200 23534 12209
rect 23478 12135 23534 12144
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 22616 11452 22924 11461
rect 22616 11450 22622 11452
rect 22678 11450 22702 11452
rect 22758 11450 22782 11452
rect 22838 11450 22862 11452
rect 22918 11450 22924 11452
rect 22678 11398 22680 11450
rect 22860 11398 22862 11450
rect 22616 11396 22622 11398
rect 22678 11396 22702 11398
rect 22758 11396 22782 11398
rect 22838 11396 22862 11398
rect 22918 11396 22924 11398
rect 22616 11387 22924 11396
rect 22112 11206 22324 11234
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10169 22048 10950
rect 22112 10470 22140 11206
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22006 10160 22062 10169
rect 22006 10095 22062 10104
rect 21836 9646 21956 9674
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 7002 21036 7142
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21008 6458 21036 6598
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21192 6254 21220 8366
rect 21284 7410 21312 9386
rect 21560 8634 21588 9454
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21652 7002 21680 9318
rect 21836 8294 21864 9646
rect 22020 9586 22048 10095
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22112 8922 22140 10406
rect 22204 9654 22232 11086
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22296 9722 22324 9998
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22204 9058 22232 9386
rect 22296 9178 22324 9658
rect 22388 9178 22416 11222
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22940 10674 22968 10950
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22616 10364 22924 10373
rect 22616 10362 22622 10364
rect 22678 10362 22702 10364
rect 22758 10362 22782 10364
rect 22838 10362 22862 10364
rect 22918 10362 22924 10364
rect 22678 10310 22680 10362
rect 22860 10310 22862 10362
rect 22616 10308 22622 10310
rect 22678 10308 22702 10310
rect 22758 10308 22782 10310
rect 22838 10308 22862 10310
rect 22918 10308 22924 10310
rect 22616 10299 22924 10308
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22480 9722 22508 10202
rect 22558 10160 22614 10169
rect 22614 10130 22692 10146
rect 22614 10124 22704 10130
rect 22614 10118 22652 10124
rect 22558 10095 22614 10104
rect 22652 10066 22704 10072
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22616 9276 22924 9285
rect 22616 9274 22622 9276
rect 22678 9274 22702 9276
rect 22758 9274 22782 9276
rect 22838 9274 22862 9276
rect 22918 9274 22924 9276
rect 22678 9222 22680 9274
rect 22860 9222 22862 9274
rect 22616 9220 22622 9222
rect 22678 9220 22702 9222
rect 22758 9220 22782 9222
rect 22838 9220 22862 9222
rect 22918 9220 22924 9222
rect 22616 9211 22924 9220
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22204 9030 22324 9058
rect 22388 9042 22416 9114
rect 22112 8894 22232 8922
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 8090 21864 8230
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 22008 7744 22060 7750
rect 22006 7712 22008 7721
rect 22060 7712 22062 7721
rect 22006 7647 22062 7656
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21652 6798 21680 6938
rect 21928 6798 21956 7482
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21744 6322 21772 6734
rect 22112 6390 22140 8298
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21192 5234 21220 6190
rect 21744 5914 21772 6258
rect 22204 6236 22232 8894
rect 22296 8838 22324 9030
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22296 7750 22324 8774
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7886 22416 8230
rect 22480 8090 22508 8366
rect 22616 8188 22924 8197
rect 22616 8186 22622 8188
rect 22678 8186 22702 8188
rect 22758 8186 22782 8188
rect 22838 8186 22862 8188
rect 22918 8186 22924 8188
rect 22678 8134 22680 8186
rect 22860 8134 22862 8186
rect 22616 8132 22622 8134
rect 22678 8132 22702 8134
rect 22758 8132 22782 8134
rect 22838 8132 22862 8134
rect 22918 8132 22924 8134
rect 22616 8123 22924 8132
rect 23032 8090 23060 12038
rect 23492 11354 23520 12135
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 23216 10130 23244 11018
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23124 8974 23152 10066
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 6662 22324 7686
rect 22388 6848 22416 7822
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 7002 22508 7142
rect 22616 7100 22924 7109
rect 22616 7098 22622 7100
rect 22678 7098 22702 7100
rect 22758 7098 22782 7100
rect 22838 7098 22862 7100
rect 22918 7098 22924 7100
rect 22678 7046 22680 7098
rect 22860 7046 22862 7098
rect 22616 7044 22622 7046
rect 22678 7044 22702 7046
rect 22758 7044 22782 7046
rect 22838 7044 22862 7046
rect 22918 7044 22924 7046
rect 22616 7035 22924 7044
rect 23032 7002 23060 7278
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 22560 6860 22612 6866
rect 22388 6820 22560 6848
rect 22560 6802 22612 6808
rect 23124 6730 23152 8910
rect 23216 8838 23244 9930
rect 23308 9178 23336 11222
rect 23584 10198 23612 13942
rect 23676 13870 23704 14214
rect 23860 14006 23888 15030
rect 24228 14618 24256 15030
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 24308 14000 24360 14006
rect 24308 13942 24360 13948
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23860 13734 23888 13942
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23952 13530 23980 13806
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 24320 12850 24348 13942
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 23848 12776 23900 12782
rect 23768 12724 23848 12730
rect 23768 12718 23900 12724
rect 23768 12702 23888 12718
rect 23768 11898 23796 12702
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23860 12306 23888 12582
rect 24412 12434 24440 14214
rect 24780 13394 24808 15982
rect 24872 15570 24900 16594
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24964 14482 24992 17002
rect 25332 16522 25360 17478
rect 25884 17338 25912 17614
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25976 17270 26004 18022
rect 26068 17882 26096 19110
rect 26620 18766 26648 20334
rect 26804 19990 26832 20998
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26792 19984 26844 19990
rect 26792 19926 26844 19932
rect 26896 19922 26924 20742
rect 27252 20392 27304 20398
rect 27252 20334 27304 20340
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26712 19514 26740 19858
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 26988 19378 27016 19654
rect 27264 19514 27292 20334
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 26988 18970 27016 19314
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26700 18148 26752 18154
rect 26700 18090 26752 18096
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25228 16040 25280 16046
rect 25056 15988 25228 15994
rect 25056 15982 25280 15988
rect 25056 15966 25268 15982
rect 25056 15366 25084 15966
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25056 15162 25084 15302
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24228 12406 24440 12434
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23676 11354 23704 11766
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23676 10130 23704 10950
rect 24228 10674 24256 12406
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24504 11558 24532 12038
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24504 11354 24532 11494
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23400 9382 23428 9998
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23400 9042 23428 9318
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23216 6866 23244 7686
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 23124 6458 23152 6666
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23216 6254 23244 6598
rect 23308 6322 23336 7142
rect 23400 6458 23428 8366
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23492 6866 23520 8026
rect 23676 7410 23704 9862
rect 23768 9518 23796 10542
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9586 23888 10406
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24412 9654 24440 9862
rect 24780 9722 24808 13330
rect 25148 12238 25176 13806
rect 25332 13410 25360 16186
rect 25424 16114 25452 17138
rect 25976 16658 26004 17206
rect 26068 17134 26096 17818
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26252 16794 26280 17614
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17134 26372 17478
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 25700 15162 25728 15914
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25700 14362 25728 15098
rect 25976 14414 26004 15846
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25964 14408 26016 14414
rect 25700 14334 25820 14362
rect 25964 14350 26016 14356
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25608 14074 25636 14214
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25424 13546 25452 14010
rect 25424 13518 25636 13546
rect 25332 13382 25544 13410
rect 25608 13394 25636 13518
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12986 25360 13262
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23768 9178 23796 9454
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24780 8090 24808 8230
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24872 8022 24900 12038
rect 24964 11898 24992 12038
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 25056 9586 25084 9998
rect 25148 9994 25176 10406
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8090 25176 8910
rect 25240 8634 25268 12038
rect 25424 11626 25452 12718
rect 25516 12306 25544 13382
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25700 13190 25728 14214
rect 25792 13394 25820 14334
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25884 12170 25912 13874
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25964 11552 26016 11558
rect 25964 11494 26016 11500
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 24860 8016 24912 8022
rect 24860 7958 24912 7964
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23860 7546 23888 7822
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23952 7342 23980 7754
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 23952 6866 23980 7278
rect 24412 7002 24440 7278
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 22112 6208 22232 6236
rect 23204 6248 23256 6254
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 22020 5137 22048 5306
rect 22006 5128 22062 5137
rect 22006 5063 22062 5072
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21008 4826 21036 4966
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 20916 4678 21036 4706
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20916 4282 20944 4558
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20732 2650 20760 3470
rect 21008 3194 21036 4678
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21100 2650 21128 2994
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21088 2644 21140 2650
rect 21088 2586 21140 2592
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20076 2440 20128 2446
rect 20128 2400 20300 2428
rect 20076 2382 20128 2388
rect 18156 734 18368 762
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19444 762 19472 2382
rect 19628 870 19748 898
rect 19628 762 19656 870
rect 19720 800 19748 870
rect 20272 800 20300 2400
rect 20824 800 20852 2450
rect 21284 2394 21312 4558
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3466 21404 3878
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21468 3097 21496 4762
rect 21744 4554 21772 4966
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 21744 4214 21772 4490
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21560 3194 21588 4014
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21652 3466 21680 3878
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 21638 3360 21694 3369
rect 21638 3295 21694 3304
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21454 3088 21510 3097
rect 21652 3058 21680 3295
rect 21454 3023 21456 3032
rect 21508 3023 21510 3032
rect 21640 3052 21692 3058
rect 21456 2994 21508 3000
rect 21640 2994 21692 3000
rect 21744 2854 21772 4014
rect 22112 3369 22140 6208
rect 23204 6190 23256 6196
rect 22192 6112 22244 6118
rect 23296 6112 23348 6118
rect 22244 6060 22324 6066
rect 22192 6054 22324 6060
rect 23296 6054 23348 6060
rect 22204 6038 22324 6054
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22204 4146 22232 5510
rect 22296 4486 22324 6038
rect 22616 6012 22924 6021
rect 22616 6010 22622 6012
rect 22678 6010 22702 6012
rect 22758 6010 22782 6012
rect 22838 6010 22862 6012
rect 22918 6010 22924 6012
rect 22678 5958 22680 6010
rect 22860 5958 22862 6010
rect 22616 5956 22622 5958
rect 22678 5956 22702 5958
rect 22758 5956 22782 5958
rect 22838 5956 22862 5958
rect 22918 5956 22924 5958
rect 22616 5947 22924 5956
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22848 5370 22876 5646
rect 23308 5370 23336 6054
rect 23492 5778 23520 6802
rect 24688 6730 24716 7414
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 22616 4924 22924 4933
rect 22616 4922 22622 4924
rect 22678 4922 22702 4924
rect 22758 4922 22782 4924
rect 22838 4922 22862 4924
rect 22918 4922 22924 4924
rect 22678 4870 22680 4922
rect 22860 4870 22862 4922
rect 22616 4868 22622 4870
rect 22678 4868 22702 4870
rect 22758 4868 22782 4870
rect 22838 4868 22862 4870
rect 22918 4868 22924 4870
rect 22616 4859 22924 4868
rect 23308 4486 23336 4966
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 22296 4214 22324 4422
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22296 3534 22324 4150
rect 22616 3836 22924 3845
rect 22616 3834 22622 3836
rect 22678 3834 22702 3836
rect 22758 3834 22782 3836
rect 22838 3834 22862 3836
rect 22918 3834 22924 3836
rect 22678 3782 22680 3834
rect 22860 3782 22862 3834
rect 22616 3780 22622 3782
rect 22678 3780 22702 3782
rect 22758 3780 22782 3782
rect 22838 3780 22862 3782
rect 22918 3780 22924 3782
rect 22616 3771 22924 3780
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22756 3590 23060 3618
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22098 3360 22154 3369
rect 22098 3295 22154 3304
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21836 2514 21864 2994
rect 22480 2514 22508 3538
rect 22756 3534 22784 3590
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22744 3120 22796 3126
rect 22742 3088 22744 3097
rect 22796 3088 22798 3097
rect 22742 3023 22798 3032
rect 22616 2748 22924 2757
rect 22616 2746 22622 2748
rect 22678 2746 22702 2748
rect 22758 2746 22782 2748
rect 22838 2746 22862 2748
rect 22918 2746 22924 2748
rect 22678 2694 22680 2746
rect 22860 2694 22862 2746
rect 22616 2692 22622 2694
rect 22678 2692 22702 2694
rect 22758 2692 22782 2694
rect 22838 2692 22862 2694
rect 22918 2692 22924 2694
rect 22616 2683 22924 2692
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22192 2440 22244 2446
rect 21928 2400 22192 2428
rect 21284 2366 21404 2394
rect 21376 800 21404 2366
rect 21928 800 21956 2400
rect 22192 2382 22244 2388
rect 22480 870 22600 898
rect 22480 800 22508 870
rect 19444 734 19656 762
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 22572 762 22600 870
rect 22756 762 22784 2450
rect 23032 800 23060 3590
rect 23308 3058 23336 4422
rect 23400 4282 23428 5170
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4554 24072 4966
rect 24032 4548 24084 4554
rect 24032 4490 24084 4496
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23400 3194 23428 4218
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23492 2582 23520 4082
rect 24044 3058 24072 4490
rect 24596 4486 24624 6258
rect 24688 6254 24716 6666
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24688 5778 24716 6190
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24228 4214 24256 4422
rect 24216 4208 24268 4214
rect 24216 4150 24268 4156
rect 24780 4078 24808 4762
rect 24964 4690 24992 7346
rect 25056 4826 25084 7754
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25240 4706 25268 8570
rect 25516 8498 25544 11494
rect 25976 10062 26004 11494
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25608 8634 25636 9522
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25608 7546 25636 7822
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25700 6780 25728 8774
rect 25792 8498 25820 8774
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25964 8356 26016 8362
rect 25964 8298 26016 8304
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25884 7970 25912 8026
rect 25792 7954 25912 7970
rect 25976 7954 26004 8298
rect 25780 7948 25912 7954
rect 25832 7942 25912 7948
rect 25964 7948 26016 7954
rect 25780 7890 25832 7896
rect 25964 7890 26016 7896
rect 26068 7449 26096 14554
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 14074 26188 14214
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26160 13394 26188 14010
rect 26252 13802 26280 16594
rect 26344 16114 26372 17070
rect 26712 16114 26740 18090
rect 26988 17202 27016 18906
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27172 18154 27200 18770
rect 27264 18426 27292 19314
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27160 18148 27212 18154
rect 27160 18090 27212 18096
rect 27356 17338 27384 20198
rect 27540 20058 27568 20878
rect 28092 20534 28120 23122
rect 28920 22098 28948 25978
rect 29000 25424 29052 25430
rect 29000 25366 29052 25372
rect 29012 24818 29040 25366
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24886 29132 25094
rect 29092 24880 29144 24886
rect 29092 24822 29144 24828
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 29000 22976 29052 22982
rect 29000 22918 29052 22924
rect 29012 22760 29040 22918
rect 29104 22760 29132 24822
rect 29288 24818 29316 26182
rect 29656 26042 29684 26318
rect 29838 26140 30146 26149
rect 29838 26138 29844 26140
rect 29900 26138 29924 26140
rect 29980 26138 30004 26140
rect 30060 26138 30084 26140
rect 30140 26138 30146 26140
rect 29900 26086 29902 26138
rect 30082 26086 30084 26138
rect 29838 26084 29844 26086
rect 29900 26084 29924 26086
rect 29980 26084 30004 26086
rect 30060 26084 30084 26086
rect 30140 26084 30146 26086
rect 29838 26075 30146 26084
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 29840 25922 29868 25978
rect 30208 25922 30236 26862
rect 29748 25894 29868 25922
rect 30024 25906 30236 25922
rect 29920 25900 29972 25906
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 29564 25226 29592 25774
rect 29552 25220 29604 25226
rect 29552 25162 29604 25168
rect 29564 24954 29592 25162
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 29748 24886 29776 25894
rect 29920 25842 29972 25848
rect 30012 25900 30236 25906
rect 30064 25894 30236 25900
rect 30012 25842 30064 25848
rect 29932 25498 29960 25842
rect 29920 25492 29972 25498
rect 29920 25434 29972 25440
rect 30208 25294 30236 25894
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 29838 25052 30146 25061
rect 29838 25050 29844 25052
rect 29900 25050 29924 25052
rect 29980 25050 30004 25052
rect 30060 25050 30084 25052
rect 30140 25050 30146 25052
rect 29900 24998 29902 25050
rect 30082 24998 30084 25050
rect 29838 24996 29844 24998
rect 29900 24996 29924 24998
rect 29980 24996 30004 24998
rect 30060 24996 30084 24998
rect 30140 24996 30146 24998
rect 29838 24987 30146 24996
rect 29736 24880 29788 24886
rect 29736 24822 29788 24828
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 30300 24614 30328 26862
rect 30392 25498 30420 26998
rect 45192 26920 45244 26926
rect 45192 26862 45244 26868
rect 46296 26920 46348 26926
rect 46296 26862 46348 26868
rect 46664 26920 46716 26926
rect 46664 26862 46716 26868
rect 48136 26920 48188 26926
rect 48136 26862 48188 26868
rect 49240 26920 49292 26926
rect 49240 26862 49292 26868
rect 50804 26920 50856 26926
rect 50804 26862 50856 26868
rect 51080 26920 51132 26926
rect 51080 26862 51132 26868
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 30840 26240 30892 26246
rect 31220 26234 31248 26726
rect 37060 26684 37368 26693
rect 37060 26682 37066 26684
rect 37122 26682 37146 26684
rect 37202 26682 37226 26684
rect 37282 26682 37306 26684
rect 37362 26682 37368 26684
rect 37122 26630 37124 26682
rect 37304 26630 37306 26682
rect 37060 26628 37066 26630
rect 37122 26628 37146 26630
rect 37202 26628 37226 26630
rect 37282 26628 37306 26630
rect 37362 26628 37368 26630
rect 37060 26619 37368 26628
rect 44180 26308 44232 26314
rect 44180 26250 44232 26256
rect 31576 26240 31628 26246
rect 31220 26206 31340 26234
rect 30840 26182 30892 26188
rect 30852 25838 30880 26182
rect 31312 25838 31340 26206
rect 31576 26182 31628 26188
rect 30840 25832 30892 25838
rect 30840 25774 30892 25780
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 30656 25696 30708 25702
rect 30656 25638 30708 25644
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30288 24608 30340 24614
rect 30288 24550 30340 24556
rect 29838 23964 30146 23973
rect 29838 23962 29844 23964
rect 29900 23962 29924 23964
rect 29980 23962 30004 23964
rect 30060 23962 30084 23964
rect 30140 23962 30146 23964
rect 29900 23910 29902 23962
rect 30082 23910 30084 23962
rect 29838 23908 29844 23910
rect 29900 23908 29924 23910
rect 29980 23908 30004 23910
rect 30060 23908 30084 23910
rect 30140 23908 30146 23910
rect 29838 23899 30146 23908
rect 30392 23798 30420 25434
rect 29736 23792 29788 23798
rect 29736 23734 29788 23740
rect 30380 23792 30432 23798
rect 30380 23734 30432 23740
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 29196 22778 29224 23598
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 29656 22982 29684 23122
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 29012 22732 29132 22760
rect 29104 22506 29132 22732
rect 29184 22772 29236 22778
rect 29184 22714 29236 22720
rect 29092 22500 29144 22506
rect 29092 22442 29144 22448
rect 28908 22092 28960 22098
rect 29104 22094 29132 22442
rect 28908 22034 28960 22040
rect 29012 22066 29132 22094
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28276 21146 28304 21898
rect 29012 21622 29040 22066
rect 29276 21888 29328 21894
rect 29276 21830 29328 21836
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28080 20528 28132 20534
rect 28080 20470 28132 20476
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27540 18630 27568 19314
rect 27816 18766 27844 19858
rect 28368 19666 28396 21286
rect 28460 21146 28488 21286
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 29012 20398 29040 21558
rect 29288 21554 29316 21830
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29656 21418 29684 22918
rect 29748 22574 29776 23734
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30484 23050 30512 23462
rect 30668 23186 30696 25638
rect 30852 24954 30880 25774
rect 30840 24948 30892 24954
rect 30840 24890 30892 24896
rect 30840 24744 30892 24750
rect 30840 24686 30892 24692
rect 30748 23520 30800 23526
rect 30748 23462 30800 23468
rect 30656 23180 30708 23186
rect 30656 23122 30708 23128
rect 30472 23044 30524 23050
rect 30472 22986 30524 22992
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 29838 22876 30146 22885
rect 29838 22874 29844 22876
rect 29900 22874 29924 22876
rect 29980 22874 30004 22876
rect 30060 22874 30084 22876
rect 30140 22874 30146 22876
rect 29900 22822 29902 22874
rect 30082 22822 30084 22874
rect 29838 22820 29844 22822
rect 29900 22820 29924 22822
rect 29980 22820 30004 22822
rect 30060 22820 30084 22822
rect 30140 22820 30146 22822
rect 29838 22811 30146 22820
rect 29736 22568 29788 22574
rect 29736 22510 29788 22516
rect 30104 22568 30156 22574
rect 30156 22528 30236 22556
rect 30104 22510 30156 22516
rect 29838 21788 30146 21797
rect 29838 21786 29844 21788
rect 29900 21786 29924 21788
rect 29980 21786 30004 21788
rect 30060 21786 30084 21788
rect 30140 21786 30146 21788
rect 29900 21734 29902 21786
rect 30082 21734 30084 21786
rect 29838 21732 29844 21734
rect 29900 21732 29924 21734
rect 29980 21732 30004 21734
rect 30060 21732 30084 21734
rect 30140 21732 30146 21734
rect 29838 21723 30146 21732
rect 30208 21690 30236 22528
rect 30196 21684 30248 21690
rect 30196 21626 30248 21632
rect 30392 21554 30420 22918
rect 30484 22556 30512 22986
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30576 22778 30604 22918
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30564 22568 30616 22574
rect 30484 22528 30564 22556
rect 30760 22522 30788 23462
rect 30564 22510 30616 22516
rect 30668 22506 30788 22522
rect 30656 22500 30788 22506
rect 30708 22494 30788 22500
rect 30656 22442 30708 22448
rect 30852 21962 30880 24686
rect 31312 23866 31340 25774
rect 31588 25770 31616 26182
rect 31576 25764 31628 25770
rect 31576 25706 31628 25712
rect 31588 23866 31616 25706
rect 31668 25696 31720 25702
rect 31668 25638 31720 25644
rect 32128 25696 32180 25702
rect 32128 25638 32180 25644
rect 31680 25498 31708 25638
rect 31668 25492 31720 25498
rect 31668 25434 31720 25440
rect 32140 25294 32168 25638
rect 37060 25596 37368 25605
rect 37060 25594 37066 25596
rect 37122 25594 37146 25596
rect 37202 25594 37226 25596
rect 37282 25594 37306 25596
rect 37362 25594 37368 25596
rect 37122 25542 37124 25594
rect 37304 25542 37306 25594
rect 37060 25540 37066 25542
rect 37122 25540 37146 25542
rect 37202 25540 37226 25542
rect 37282 25540 37306 25542
rect 37362 25540 37368 25542
rect 37060 25531 37368 25540
rect 38384 25356 38436 25362
rect 38384 25298 38436 25304
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 37060 24508 37368 24517
rect 37060 24506 37066 24508
rect 37122 24506 37146 24508
rect 37202 24506 37226 24508
rect 37282 24506 37306 24508
rect 37362 24506 37368 24508
rect 37122 24454 37124 24506
rect 37304 24454 37306 24506
rect 37060 24452 37066 24454
rect 37122 24452 37146 24454
rect 37202 24452 37226 24454
rect 37282 24452 37306 24454
rect 37362 24452 37368 24454
rect 37060 24443 37368 24452
rect 33508 24200 33560 24206
rect 33508 24142 33560 24148
rect 33692 24200 33744 24206
rect 33692 24142 33744 24148
rect 35992 24200 36044 24206
rect 35992 24142 36044 24148
rect 37556 24200 37608 24206
rect 37556 24142 37608 24148
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 31588 23526 31616 23802
rect 32968 23730 32996 24006
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 32036 23724 32088 23730
rect 32036 23666 32088 23672
rect 32956 23724 33008 23730
rect 32956 23666 33008 23672
rect 31576 23520 31628 23526
rect 31576 23462 31628 23468
rect 31588 23254 31616 23462
rect 31576 23248 31628 23254
rect 31496 23196 31576 23202
rect 31496 23190 31628 23196
rect 31496 23174 31616 23190
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30840 21956 30892 21962
rect 30840 21898 30892 21904
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30380 21548 30432 21554
rect 30380 21490 30432 21496
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28460 19786 28488 20198
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 28368 19638 28488 19666
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18834 28396 19110
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 27804 18760 27856 18766
rect 27804 18702 27856 18708
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27448 18426 27476 18566
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26792 17060 26844 17066
rect 26792 17002 26844 17008
rect 26804 16250 26832 17002
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26896 16590 26924 16934
rect 26988 16794 27016 17138
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26436 13530 26464 14350
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26252 12986 26280 13262
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26252 12306 26280 12922
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26436 12442 26464 12786
rect 26424 12436 26476 12442
rect 26712 12434 26740 16050
rect 27264 13870 27292 16186
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26896 12434 26924 12650
rect 26424 12378 26476 12384
rect 26528 12406 26924 12434
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26528 11694 26556 12406
rect 26516 11688 26568 11694
rect 26516 11630 26568 11636
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26344 8838 26372 10610
rect 26436 10606 26464 11086
rect 26528 11082 26556 11630
rect 26516 11076 26568 11082
rect 26516 11018 26568 11024
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26436 10266 26464 10542
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 7954 26188 8230
rect 26148 7948 26200 7954
rect 26148 7890 26200 7896
rect 26344 7834 26372 8774
rect 26436 8498 26464 9318
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26344 7818 26464 7834
rect 26344 7812 26476 7818
rect 26344 7806 26424 7812
rect 26424 7754 26476 7760
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26422 7712 26478 7721
rect 26054 7440 26110 7449
rect 26054 7375 26110 7384
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25884 6798 25912 7142
rect 26344 6866 26372 7686
rect 26422 7647 26478 7656
rect 26436 7546 26464 7647
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 25780 6792 25832 6798
rect 25700 6752 25780 6780
rect 25780 6734 25832 6740
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25608 5370 25636 5578
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25884 5234 25912 6734
rect 26344 6458 26372 6802
rect 26332 6452 26384 6458
rect 26332 6394 26384 6400
rect 26528 6322 26556 9318
rect 26620 9042 26648 9862
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26620 6866 26648 7686
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26608 5772 26660 5778
rect 26608 5714 26660 5720
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26252 5234 26280 5510
rect 26620 5370 26648 5714
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 25332 4826 25360 5102
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 25044 4684 25096 4690
rect 25240 4678 25452 4706
rect 25044 4626 25096 4632
rect 25056 4570 25084 4626
rect 24964 4542 25084 4570
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 24964 4146 24992 4542
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 25044 4140 25096 4146
rect 25096 4100 25176 4128
rect 25044 4082 25096 4088
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24136 3738 24164 4014
rect 25044 4004 25096 4010
rect 25044 3946 25096 3952
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24136 3194 24164 3402
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24228 3058 24256 3334
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23584 800 23612 2858
rect 24320 2774 24348 3062
rect 24136 2746 24348 2774
rect 24136 800 24164 2746
rect 24412 2650 24440 3878
rect 25056 3194 25084 3946
rect 25148 3738 25176 4100
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25240 3194 25268 4558
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24676 3120 24728 3126
rect 24676 3062 24728 3068
rect 24688 2990 24716 3062
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 25332 2774 25360 4558
rect 25424 4146 25452 4678
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25332 2746 25452 2774
rect 25424 2650 25452 2746
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25516 2446 25544 3674
rect 26252 3466 26280 4422
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 26528 3194 26556 4558
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26620 2961 26648 3878
rect 26606 2952 26662 2961
rect 26712 2922 26740 11018
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10674 27292 10950
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27172 10130 27200 10406
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27172 9654 27200 10066
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26804 7478 26832 7686
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26804 6662 26832 6802
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26896 5778 26924 7686
rect 26988 6866 27016 7822
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 27080 6662 27108 8842
rect 27172 8634 27200 9590
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27448 8294 27476 17070
rect 27540 11354 27568 18566
rect 28460 16658 28488 19638
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 27620 16040 27672 16046
rect 27620 15982 27672 15988
rect 27632 15638 27660 15982
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27724 15638 27752 15846
rect 27620 15632 27672 15638
rect 27620 15574 27672 15580
rect 27712 15632 27764 15638
rect 27712 15574 27764 15580
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27632 12434 27660 13738
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27724 13258 27752 13670
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27712 13252 27764 13258
rect 27712 13194 27764 13200
rect 27632 12406 27752 12434
rect 27620 12232 27672 12238
rect 27618 12200 27620 12209
rect 27672 12200 27674 12209
rect 27618 12135 27674 12144
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27632 10742 27660 12038
rect 27724 11558 27752 12406
rect 27816 12102 27844 13262
rect 28000 12850 28028 16390
rect 28460 15026 28488 16594
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28644 15026 28672 16390
rect 28736 15570 28764 19450
rect 28816 17128 28868 17134
rect 28816 17070 28868 17076
rect 28828 16250 28856 17070
rect 28816 16244 28868 16250
rect 28816 16186 28868 16192
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28724 14272 28776 14278
rect 28724 14214 28776 14220
rect 28736 14006 28764 14214
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28092 13326 28120 13670
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 28448 12640 28500 12646
rect 28448 12582 28500 12588
rect 28460 12434 28488 12582
rect 28644 12442 28672 13194
rect 29012 12986 29040 20334
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 29104 17134 29132 18906
rect 29472 18902 29500 20198
rect 29460 18896 29512 18902
rect 29460 18838 29512 18844
rect 29656 17218 29684 21354
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20602 29776 20878
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 29838 20700 30146 20709
rect 29838 20698 29844 20700
rect 29900 20698 29924 20700
rect 29980 20698 30004 20700
rect 30060 20698 30084 20700
rect 30140 20698 30146 20700
rect 29900 20646 29902 20698
rect 30082 20646 30084 20698
rect 29838 20644 29844 20646
rect 29900 20644 29924 20646
rect 29980 20644 30004 20646
rect 30060 20644 30084 20646
rect 30140 20644 30146 20646
rect 29838 20635 30146 20644
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 30392 19854 30420 20742
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 29838 19612 30146 19621
rect 29838 19610 29844 19612
rect 29900 19610 29924 19612
rect 29980 19610 30004 19612
rect 30060 19610 30084 19612
rect 30140 19610 30146 19612
rect 29900 19558 29902 19610
rect 30082 19558 30084 19610
rect 29838 19556 29844 19558
rect 29900 19556 29924 19558
rect 29980 19556 30004 19558
rect 30060 19556 30084 19558
rect 30140 19556 30146 19558
rect 29838 19547 30146 19556
rect 30564 19372 30616 19378
rect 30564 19314 30616 19320
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30116 18970 30144 19246
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 29838 18524 30146 18533
rect 29838 18522 29844 18524
rect 29900 18522 29924 18524
rect 29980 18522 30004 18524
rect 30060 18522 30084 18524
rect 30140 18522 30146 18524
rect 29900 18470 29902 18522
rect 30082 18470 30084 18522
rect 29838 18468 29844 18470
rect 29900 18468 29924 18470
rect 29980 18468 30004 18470
rect 30060 18468 30084 18470
rect 30140 18468 30146 18470
rect 29838 18459 30146 18468
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29748 17338 29776 17478
rect 29838 17436 30146 17445
rect 29838 17434 29844 17436
rect 29900 17434 29924 17436
rect 29980 17434 30004 17436
rect 30060 17434 30084 17436
rect 30140 17434 30146 17436
rect 29900 17382 29902 17434
rect 30082 17382 30084 17434
rect 29838 17380 29844 17382
rect 29900 17380 29924 17382
rect 29980 17380 30004 17382
rect 30060 17380 30084 17382
rect 30140 17380 30146 17382
rect 29838 17371 30146 17380
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29552 17196 29604 17202
rect 29656 17190 29776 17218
rect 29552 17138 29604 17144
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 16590 29500 16934
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29564 16250 29592 17138
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29552 16244 29604 16250
rect 29552 16186 29604 16192
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 28908 12708 28960 12714
rect 28908 12650 28960 12656
rect 28368 12406 28488 12434
rect 28632 12436 28684 12442
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27724 10674 27752 11494
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27724 10554 27752 10610
rect 27632 10526 27752 10554
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27540 9382 27568 9998
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27436 8288 27488 8294
rect 27632 8276 27660 10526
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27724 8974 27752 9998
rect 27816 9178 27844 11086
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27908 9586 27936 11018
rect 27988 10804 28040 10810
rect 27988 10746 28040 10752
rect 28000 10130 28028 10746
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 28000 9042 28028 10066
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 27988 9036 28040 9042
rect 27988 8978 28040 8984
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27724 8634 27752 8910
rect 27908 8634 27936 8910
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27436 8230 27488 8236
rect 27540 8248 27660 8276
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 27172 5710 27200 6734
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27158 4176 27214 4185
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26976 4140 27028 4146
rect 27158 4111 27214 4120
rect 26976 4082 27028 4088
rect 26804 3641 26832 4082
rect 26790 3632 26846 3641
rect 26790 3567 26846 3576
rect 26606 2887 26662 2896
rect 26700 2916 26752 2922
rect 26700 2858 26752 2864
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 24584 2440 24636 2446
rect 25228 2440 25280 2446
rect 24636 2400 24716 2428
rect 24584 2382 24636 2388
rect 24688 800 24716 2400
rect 25228 2382 25280 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25240 800 25268 2382
rect 25884 1170 25912 2450
rect 26332 2100 26384 2106
rect 26332 2042 26384 2048
rect 25792 1142 25912 1170
rect 25792 800 25820 1142
rect 26344 800 26372 2042
rect 26896 800 26924 2858
rect 26988 2106 27016 4082
rect 27172 4010 27200 4111
rect 27252 4072 27304 4078
rect 27252 4014 27304 4020
rect 27160 4004 27212 4010
rect 27160 3946 27212 3952
rect 27264 2446 27292 4014
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 2446 27384 3334
rect 27448 2446 27476 8230
rect 27540 7410 27568 8248
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 28000 7410 28028 7890
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 27620 6860 27672 6866
rect 27540 6820 27620 6848
rect 27540 6322 27568 6820
rect 27620 6802 27672 6808
rect 27988 6860 28040 6866
rect 27988 6802 28040 6808
rect 28000 6458 28028 6802
rect 28092 6798 28120 9862
rect 28184 8922 28212 10066
rect 28276 9042 28304 12174
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 28184 8906 28304 8922
rect 28184 8900 28316 8906
rect 28184 8894 28264 8900
rect 28264 8842 28316 8848
rect 28368 8498 28396 12406
rect 28632 12378 28684 12384
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28736 11286 28764 11630
rect 28920 11286 28948 12650
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 29012 12322 29040 12582
rect 29196 12442 29224 12718
rect 29184 12436 29236 12442
rect 29184 12378 29236 12384
rect 29012 12306 29224 12322
rect 29012 12300 29236 12306
rect 29012 12294 29184 12300
rect 29184 12242 29236 12248
rect 29288 12050 29316 15302
rect 29380 15162 29408 16050
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29656 12866 29684 16730
rect 29748 14618 29776 17190
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30116 16658 30144 16730
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 29838 16348 30146 16357
rect 29838 16346 29844 16348
rect 29900 16346 29924 16348
rect 29980 16346 30004 16348
rect 30060 16346 30084 16348
rect 30140 16346 30146 16348
rect 29900 16294 29902 16346
rect 30082 16294 30084 16346
rect 29838 16292 29844 16294
rect 29900 16292 29924 16294
rect 29980 16292 30004 16294
rect 30060 16292 30084 16294
rect 30140 16292 30146 16294
rect 29838 16283 30146 16292
rect 30392 15638 30420 17614
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30484 16590 30512 17206
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30380 15632 30432 15638
rect 30380 15574 30432 15580
rect 30484 15502 30512 16526
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 29838 15260 30146 15269
rect 29838 15258 29844 15260
rect 29900 15258 29924 15260
rect 29980 15258 30004 15260
rect 30060 15258 30084 15260
rect 30140 15258 30146 15260
rect 29900 15206 29902 15258
rect 30082 15206 30084 15258
rect 29838 15204 29844 15206
rect 29900 15204 29924 15206
rect 29980 15204 30004 15206
rect 30060 15204 30084 15206
rect 30140 15204 30146 15206
rect 29838 15195 30146 15204
rect 30484 15178 30512 15438
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30392 15150 30512 15178
rect 30116 14618 30144 15098
rect 30196 15020 30248 15026
rect 30196 14962 30248 14968
rect 29736 14612 29788 14618
rect 29736 14554 29788 14560
rect 30104 14612 30156 14618
rect 30104 14554 30156 14560
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 14074 29776 14350
rect 29838 14172 30146 14181
rect 29838 14170 29844 14172
rect 29900 14170 29924 14172
rect 29980 14170 30004 14172
rect 30060 14170 30084 14172
rect 30140 14170 30146 14172
rect 29900 14118 29902 14170
rect 30082 14118 30084 14170
rect 29838 14116 29844 14118
rect 29900 14116 29924 14118
rect 29980 14116 30004 14118
rect 30060 14116 30084 14118
rect 30140 14116 30146 14118
rect 29838 14107 30146 14116
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29920 13728 29972 13734
rect 29920 13670 29972 13676
rect 29932 13530 29960 13670
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29564 12838 29684 12866
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 29196 12022 29316 12050
rect 29196 11762 29224 12022
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 28724 11280 28776 11286
rect 28724 11222 28776 11228
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28540 10464 28592 10470
rect 28540 10406 28592 10412
rect 28552 9042 28580 10406
rect 29012 10130 29040 10950
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28736 8974 28764 9998
rect 29012 9586 29040 10066
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29104 9466 29132 11494
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29012 9438 29132 9466
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7002 28580 7822
rect 28644 7818 28672 8774
rect 28908 8424 28960 8430
rect 28908 8366 28960 8372
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28632 7812 28684 7818
rect 28632 7754 28684 7760
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28644 6458 28672 7754
rect 28736 7410 28764 8230
rect 28920 8090 28948 8366
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 28644 5778 28672 6394
rect 28920 5914 28948 6598
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 28632 5772 28684 5778
rect 28632 5714 28684 5720
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28276 5302 28304 5510
rect 28264 5296 28316 5302
rect 28264 5238 28316 5244
rect 28828 4826 28856 5646
rect 28906 5128 28962 5137
rect 28906 5063 28962 5072
rect 28920 4826 28948 5063
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 28172 4752 28224 4758
rect 28172 4694 28224 4700
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27540 4146 27568 4626
rect 28184 4622 28212 4694
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 27620 4480 27672 4486
rect 28356 4480 28408 4486
rect 27672 4440 27752 4468
rect 27620 4422 27672 4428
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27540 2582 27568 4082
rect 27724 3618 27752 4440
rect 28356 4422 28408 4428
rect 27896 4276 27948 4282
rect 28080 4276 28132 4282
rect 27948 4236 28080 4264
rect 27896 4218 27948 4224
rect 28080 4218 28132 4224
rect 28368 4146 28396 4422
rect 29012 4162 29040 9438
rect 29196 8838 29224 11018
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 29104 6390 29132 7142
rect 29092 6384 29144 6390
rect 29092 6326 29144 6332
rect 29184 4480 29236 4486
rect 29184 4422 29236 4428
rect 29196 4214 29224 4422
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28724 4140 28776 4146
rect 28920 4134 29040 4162
rect 29184 4208 29236 4214
rect 29184 4150 29236 4156
rect 28920 4128 28948 4134
rect 28776 4100 28948 4128
rect 28724 4082 28776 4088
rect 28080 4004 28132 4010
rect 28080 3946 28132 3952
rect 28092 3618 28120 3946
rect 27724 3590 28120 3618
rect 27724 3534 27752 3590
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27632 2650 27660 2926
rect 28184 2774 28212 4082
rect 28460 3466 28488 4082
rect 28816 4004 28868 4010
rect 28816 3946 28868 3952
rect 28828 3738 28856 3946
rect 28816 3732 28868 3738
rect 28816 3674 28868 3680
rect 28448 3460 28500 3466
rect 28448 3402 28500 3408
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29288 3194 29316 3334
rect 29276 3188 29328 3194
rect 29276 3130 29328 3136
rect 28540 2984 28592 2990
rect 29368 2984 29420 2990
rect 28540 2926 28592 2932
rect 29196 2944 29368 2972
rect 28000 2746 28212 2774
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 26976 2100 27028 2106
rect 26976 2042 27028 2048
rect 27724 1442 27752 2450
rect 27448 1414 27752 1442
rect 27448 800 27476 1414
rect 28000 800 28028 2746
rect 28552 800 28580 2926
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 29104 2446 29132 2790
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 29196 1442 29224 2944
rect 29368 2926 29420 2932
rect 29472 2774 29500 12378
rect 29564 10470 29592 12838
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29656 11830 29684 12718
rect 29748 12646 29776 13262
rect 29838 13084 30146 13093
rect 29838 13082 29844 13084
rect 29900 13082 29924 13084
rect 29980 13082 30004 13084
rect 30060 13082 30084 13084
rect 30140 13082 30146 13084
rect 29900 13030 29902 13082
rect 30082 13030 30084 13082
rect 29838 13028 29844 13030
rect 29900 13028 29924 13030
rect 29980 13028 30004 13030
rect 30060 13028 30084 13030
rect 30140 13028 30146 13030
rect 29838 13019 30146 13028
rect 29736 12640 29788 12646
rect 29736 12582 29788 12588
rect 29748 12442 29776 12582
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29748 11898 29776 12378
rect 29838 11996 30146 12005
rect 29838 11994 29844 11996
rect 29900 11994 29924 11996
rect 29980 11994 30004 11996
rect 30060 11994 30084 11996
rect 30140 11994 30146 11996
rect 29900 11942 29902 11994
rect 30082 11942 30084 11994
rect 29838 11940 29844 11942
rect 29900 11940 29924 11942
rect 29980 11940 30004 11942
rect 30060 11940 30084 11942
rect 30140 11940 30146 11942
rect 29838 11931 30146 11940
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 29644 11824 29696 11830
rect 29644 11766 29696 11772
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29656 8090 29684 11766
rect 30104 11688 30156 11694
rect 30104 11630 30156 11636
rect 30116 11354 30144 11630
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 29838 10908 30146 10917
rect 29838 10906 29844 10908
rect 29900 10906 29924 10908
rect 29980 10906 30004 10908
rect 30060 10906 30084 10908
rect 30140 10906 30146 10908
rect 29900 10854 29902 10906
rect 30082 10854 30084 10906
rect 29838 10852 29844 10854
rect 29900 10852 29924 10854
rect 29980 10852 30004 10854
rect 30060 10852 30084 10854
rect 30140 10852 30146 10854
rect 29838 10843 30146 10852
rect 29736 10736 29788 10742
rect 29736 10678 29788 10684
rect 29748 10130 29776 10678
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29748 9178 29776 10066
rect 29838 9820 30146 9829
rect 29838 9818 29844 9820
rect 29900 9818 29924 9820
rect 29980 9818 30004 9820
rect 30060 9818 30084 9820
rect 30140 9818 30146 9820
rect 29900 9766 29902 9818
rect 30082 9766 30084 9818
rect 29838 9764 29844 9766
rect 29900 9764 29924 9766
rect 29980 9764 30004 9766
rect 30060 9764 30084 9766
rect 30140 9764 30146 9766
rect 29838 9755 30146 9764
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29838 8732 30146 8741
rect 29838 8730 29844 8732
rect 29900 8730 29924 8732
rect 29980 8730 30004 8732
rect 30060 8730 30084 8732
rect 30140 8730 30146 8732
rect 29900 8678 29902 8730
rect 30082 8678 30084 8730
rect 29838 8676 29844 8678
rect 29900 8676 29924 8678
rect 29980 8676 30004 8678
rect 30060 8676 30084 8678
rect 30140 8676 30146 8678
rect 29838 8667 30146 8676
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29656 7954 29684 8026
rect 29644 7948 29696 7954
rect 29644 7890 29696 7896
rect 30116 7750 30144 8366
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 29838 7644 30146 7653
rect 29838 7642 29844 7644
rect 29900 7642 29924 7644
rect 29980 7642 30004 7644
rect 30060 7642 30084 7644
rect 30140 7642 30146 7644
rect 29900 7590 29902 7642
rect 30082 7590 30084 7642
rect 29838 7588 29844 7590
rect 29900 7588 29924 7590
rect 29980 7588 30004 7590
rect 30060 7588 30084 7590
rect 30140 7588 30146 7590
rect 29838 7579 30146 7588
rect 29838 6556 30146 6565
rect 29838 6554 29844 6556
rect 29900 6554 29924 6556
rect 29980 6554 30004 6556
rect 30060 6554 30084 6556
rect 30140 6554 30146 6556
rect 29900 6502 29902 6554
rect 30082 6502 30084 6554
rect 29838 6500 29844 6502
rect 29900 6500 29924 6502
rect 29980 6500 30004 6502
rect 30060 6500 30084 6502
rect 30140 6500 30146 6502
rect 29838 6491 30146 6500
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 4622 29592 5510
rect 29838 5468 30146 5477
rect 29838 5466 29844 5468
rect 29900 5466 29924 5468
rect 29980 5466 30004 5468
rect 30060 5466 30084 5468
rect 30140 5466 30146 5468
rect 29900 5414 29902 5466
rect 30082 5414 30084 5466
rect 29838 5412 29844 5414
rect 29900 5412 29924 5414
rect 29980 5412 30004 5414
rect 30060 5412 30084 5414
rect 30140 5412 30146 5414
rect 29838 5403 30146 5412
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29656 4214 29684 4422
rect 29644 4208 29696 4214
rect 29644 4150 29696 4156
rect 29656 4010 29684 4150
rect 29748 4010 29776 4558
rect 29838 4380 30146 4389
rect 29838 4378 29844 4380
rect 29900 4378 29924 4380
rect 29980 4378 30004 4380
rect 30060 4378 30084 4380
rect 30140 4378 30146 4380
rect 29900 4326 29902 4378
rect 30082 4326 30084 4378
rect 29838 4324 29844 4326
rect 29900 4324 29924 4326
rect 29980 4324 30004 4326
rect 30060 4324 30084 4326
rect 30140 4324 30146 4326
rect 29838 4315 30146 4324
rect 30010 4176 30066 4185
rect 30010 4111 30012 4120
rect 30064 4111 30066 4120
rect 30012 4082 30064 4088
rect 29644 4004 29696 4010
rect 29644 3946 29696 3952
rect 29736 4004 29788 4010
rect 29736 3946 29788 3952
rect 30208 3505 30236 14962
rect 30288 14408 30340 14414
rect 30392 14362 30420 15150
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30340 14356 30420 14362
rect 30288 14350 30420 14356
rect 30300 14334 30420 14350
rect 30300 14278 30328 14334
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30484 13802 30512 15030
rect 30472 13796 30524 13802
rect 30472 13738 30524 13744
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30392 12918 30420 13466
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30484 12730 30512 13194
rect 30300 12702 30512 12730
rect 30300 12442 30328 12702
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30576 11558 30604 19314
rect 30668 19174 30696 21626
rect 30944 20602 30972 22510
rect 31036 22030 31064 22918
rect 31392 22500 31444 22506
rect 31392 22442 31444 22448
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 31036 19514 31064 21286
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 31128 20058 31156 20334
rect 31116 20052 31168 20058
rect 31116 19994 31168 20000
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31128 19446 31156 19654
rect 31116 19440 31168 19446
rect 31116 19382 31168 19388
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30668 16794 30696 19110
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30852 17338 30880 17614
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 30840 17332 30892 17338
rect 30840 17274 30892 17280
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 30944 16794 30972 16934
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 31220 16658 31248 17478
rect 31208 16652 31260 16658
rect 31208 16594 31260 16600
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 15638 30788 16390
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 30852 15638 30880 16050
rect 30748 15632 30800 15638
rect 30748 15574 30800 15580
rect 30840 15632 30892 15638
rect 30840 15574 30892 15580
rect 30748 15496 30800 15502
rect 30748 15438 30800 15444
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 30668 14074 30696 14214
rect 30656 14068 30708 14074
rect 30656 14010 30708 14016
rect 30668 12986 30696 14010
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30668 12306 30696 12582
rect 30656 12300 30708 12306
rect 30656 12242 30708 12248
rect 30564 11552 30616 11558
rect 30564 11494 30616 11500
rect 30760 11218 30788 15438
rect 31220 15434 31248 16594
rect 31208 15428 31260 15434
rect 31208 15370 31260 15376
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30852 13870 30880 14010
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 30944 13258 30972 14350
rect 31024 14340 31076 14346
rect 31024 14282 31076 14288
rect 31036 13938 31064 14282
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 30932 13252 30984 13258
rect 30932 13194 30984 13200
rect 30944 12986 30972 13194
rect 31024 13184 31076 13190
rect 31024 13126 31076 13132
rect 31036 12986 31064 13126
rect 30932 12980 30984 12986
rect 30932 12922 30984 12928
rect 31024 12980 31076 12986
rect 31024 12922 31076 12928
rect 31128 12714 31156 13806
rect 31220 13462 31248 14350
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 31312 12782 31340 21898
rect 31404 21690 31432 22442
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31404 19854 31432 20198
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31392 19304 31444 19310
rect 31392 19246 31444 19252
rect 31404 18970 31432 19246
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31496 16658 31524 23174
rect 32048 23118 32076 23666
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 31588 22778 31616 23054
rect 32312 23044 32364 23050
rect 32312 22986 32364 22992
rect 31576 22772 31628 22778
rect 31576 22714 31628 22720
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32140 22166 32168 22510
rect 32324 22166 32352 22986
rect 33152 22710 33180 23802
rect 33520 23322 33548 24142
rect 33704 23866 33732 24142
rect 34336 24064 34388 24070
rect 34336 24006 34388 24012
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 33692 23860 33744 23866
rect 33692 23802 33744 23808
rect 34152 23860 34204 23866
rect 34152 23802 34204 23808
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 34072 23186 34100 23462
rect 34060 23180 34112 23186
rect 34060 23122 34112 23128
rect 34164 23066 34192 23802
rect 34348 23118 34376 24006
rect 35452 23798 35480 24006
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 23118 34560 23462
rect 34072 23038 34192 23066
rect 34336 23112 34388 23118
rect 34336 23054 34388 23060
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 33324 22976 33376 22982
rect 33324 22918 33376 22924
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 33048 22568 33100 22574
rect 33048 22510 33100 22516
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32128 22160 32180 22166
rect 32128 22102 32180 22108
rect 32312 22160 32364 22166
rect 32312 22102 32364 22108
rect 32416 22098 32444 22374
rect 33060 22098 33088 22510
rect 33336 22098 33364 22918
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 22166 33456 22578
rect 34072 22574 34100 23038
rect 34348 22642 34376 23054
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34336 22636 34388 22642
rect 34336 22578 34388 22584
rect 34624 22574 34652 22986
rect 35544 22982 35572 23666
rect 35716 23520 35768 23526
rect 35716 23462 35768 23468
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 35532 22976 35584 22982
rect 35584 22936 35664 22964
rect 35532 22918 35584 22924
rect 34808 22778 34836 22918
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34060 22568 34112 22574
rect 34060 22510 34112 22516
rect 34152 22568 34204 22574
rect 34152 22510 34204 22516
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 32404 22092 32456 22098
rect 32404 22034 32456 22040
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33060 21690 33088 22034
rect 34072 21894 34100 22510
rect 34164 22166 34192 22510
rect 34808 22506 34836 22714
rect 35256 22568 35308 22574
rect 35256 22510 35308 22516
rect 34796 22500 34848 22506
rect 34796 22442 34848 22448
rect 34152 22160 34204 22166
rect 34152 22102 34204 22108
rect 34808 22094 34836 22442
rect 35268 22166 35296 22510
rect 35532 22432 35584 22438
rect 35532 22374 35584 22380
rect 35256 22160 35308 22166
rect 35256 22102 35308 22108
rect 34808 22066 34928 22094
rect 34900 21894 34928 22066
rect 34060 21888 34112 21894
rect 34060 21830 34112 21836
rect 34888 21888 34940 21894
rect 34888 21830 34940 21836
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 34072 21146 34100 21830
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 34060 21140 34112 21146
rect 34060 21082 34112 21088
rect 32680 20800 32732 20806
rect 32680 20742 32732 20748
rect 32692 20398 32720 20742
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 32956 20392 33008 20398
rect 32956 20334 33008 20340
rect 31944 18828 31996 18834
rect 31944 18770 31996 18776
rect 31576 17128 31628 17134
rect 31576 17070 31628 17076
rect 31484 16652 31536 16658
rect 31484 16594 31536 16600
rect 31496 15094 31524 16594
rect 31588 16250 31616 17070
rect 31852 17060 31904 17066
rect 31852 17002 31904 17008
rect 31864 16658 31892 17002
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31956 15638 31984 18770
rect 32600 18698 32628 20334
rect 32968 20058 32996 20334
rect 32956 20052 33008 20058
rect 32956 19994 33008 20000
rect 33336 19922 33364 21082
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 33600 20800 33652 20806
rect 33600 20742 33652 20748
rect 33508 20460 33560 20466
rect 33508 20402 33560 20408
rect 33520 19922 33548 20402
rect 33324 19916 33376 19922
rect 33324 19858 33376 19864
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33612 19854 33640 20742
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33600 19848 33652 19854
rect 33520 19796 33600 19802
rect 33520 19790 33652 19796
rect 33520 19774 33640 19790
rect 32680 19712 32732 19718
rect 32680 19654 32732 19660
rect 32692 19514 32720 19654
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 33520 18766 33548 19774
rect 33888 19446 33916 20402
rect 33876 19440 33928 19446
rect 33876 19382 33928 19388
rect 33600 19168 33652 19174
rect 33600 19110 33652 19116
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 32588 18692 32640 18698
rect 32588 18634 32640 18640
rect 33612 18290 33640 19110
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33048 17672 33100 17678
rect 33048 17614 33100 17620
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32692 16794 32720 16934
rect 33060 16794 33088 17614
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 33152 17202 33180 17478
rect 33796 17338 33824 17614
rect 33784 17332 33836 17338
rect 33784 17274 33836 17280
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 33888 16794 33916 19382
rect 34164 19378 34192 20878
rect 34796 19916 34848 19922
rect 34796 19858 34848 19864
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34532 18834 34560 19790
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34532 18426 34560 18770
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34520 18420 34572 18426
rect 34520 18362 34572 18368
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34244 17128 34296 17134
rect 34244 17070 34296 17076
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34060 16992 34112 16998
rect 34060 16934 34112 16940
rect 32680 16788 32732 16794
rect 32680 16730 32732 16736
rect 33048 16788 33100 16794
rect 33048 16730 33100 16736
rect 33876 16788 33928 16794
rect 33876 16730 33928 16736
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 32048 16250 32076 16526
rect 32036 16244 32088 16250
rect 32036 16186 32088 16192
rect 31944 15632 31996 15638
rect 31944 15574 31996 15580
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31496 13530 31524 14758
rect 32048 13870 32076 16186
rect 32312 15156 32364 15162
rect 32312 15098 32364 15104
rect 32128 14000 32180 14006
rect 32128 13942 32180 13948
rect 32036 13864 32088 13870
rect 32036 13806 32088 13812
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 32048 12986 32076 13806
rect 32140 13190 32168 13942
rect 32128 13184 32180 13190
rect 32128 13126 32180 13132
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31116 12708 31168 12714
rect 31116 12650 31168 12656
rect 31312 12434 31340 12718
rect 31128 12406 31340 12434
rect 31128 12102 31156 12406
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 31024 11552 31076 11558
rect 31024 11494 31076 11500
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 30484 9042 30512 11018
rect 30760 10742 30788 11154
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30852 10062 30880 11494
rect 31036 11082 31064 11494
rect 31024 11076 31076 11082
rect 31024 11018 31076 11024
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30944 10266 30972 10610
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30484 8514 30512 8978
rect 30484 8486 30604 8514
rect 30472 8356 30524 8362
rect 30472 8298 30524 8304
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30300 7478 30328 8230
rect 30484 7886 30512 8298
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30576 7750 30604 8486
rect 30656 8424 30708 8430
rect 30656 8366 30708 8372
rect 30668 8090 30696 8366
rect 30932 8288 30984 8294
rect 30932 8230 30984 8236
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 30748 8016 30800 8022
rect 30748 7958 30800 7964
rect 30760 7750 30788 7958
rect 30944 7818 30972 8230
rect 30932 7812 30984 7818
rect 30932 7754 30984 7760
rect 30564 7744 30616 7750
rect 30748 7744 30800 7750
rect 30616 7704 30696 7732
rect 30564 7686 30616 7692
rect 30288 7472 30340 7478
rect 30288 7414 30340 7420
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30300 4554 30328 4966
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 30300 4282 30328 4490
rect 30392 4282 30420 4558
rect 30288 4276 30340 4282
rect 30288 4218 30340 4224
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30484 4162 30512 6258
rect 30576 5914 30604 6598
rect 30668 6458 30696 7704
rect 30748 7686 30800 7692
rect 30656 6452 30708 6458
rect 30656 6394 30708 6400
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30668 5642 30696 6394
rect 31128 5846 31156 12038
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31588 10266 31616 11630
rect 31680 11218 31708 11766
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 31680 9042 31708 11154
rect 32048 10146 32076 12922
rect 32128 11620 32180 11626
rect 32128 11562 32180 11568
rect 32140 10674 32168 11562
rect 32220 11008 32272 11014
rect 32220 10950 32272 10956
rect 32128 10668 32180 10674
rect 32128 10610 32180 10616
rect 31944 10124 31996 10130
rect 32048 10118 32168 10146
rect 31944 10066 31996 10072
rect 31956 9722 31984 10066
rect 32140 10062 32168 10118
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32140 9722 32168 9998
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 32128 9716 32180 9722
rect 32128 9658 32180 9664
rect 31668 9036 31720 9042
rect 31668 8978 31720 8984
rect 31956 8906 31984 9658
rect 32232 9586 32260 10950
rect 32220 9580 32272 9586
rect 32220 9522 32272 9528
rect 31944 8900 31996 8906
rect 31944 8842 31996 8848
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31404 7546 31432 8366
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31312 6798 31340 7142
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31208 6316 31260 6322
rect 31208 6258 31260 6264
rect 31220 5914 31248 6258
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31116 5840 31168 5846
rect 31116 5782 31168 5788
rect 30656 5636 30708 5642
rect 30656 5578 30708 5584
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30484 4134 30604 4162
rect 30668 4146 30696 4966
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31404 4554 31432 4762
rect 31392 4548 31444 4554
rect 31392 4490 31444 4496
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 30472 4072 30524 4078
rect 30472 4014 30524 4020
rect 30380 4004 30432 4010
rect 30380 3946 30432 3952
rect 30194 3496 30250 3505
rect 30392 3466 30420 3946
rect 30194 3431 30250 3440
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 29838 3292 30146 3301
rect 29838 3290 29844 3292
rect 29900 3290 29924 3292
rect 29980 3290 30004 3292
rect 30060 3290 30084 3292
rect 30140 3290 30146 3292
rect 29900 3238 29902 3290
rect 30082 3238 30084 3290
rect 29838 3236 29844 3238
rect 29900 3236 29924 3238
rect 29980 3236 30004 3238
rect 30060 3236 30084 3238
rect 30140 3236 30146 3238
rect 29838 3227 30146 3236
rect 30484 2774 30512 4014
rect 30576 2990 30604 4134
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30668 3194 30696 3878
rect 30760 3738 30788 3878
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30840 3460 30892 3466
rect 30840 3402 30892 3408
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30564 2984 30616 2990
rect 30564 2926 30616 2932
rect 29380 2746 29500 2774
rect 30392 2746 30512 2774
rect 29380 2650 29408 2746
rect 30392 2650 30420 2746
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30852 2446 30880 3402
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30944 2650 30972 2994
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31128 2514 31156 4422
rect 31496 3602 31524 6734
rect 31680 6662 31708 8774
rect 31944 8356 31996 8362
rect 31944 8298 31996 8304
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 31772 6254 31800 7890
rect 31956 7886 31984 8298
rect 32324 7954 32352 15098
rect 32404 14476 32456 14482
rect 32404 14418 32456 14424
rect 32416 13462 32444 14418
rect 32692 14414 32720 16594
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 33152 14890 33180 15846
rect 33140 14884 33192 14890
rect 33140 14826 33192 14832
rect 32772 14816 32824 14822
rect 32772 14758 32824 14764
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 32680 14408 32732 14414
rect 32680 14350 32732 14356
rect 32496 14272 32548 14278
rect 32496 14214 32548 14220
rect 32508 14074 32536 14214
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32404 13456 32456 13462
rect 32404 13398 32456 13404
rect 32680 13252 32732 13258
rect 32680 13194 32732 13200
rect 32692 12646 32720 13194
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 32692 11626 32720 12582
rect 32680 11620 32732 11626
rect 32680 11562 32732 11568
rect 32784 11234 32812 14758
rect 33244 14346 33272 14758
rect 33232 14340 33284 14346
rect 33232 14282 33284 14288
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32876 12986 32904 13194
rect 32956 13184 33008 13190
rect 32956 13126 33008 13132
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32692 11206 32812 11234
rect 32416 10130 32444 11154
rect 32692 10198 32720 11206
rect 32680 10192 32732 10198
rect 32680 10134 32732 10140
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 32968 10010 32996 13126
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33060 10742 33088 11494
rect 33048 10736 33100 10742
rect 33048 10678 33100 10684
rect 32968 9982 33088 10010
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32680 9512 32732 9518
rect 32680 9454 32732 9460
rect 32692 9178 32720 9454
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32968 8974 32996 9862
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 33060 8566 33088 9982
rect 33244 9042 33272 14282
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33520 14074 33548 14214
rect 33612 14074 33640 14758
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33416 14068 33468 14074
rect 33416 14010 33468 14016
rect 33508 14068 33560 14074
rect 33508 14010 33560 14016
rect 33600 14068 33652 14074
rect 33600 14010 33652 14016
rect 33428 13716 33456 14010
rect 33600 13728 33652 13734
rect 33428 13688 33600 13716
rect 33600 13670 33652 13676
rect 33796 12986 33824 14214
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 33968 12980 34020 12986
rect 33968 12922 34020 12928
rect 33980 12782 34008 12922
rect 33968 12776 34020 12782
rect 33968 12718 34020 12724
rect 33600 11688 33652 11694
rect 33600 11630 33652 11636
rect 33784 11688 33836 11694
rect 33784 11630 33836 11636
rect 33508 11076 33560 11082
rect 33508 11018 33560 11024
rect 33520 9654 33548 11018
rect 33612 10810 33640 11630
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33796 10606 33824 11630
rect 33980 10826 34008 12718
rect 34072 11082 34100 16934
rect 34256 16697 34284 17070
rect 34348 16794 34376 17070
rect 34336 16788 34388 16794
rect 34336 16730 34388 16736
rect 34242 16688 34298 16697
rect 34242 16623 34298 16632
rect 34348 13274 34376 16730
rect 34440 16590 34468 17478
rect 34716 17338 34744 18566
rect 34704 17332 34756 17338
rect 34704 17274 34756 17280
rect 34808 17066 34836 19858
rect 34900 19718 34928 21830
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34900 18630 34928 19654
rect 35072 19168 35124 19174
rect 35072 19110 35124 19116
rect 35084 18834 35112 19110
rect 35072 18828 35124 18834
rect 35072 18770 35124 18776
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34796 17060 34848 17066
rect 34796 17002 34848 17008
rect 34704 16992 34756 16998
rect 34704 16934 34756 16940
rect 34428 16584 34480 16590
rect 34428 16526 34480 16532
rect 34716 16182 34744 16934
rect 34704 16176 34756 16182
rect 34704 16118 34756 16124
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34532 14226 34560 15846
rect 34532 14198 34744 14226
rect 34612 13932 34664 13938
rect 34612 13874 34664 13880
rect 34520 13456 34572 13462
rect 34520 13398 34572 13404
rect 34256 13246 34376 13274
rect 34256 12986 34284 13246
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34244 12980 34296 12986
rect 34244 12922 34296 12928
rect 34348 12434 34376 13126
rect 34256 12406 34376 12434
rect 34060 11076 34112 11082
rect 34060 11018 34112 11024
rect 33980 10798 34100 10826
rect 33968 10668 34020 10674
rect 33968 10610 34020 10616
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33980 10130 34008 10610
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33600 9988 33652 9994
rect 33600 9930 33652 9936
rect 33612 9722 33640 9930
rect 33600 9716 33652 9722
rect 33600 9658 33652 9664
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33416 9580 33468 9586
rect 33416 9522 33468 9528
rect 33232 9036 33284 9042
rect 33232 8978 33284 8984
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 33244 8430 33272 8978
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 33232 8424 33284 8430
rect 33232 8366 33284 8372
rect 32680 8288 32732 8294
rect 32680 8230 32732 8236
rect 32312 7948 32364 7954
rect 32312 7890 32364 7896
rect 31944 7880 31996 7886
rect 32692 7857 32720 8230
rect 33232 8016 33284 8022
rect 33336 8004 33364 8910
rect 33428 8838 33456 9522
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33428 8430 33456 8774
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 33284 7976 33364 8004
rect 33232 7958 33284 7964
rect 31944 7822 31996 7828
rect 32678 7848 32734 7857
rect 32312 7812 32364 7818
rect 32678 7783 32734 7792
rect 32312 7754 32364 7760
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 31864 6390 31892 7278
rect 32232 6882 32260 7346
rect 31956 6866 32260 6882
rect 31944 6860 32260 6866
rect 31996 6854 32260 6860
rect 31944 6802 31996 6808
rect 32232 6390 32260 6854
rect 32324 6798 32352 7754
rect 32588 6996 32640 7002
rect 32588 6938 32640 6944
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 31852 6384 31904 6390
rect 31852 6326 31904 6332
rect 32220 6384 32272 6390
rect 32220 6326 32272 6332
rect 32312 6316 32364 6322
rect 32416 6304 32444 6734
rect 32600 6662 32628 6938
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32364 6276 32444 6304
rect 32496 6316 32548 6322
rect 32312 6258 32364 6264
rect 32496 6258 32548 6264
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 32508 5370 32536 6258
rect 32600 5914 32628 6598
rect 32588 5908 32640 5914
rect 32588 5850 32640 5856
rect 33152 5710 33180 6734
rect 33244 5778 33272 7958
rect 33428 7834 33456 8366
rect 33876 8356 33928 8362
rect 33876 8298 33928 8304
rect 33336 7806 33456 7834
rect 33336 6934 33364 7806
rect 33598 7440 33654 7449
rect 33888 7410 33916 8298
rect 33598 7375 33600 7384
rect 33652 7375 33654 7384
rect 33876 7404 33928 7410
rect 33600 7346 33652 7352
rect 33876 7346 33928 7352
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 33324 6928 33376 6934
rect 33376 6876 33456 6882
rect 33324 6870 33456 6876
rect 33336 6854 33456 6870
rect 33324 6792 33376 6798
rect 33324 6734 33376 6740
rect 33336 5778 33364 6734
rect 33232 5772 33284 5778
rect 33232 5714 33284 5720
rect 33324 5772 33376 5778
rect 33324 5714 33376 5720
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33152 5370 33180 5646
rect 33428 5574 33456 6854
rect 33324 5568 33376 5574
rect 33324 5510 33376 5516
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 32496 5364 32548 5370
rect 32496 5306 32548 5312
rect 33140 5364 33192 5370
rect 33140 5306 33192 5312
rect 33336 5234 33364 5510
rect 33520 5234 33548 7142
rect 33612 7002 33640 7346
rect 33692 7336 33744 7342
rect 33692 7278 33744 7284
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33704 6866 33732 7278
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33980 6798 34008 10066
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 33876 6112 33928 6118
rect 33876 6054 33928 6060
rect 33784 5772 33836 5778
rect 33784 5714 33836 5720
rect 33796 5370 33824 5714
rect 33784 5364 33836 5370
rect 33784 5306 33836 5312
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33508 5228 33560 5234
rect 33508 5170 33560 5176
rect 32404 5024 32456 5030
rect 32404 4966 32456 4972
rect 32416 4690 32444 4966
rect 32404 4684 32456 4690
rect 32404 4626 32456 4632
rect 33888 4622 33916 6054
rect 33980 5710 34008 6734
rect 33968 5704 34020 5710
rect 33968 5646 34020 5652
rect 34072 5030 34100 10798
rect 34152 10464 34204 10470
rect 34152 10406 34204 10412
rect 34164 10266 34192 10406
rect 34152 10260 34204 10266
rect 34152 10202 34204 10208
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34256 9874 34284 12406
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34336 11076 34388 11082
rect 34336 11018 34388 11024
rect 34348 10130 34376 11018
rect 34440 10810 34468 11494
rect 34428 10804 34480 10810
rect 34428 10746 34480 10752
rect 34440 10130 34468 10746
rect 34336 10124 34388 10130
rect 34336 10066 34388 10072
rect 34428 10124 34480 10130
rect 34428 10066 34480 10072
rect 34348 10010 34376 10066
rect 34348 9982 34468 10010
rect 34440 9926 34468 9982
rect 34428 9920 34480 9926
rect 34164 9586 34192 9862
rect 34256 9846 34376 9874
rect 34428 9862 34480 9868
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 34348 8974 34376 9846
rect 34440 9178 34468 9862
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34164 6934 34192 8774
rect 34532 8498 34560 13398
rect 34624 13394 34652 13874
rect 34612 13388 34664 13394
rect 34612 13330 34664 13336
rect 34716 9586 34744 14198
rect 34900 11898 34928 18566
rect 35256 16992 35308 16998
rect 35256 16934 35308 16940
rect 35164 13252 35216 13258
rect 35164 13194 35216 13200
rect 35176 12986 35204 13194
rect 35164 12980 35216 12986
rect 35164 12922 35216 12928
rect 34980 12912 35032 12918
rect 34980 12854 35032 12860
rect 34992 12434 35020 12854
rect 34992 12406 35204 12434
rect 34888 11892 34940 11898
rect 34888 11834 34940 11840
rect 35072 11756 35124 11762
rect 35072 11698 35124 11704
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 34808 11218 34836 11630
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 34808 10674 34836 11154
rect 35084 10810 35112 11698
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34808 10062 34836 10610
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34808 9178 34836 9998
rect 34978 9616 35034 9625
rect 34978 9551 34980 9560
rect 35032 9551 35034 9560
rect 34980 9522 35032 9528
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 34612 8900 34664 8906
rect 34612 8842 34664 8848
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 34060 5024 34112 5030
rect 34060 4966 34112 4972
rect 34072 4622 34100 4966
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 34164 4554 34192 4762
rect 34152 4548 34204 4554
rect 34152 4490 34204 4496
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33876 4480 33928 4486
rect 33876 4422 33928 4428
rect 32140 4282 32168 4422
rect 33520 4282 33548 4422
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33508 4276 33560 4282
rect 33508 4218 33560 4224
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 31680 3738 31708 3878
rect 31668 3732 31720 3738
rect 31668 3674 31720 3680
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 31404 3194 31432 3470
rect 32876 3194 32904 3878
rect 31392 3188 31444 3194
rect 31392 3130 31444 3136
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 33428 3058 33456 4218
rect 33888 4214 33916 4422
rect 33968 4276 34020 4282
rect 33968 4218 34020 4224
rect 33876 4208 33928 4214
rect 33876 4150 33928 4156
rect 33508 4140 33560 4146
rect 33508 4082 33560 4088
rect 33520 3738 33548 4082
rect 33508 3732 33560 3738
rect 33508 3674 33560 3680
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33506 3088 33562 3097
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 33416 3052 33468 3058
rect 33468 3032 33506 3040
rect 33468 3023 33562 3032
rect 33468 3012 33548 3023
rect 33416 2994 33468 3000
rect 31220 2774 31248 2994
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 31220 2746 31340 2774
rect 31024 2508 31076 2514
rect 31024 2450 31076 2456
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 29552 2440 29604 2446
rect 30196 2440 30248 2446
rect 29604 2400 29684 2428
rect 29552 2382 29604 2388
rect 29104 1414 29224 1442
rect 29104 800 29132 1414
rect 29656 800 29684 2400
rect 30196 2382 30248 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 29838 2204 30146 2213
rect 29838 2202 29844 2204
rect 29900 2202 29924 2204
rect 29980 2202 30004 2204
rect 30060 2202 30084 2204
rect 30140 2202 30146 2204
rect 29900 2150 29902 2202
rect 30082 2150 30084 2202
rect 29838 2148 29844 2150
rect 29900 2148 29924 2150
rect 29980 2148 30004 2150
rect 30060 2148 30084 2150
rect 30140 2148 30146 2150
rect 29838 2139 30146 2148
rect 30208 800 30236 2382
rect 30760 870 30880 898
rect 30760 800 30788 870
rect 22572 734 22784 762
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 30852 762 30880 870
rect 31036 762 31064 2450
rect 31312 800 31340 2746
rect 31864 800 31892 2926
rect 32956 2916 33008 2922
rect 32956 2858 33008 2864
rect 31944 2848 31996 2854
rect 31944 2790 31996 2796
rect 31956 2632 31984 2790
rect 31956 2604 32168 2632
rect 32140 2446 32168 2604
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 32416 800 32444 2314
rect 32968 800 32996 2858
rect 33152 2650 33180 2926
rect 33612 2774 33640 2926
rect 33520 2746 33640 2774
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33520 800 33548 2746
rect 33704 2446 33732 3334
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33980 2378 34008 4218
rect 34348 3194 34376 8434
rect 34624 6322 34652 8842
rect 34900 8566 34928 8978
rect 34888 8560 34940 8566
rect 34888 8502 34940 8508
rect 34888 7880 34940 7886
rect 34888 7822 34940 7828
rect 34704 6724 34756 6730
rect 34704 6666 34756 6672
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34520 6180 34572 6186
rect 34520 6122 34572 6128
rect 34532 5234 34560 6122
rect 34716 5778 34744 6666
rect 34900 6458 34928 7822
rect 34888 6452 34940 6458
rect 34888 6394 34940 6400
rect 34900 5778 34928 6394
rect 34704 5772 34756 5778
rect 34704 5714 34756 5720
rect 34888 5772 34940 5778
rect 34888 5714 34940 5720
rect 34716 5370 34744 5714
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34520 5228 34572 5234
rect 34520 5170 34572 5176
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 33968 2372 34020 2378
rect 33968 2314 34020 2320
rect 34520 2372 34572 2378
rect 34520 2314 34572 2320
rect 34532 1442 34560 2314
rect 34440 1414 34560 1442
rect 34072 870 34192 898
rect 34072 800 34100 870
rect 30852 734 31064 762
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34164 762 34192 870
rect 34440 762 34468 1414
rect 34624 800 34652 3606
rect 34716 2854 34744 5170
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34808 4214 34836 4966
rect 34900 4826 34928 5170
rect 34888 4820 34940 4826
rect 34888 4762 34940 4768
rect 34992 4622 35020 9522
rect 35176 8362 35204 12406
rect 35268 10146 35296 16934
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 35360 12850 35388 14214
rect 35452 13258 35480 21626
rect 35544 19514 35572 22374
rect 35636 21350 35664 22936
rect 35728 22778 35756 23462
rect 35716 22772 35768 22778
rect 35716 22714 35768 22720
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35820 22094 35848 22646
rect 35728 22066 35848 22094
rect 35728 21690 35756 22066
rect 35808 22024 35860 22030
rect 35912 21978 35940 23462
rect 36004 22506 36032 24142
rect 36820 24064 36872 24070
rect 36820 24006 36872 24012
rect 36636 23316 36688 23322
rect 36636 23258 36688 23264
rect 36176 23044 36228 23050
rect 36176 22986 36228 22992
rect 36084 22976 36136 22982
rect 36084 22918 36136 22924
rect 35992 22500 36044 22506
rect 35992 22442 36044 22448
rect 36096 22098 36124 22918
rect 36188 22778 36216 22986
rect 36176 22772 36228 22778
rect 36176 22714 36228 22720
rect 36648 22166 36676 23258
rect 36832 23050 36860 24006
rect 37568 23866 37596 24142
rect 37556 23860 37608 23866
rect 37556 23802 37608 23808
rect 37648 23656 37700 23662
rect 37648 23598 37700 23604
rect 37060 23420 37368 23429
rect 37060 23418 37066 23420
rect 37122 23418 37146 23420
rect 37202 23418 37226 23420
rect 37282 23418 37306 23420
rect 37362 23418 37368 23420
rect 37122 23366 37124 23418
rect 37304 23366 37306 23418
rect 37060 23364 37066 23366
rect 37122 23364 37146 23366
rect 37202 23364 37226 23366
rect 37282 23364 37306 23366
rect 37362 23364 37368 23366
rect 37060 23355 37368 23364
rect 36912 23112 36964 23118
rect 36912 23054 36964 23060
rect 36820 23044 36872 23050
rect 36820 22986 36872 22992
rect 36924 22574 36952 23054
rect 36728 22568 36780 22574
rect 36728 22510 36780 22516
rect 36912 22568 36964 22574
rect 36912 22510 36964 22516
rect 36636 22160 36688 22166
rect 36636 22102 36688 22108
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 35860 21972 35940 21978
rect 35808 21966 35940 21972
rect 35820 21950 35940 21966
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35636 19990 35664 21286
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 35716 20256 35768 20262
rect 35716 20198 35768 20204
rect 35624 19984 35676 19990
rect 35624 19926 35676 19932
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35728 19310 35756 20198
rect 35820 20058 35848 20334
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35820 19514 35848 19858
rect 35808 19508 35860 19514
rect 35808 19450 35860 19456
rect 35624 19304 35676 19310
rect 35624 19246 35676 19252
rect 35716 19304 35768 19310
rect 35716 19246 35768 19252
rect 35532 19236 35584 19242
rect 35532 19178 35584 19184
rect 35544 14618 35572 19178
rect 35636 18630 35664 19246
rect 35624 18624 35676 18630
rect 35624 18566 35676 18572
rect 35636 14958 35664 18566
rect 35820 18426 35848 19450
rect 35808 18420 35860 18426
rect 35808 18362 35860 18368
rect 35716 17536 35768 17542
rect 35716 17478 35768 17484
rect 35728 16522 35756 17478
rect 35808 17264 35860 17270
rect 35808 17206 35860 17212
rect 35820 16522 35848 17206
rect 35912 16998 35940 21950
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 36004 20058 36032 20198
rect 35992 20052 36044 20058
rect 35992 19994 36044 20000
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 36188 19378 36216 19790
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 36096 18902 36124 19246
rect 36084 18896 36136 18902
rect 36084 18838 36136 18844
rect 36188 18834 36216 19314
rect 36452 19304 36504 19310
rect 36452 19246 36504 19252
rect 36464 18970 36492 19246
rect 36452 18964 36504 18970
rect 36452 18906 36504 18912
rect 36176 18828 36228 18834
rect 36176 18770 36228 18776
rect 36648 17762 36676 22102
rect 36740 21894 36768 22510
rect 36924 22094 36952 22510
rect 37060 22332 37368 22341
rect 37060 22330 37066 22332
rect 37122 22330 37146 22332
rect 37202 22330 37226 22332
rect 37282 22330 37306 22332
rect 37362 22330 37368 22332
rect 37122 22278 37124 22330
rect 37304 22278 37306 22330
rect 37060 22276 37066 22278
rect 37122 22276 37146 22278
rect 37202 22276 37226 22278
rect 37282 22276 37306 22278
rect 37362 22276 37368 22278
rect 37060 22267 37368 22276
rect 36832 22066 36952 22094
rect 36728 21888 36780 21894
rect 36728 21830 36780 21836
rect 36728 21480 36780 21486
rect 36728 21422 36780 21428
rect 36740 21010 36768 21422
rect 36832 21026 36860 22066
rect 37660 21894 37688 23598
rect 37752 23322 37780 24142
rect 38396 23730 38424 25298
rect 42628 24818 42748 24834
rect 42628 24812 42760 24818
rect 42628 24806 42708 24812
rect 42248 24608 42300 24614
rect 42248 24550 42300 24556
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 41144 24200 41196 24206
rect 41144 24142 41196 24148
rect 38936 24064 38988 24070
rect 38936 24006 38988 24012
rect 39672 24064 39724 24070
rect 39672 24006 39724 24012
rect 39856 24064 39908 24070
rect 39856 24006 39908 24012
rect 38948 23866 38976 24006
rect 38936 23860 38988 23866
rect 38936 23802 38988 23808
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38384 23724 38436 23730
rect 38384 23666 38436 23672
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38304 23322 38332 23666
rect 38580 23474 38608 23666
rect 38580 23446 38700 23474
rect 37740 23316 37792 23322
rect 37740 23258 37792 23264
rect 38292 23316 38344 23322
rect 38292 23258 38344 23264
rect 38292 23180 38344 23186
rect 38292 23122 38344 23128
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 38028 22166 38056 22578
rect 38016 22160 38068 22166
rect 38016 22102 38068 22108
rect 37648 21888 37700 21894
rect 37648 21830 37700 21836
rect 37060 21244 37368 21253
rect 37060 21242 37066 21244
rect 37122 21242 37146 21244
rect 37202 21242 37226 21244
rect 37282 21242 37306 21244
rect 37362 21242 37368 21244
rect 37122 21190 37124 21242
rect 37304 21190 37306 21242
rect 37060 21188 37066 21190
rect 37122 21188 37146 21190
rect 37202 21188 37226 21190
rect 37282 21188 37306 21190
rect 37362 21188 37368 21190
rect 37060 21179 37368 21188
rect 36728 21004 36780 21010
rect 36832 20998 36952 21026
rect 36728 20946 36780 20952
rect 36728 20868 36780 20874
rect 36728 20810 36780 20816
rect 36740 19786 36768 20810
rect 36924 20806 36952 20998
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 36912 20800 36964 20806
rect 36912 20742 36964 20748
rect 36924 20330 36952 20742
rect 37464 20392 37516 20398
rect 37464 20334 37516 20340
rect 36912 20324 36964 20330
rect 36912 20266 36964 20272
rect 36924 19854 36952 20266
rect 37060 20156 37368 20165
rect 37060 20154 37066 20156
rect 37122 20154 37146 20156
rect 37202 20154 37226 20156
rect 37282 20154 37306 20156
rect 37362 20154 37368 20156
rect 37122 20102 37124 20154
rect 37304 20102 37306 20154
rect 37060 20100 37066 20102
rect 37122 20100 37146 20102
rect 37202 20100 37226 20102
rect 37282 20100 37306 20102
rect 37362 20100 37368 20102
rect 37060 20091 37368 20100
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36728 19780 36780 19786
rect 36728 19722 36780 19728
rect 37476 19378 37504 20334
rect 37568 19514 37596 20878
rect 37660 20466 37688 21830
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37844 21010 37872 21286
rect 38304 21078 38332 23122
rect 38672 22642 38700 23446
rect 38948 23186 38976 23802
rect 39684 23662 39712 24006
rect 39868 23866 39896 24006
rect 39856 23860 39908 23866
rect 39856 23802 39908 23808
rect 40224 23724 40276 23730
rect 40224 23666 40276 23672
rect 40316 23724 40368 23730
rect 40316 23666 40368 23672
rect 39672 23656 39724 23662
rect 39672 23598 39724 23604
rect 39028 23248 39080 23254
rect 39028 23190 39080 23196
rect 38936 23180 38988 23186
rect 38936 23122 38988 23128
rect 38752 23112 38804 23118
rect 38752 23054 38804 23060
rect 38660 22636 38712 22642
rect 38660 22578 38712 22584
rect 38660 22432 38712 22438
rect 38660 22374 38712 22380
rect 38672 22098 38700 22374
rect 38764 22166 38792 23054
rect 38752 22160 38804 22166
rect 38752 22102 38804 22108
rect 38660 22092 38712 22098
rect 38660 22034 38712 22040
rect 38292 21072 38344 21078
rect 38292 21014 38344 21020
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37648 20460 37700 20466
rect 37648 20402 37700 20408
rect 37752 20058 37780 20878
rect 37844 20398 37872 20946
rect 38108 20596 38160 20602
rect 38108 20538 38160 20544
rect 38120 20398 38148 20538
rect 37832 20392 37884 20398
rect 37832 20334 37884 20340
rect 38108 20392 38160 20398
rect 38108 20334 38160 20340
rect 37832 20256 37884 20262
rect 37832 20198 37884 20204
rect 38016 20256 38068 20262
rect 38016 20198 38068 20204
rect 37740 20052 37792 20058
rect 37740 19994 37792 20000
rect 37556 19508 37608 19514
rect 37556 19450 37608 19456
rect 37844 19446 37872 20198
rect 37832 19440 37884 19446
rect 37832 19382 37884 19388
rect 37464 19372 37516 19378
rect 37464 19314 37516 19320
rect 37060 19068 37368 19077
rect 37060 19066 37066 19068
rect 37122 19066 37146 19068
rect 37202 19066 37226 19068
rect 37282 19066 37306 19068
rect 37362 19066 37368 19068
rect 37122 19014 37124 19066
rect 37304 19014 37306 19066
rect 37060 19012 37066 19014
rect 37122 19012 37146 19014
rect 37202 19012 37226 19014
rect 37282 19012 37306 19014
rect 37362 19012 37368 19014
rect 37060 19003 37368 19012
rect 37476 18170 37504 19314
rect 37476 18142 37688 18170
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 37060 17980 37368 17989
rect 37060 17978 37066 17980
rect 37122 17978 37146 17980
rect 37202 17978 37226 17980
rect 37282 17978 37306 17980
rect 37362 17978 37368 17980
rect 37122 17926 37124 17978
rect 37304 17926 37306 17978
rect 37060 17924 37066 17926
rect 37122 17924 37146 17926
rect 37202 17924 37226 17926
rect 37282 17924 37306 17926
rect 37362 17924 37368 17926
rect 37060 17915 37368 17924
rect 37568 17814 37596 18022
rect 37556 17808 37608 17814
rect 36648 17734 36768 17762
rect 37556 17750 37608 17756
rect 36360 17672 36412 17678
rect 36360 17614 36412 17620
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 36372 17338 36400 17614
rect 36360 17332 36412 17338
rect 36360 17274 36412 17280
rect 36452 17128 36504 17134
rect 36280 17076 36452 17082
rect 36280 17070 36504 17076
rect 36280 17054 36492 17070
rect 36280 16998 36308 17054
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 36268 16992 36320 16998
rect 36268 16934 36320 16940
rect 36648 16794 36676 17614
rect 36740 17338 36768 17734
rect 37188 17604 37240 17610
rect 37188 17546 37240 17552
rect 36728 17332 36780 17338
rect 36728 17274 36780 17280
rect 36636 16788 36688 16794
rect 36636 16730 36688 16736
rect 36740 16658 36768 17274
rect 37200 17202 37228 17546
rect 37372 17536 37424 17542
rect 37372 17478 37424 17484
rect 37384 17202 37412 17478
rect 37188 17196 37240 17202
rect 37188 17138 37240 17144
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37464 16992 37516 16998
rect 37464 16934 37516 16940
rect 37060 16892 37368 16901
rect 37060 16890 37066 16892
rect 37122 16890 37146 16892
rect 37202 16890 37226 16892
rect 37282 16890 37306 16892
rect 37362 16890 37368 16892
rect 37122 16838 37124 16890
rect 37304 16838 37306 16890
rect 37060 16836 37066 16838
rect 37122 16836 37146 16838
rect 37202 16836 37226 16838
rect 37282 16836 37306 16838
rect 37362 16836 37368 16838
rect 37060 16827 37368 16836
rect 37476 16658 37504 16934
rect 37568 16794 37596 17750
rect 37556 16788 37608 16794
rect 37556 16730 37608 16736
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 35716 16516 35768 16522
rect 35716 16458 35768 16464
rect 35808 16516 35860 16522
rect 35808 16458 35860 16464
rect 35820 16114 35848 16458
rect 35808 16108 35860 16114
rect 35808 16050 35860 16056
rect 36740 15162 36768 16594
rect 37060 15804 37368 15813
rect 37060 15802 37066 15804
rect 37122 15802 37146 15804
rect 37202 15802 37226 15804
rect 37282 15802 37306 15804
rect 37362 15802 37368 15804
rect 37122 15750 37124 15802
rect 37304 15750 37306 15802
rect 37060 15748 37066 15750
rect 37122 15748 37146 15750
rect 37202 15748 37226 15750
rect 37282 15748 37306 15750
rect 37362 15748 37368 15750
rect 37060 15739 37368 15748
rect 36728 15156 36780 15162
rect 36728 15098 36780 15104
rect 36544 15088 36596 15094
rect 36544 15030 36596 15036
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35992 14952 36044 14958
rect 35992 14894 36044 14900
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 35544 12434 35572 14554
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 35912 14074 35940 14214
rect 36004 14074 36032 14894
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 36556 13870 36584 15030
rect 37060 14716 37368 14725
rect 37060 14714 37066 14716
rect 37122 14714 37146 14716
rect 37202 14714 37226 14716
rect 37282 14714 37306 14716
rect 37362 14714 37368 14716
rect 37122 14662 37124 14714
rect 37304 14662 37306 14714
rect 37060 14660 37066 14662
rect 37122 14660 37146 14662
rect 37202 14660 37226 14662
rect 37282 14660 37306 14662
rect 37362 14660 37368 14662
rect 37060 14651 37368 14660
rect 37476 14414 37504 16594
rect 37660 16538 37688 18142
rect 37568 16510 37688 16538
rect 37568 15162 37596 16510
rect 37648 16448 37700 16454
rect 37648 16390 37700 16396
rect 37660 16250 37688 16390
rect 37648 16244 37700 16250
rect 37648 16186 37700 16192
rect 37844 15502 37872 19382
rect 38028 18834 38056 20198
rect 38016 18828 38068 18834
rect 38016 18770 38068 18776
rect 38120 18766 38148 20334
rect 38304 19938 38332 21014
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 38384 20800 38436 20806
rect 38384 20742 38436 20748
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 38212 19922 38332 19938
rect 38200 19916 38332 19922
rect 38252 19910 38332 19916
rect 38200 19858 38252 19864
rect 38304 19174 38332 19910
rect 38396 19836 38424 20742
rect 38764 20602 38792 20742
rect 38948 20602 38976 20878
rect 38752 20596 38804 20602
rect 38752 20538 38804 20544
rect 38936 20596 38988 20602
rect 38936 20538 38988 20544
rect 38660 20528 38712 20534
rect 38660 20470 38712 20476
rect 38568 20460 38620 20466
rect 38568 20402 38620 20408
rect 38476 19848 38528 19854
rect 38396 19808 38476 19836
rect 38396 19514 38424 19808
rect 38476 19790 38528 19796
rect 38580 19666 38608 20402
rect 38672 19922 38700 20470
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38856 20058 38884 20334
rect 38844 20052 38896 20058
rect 38844 19994 38896 20000
rect 39040 19922 39068 23190
rect 40236 23050 40264 23666
rect 40328 23186 40356 23666
rect 40420 23322 40448 24142
rect 40592 24064 40644 24070
rect 40592 24006 40644 24012
rect 40408 23316 40460 23322
rect 40408 23258 40460 23264
rect 40316 23180 40368 23186
rect 40316 23122 40368 23128
rect 40408 23180 40460 23186
rect 40408 23122 40460 23128
rect 40224 23044 40276 23050
rect 40224 22986 40276 22992
rect 40420 22982 40448 23122
rect 40040 22976 40092 22982
rect 40040 22918 40092 22924
rect 40408 22976 40460 22982
rect 40408 22918 40460 22924
rect 39580 20800 39632 20806
rect 39580 20742 39632 20748
rect 39120 20256 39172 20262
rect 39120 20198 39172 20204
rect 39132 20058 39160 20198
rect 39120 20052 39172 20058
rect 39120 19994 39172 20000
rect 38660 19916 38712 19922
rect 38660 19858 38712 19864
rect 39028 19916 39080 19922
rect 39028 19858 39080 19864
rect 38488 19638 38608 19666
rect 38384 19508 38436 19514
rect 38384 19450 38436 19456
rect 38488 19378 38516 19638
rect 38476 19372 38528 19378
rect 38476 19314 38528 19320
rect 38292 19168 38344 19174
rect 38292 19110 38344 19116
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37556 15156 37608 15162
rect 37556 15098 37608 15104
rect 37740 14816 37792 14822
rect 37740 14758 37792 14764
rect 37752 14618 37780 14758
rect 37740 14612 37792 14618
rect 37740 14554 37792 14560
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 36636 14340 36688 14346
rect 36636 14282 36688 14288
rect 36544 13864 36596 13870
rect 36544 13806 36596 13812
rect 36648 13818 36676 14282
rect 36740 14074 36768 14350
rect 36728 14068 36780 14074
rect 36728 14010 36780 14016
rect 37292 13954 37320 14350
rect 37648 14340 37700 14346
rect 37648 14282 37700 14288
rect 37372 14272 37424 14278
rect 37372 14214 37424 14220
rect 37200 13938 37320 13954
rect 37384 13938 37412 14214
rect 37660 13938 37688 14282
rect 37188 13932 37320 13938
rect 37240 13926 37320 13932
rect 37372 13932 37424 13938
rect 37188 13874 37240 13880
rect 37372 13874 37424 13880
rect 37648 13932 37700 13938
rect 37648 13874 37700 13880
rect 36728 13864 36780 13870
rect 36648 13812 36728 13818
rect 36648 13806 36780 13812
rect 37384 13818 37412 13874
rect 37752 13818 37780 14554
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35820 12986 35848 13262
rect 36084 13184 36136 13190
rect 36084 13126 36136 13132
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 36096 12918 36124 13126
rect 36084 12912 36136 12918
rect 36084 12854 36136 12860
rect 35452 12406 35572 12434
rect 35452 11830 35480 12406
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 35440 11824 35492 11830
rect 35440 11766 35492 11772
rect 35452 11218 35480 11766
rect 36096 11694 36124 12038
rect 36084 11688 36136 11694
rect 36084 11630 36136 11636
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 36360 11688 36412 11694
rect 36360 11630 36412 11636
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35532 11280 35584 11286
rect 35532 11222 35584 11228
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35268 10118 35388 10146
rect 35256 9988 35308 9994
rect 35256 9930 35308 9936
rect 35268 9722 35296 9930
rect 35256 9716 35308 9722
rect 35256 9658 35308 9664
rect 35360 9674 35388 10118
rect 35360 9646 35480 9674
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35164 8356 35216 8362
rect 35164 8298 35216 8304
rect 35072 7336 35124 7342
rect 35072 7278 35124 7284
rect 35084 6934 35112 7278
rect 35072 6928 35124 6934
rect 35072 6870 35124 6876
rect 35084 5846 35112 6870
rect 35072 5840 35124 5846
rect 35072 5782 35124 5788
rect 34980 4616 35032 4622
rect 34980 4558 35032 4564
rect 35072 4276 35124 4282
rect 35072 4218 35124 4224
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 34794 4040 34850 4049
rect 34794 3975 34850 3984
rect 34808 3194 34836 3975
rect 34888 3460 34940 3466
rect 34888 3402 34940 3408
rect 34900 3194 34928 3402
rect 34796 3188 34848 3194
rect 34796 3130 34848 3136
rect 34888 3188 34940 3194
rect 34888 3130 34940 3136
rect 35084 2990 35112 4218
rect 35176 3466 35204 8298
rect 35268 7818 35296 8774
rect 35452 8430 35480 9646
rect 35544 9586 35572 11222
rect 35636 10742 35664 11494
rect 36096 11150 36124 11630
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35820 10826 35848 10950
rect 35820 10810 35940 10826
rect 35716 10804 35768 10810
rect 35716 10746 35768 10752
rect 35820 10804 35952 10810
rect 35820 10798 35900 10804
rect 35624 10736 35676 10742
rect 35624 10678 35676 10684
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35452 8090 35480 8366
rect 35440 8084 35492 8090
rect 35440 8026 35492 8032
rect 35256 7812 35308 7818
rect 35256 7754 35308 7760
rect 35256 6792 35308 6798
rect 35256 6734 35308 6740
rect 35268 5914 35296 6734
rect 35256 5908 35308 5914
rect 35256 5850 35308 5856
rect 35624 3936 35676 3942
rect 35624 3878 35676 3884
rect 35636 3466 35664 3878
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35624 3460 35676 3466
rect 35624 3402 35676 3408
rect 35348 3392 35400 3398
rect 35348 3334 35400 3340
rect 35360 3194 35388 3334
rect 35348 3188 35400 3194
rect 35348 3130 35400 3136
rect 35072 2984 35124 2990
rect 35072 2926 35124 2932
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 35084 2514 35112 2926
rect 35268 2774 35296 2926
rect 35176 2746 35296 2774
rect 35072 2508 35124 2514
rect 35072 2450 35124 2456
rect 35176 800 35204 2746
rect 35636 2582 35664 3402
rect 35728 3194 35756 10746
rect 35820 8566 35848 10798
rect 35900 10746 35952 10752
rect 36004 10130 36032 11018
rect 36188 10810 36216 11630
rect 36176 10804 36228 10810
rect 36176 10746 36228 10752
rect 36372 10606 36400 11630
rect 36556 10606 36584 13806
rect 36648 13790 36768 13806
rect 37384 13790 37596 13818
rect 36648 12918 36676 13790
rect 37060 13628 37368 13637
rect 37060 13626 37066 13628
rect 37122 13626 37146 13628
rect 37202 13626 37226 13628
rect 37282 13626 37306 13628
rect 37362 13626 37368 13628
rect 37122 13574 37124 13626
rect 37304 13574 37306 13626
rect 37060 13572 37066 13574
rect 37122 13572 37146 13574
rect 37202 13572 37226 13574
rect 37282 13572 37306 13574
rect 37362 13572 37368 13574
rect 37060 13563 37368 13572
rect 37568 12918 37596 13790
rect 37660 13790 37780 13818
rect 37844 13802 37872 15438
rect 38120 14890 38148 18702
rect 38304 16658 38332 19110
rect 38384 17536 38436 17542
rect 38384 17478 38436 17484
rect 38292 16652 38344 16658
rect 38292 16594 38344 16600
rect 38304 15366 38332 16594
rect 38292 15360 38344 15366
rect 38292 15302 38344 15308
rect 38108 14884 38160 14890
rect 38108 14826 38160 14832
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 37832 13796 37884 13802
rect 36636 12912 36688 12918
rect 36636 12854 36688 12860
rect 37556 12912 37608 12918
rect 37556 12854 37608 12860
rect 37060 12540 37368 12549
rect 37060 12538 37066 12540
rect 37122 12538 37146 12540
rect 37202 12538 37226 12540
rect 37282 12538 37306 12540
rect 37362 12538 37368 12540
rect 37122 12486 37124 12538
rect 37304 12486 37306 12538
rect 37060 12484 37066 12486
rect 37122 12484 37146 12486
rect 37202 12484 37226 12486
rect 37282 12484 37306 12486
rect 37362 12484 37368 12486
rect 37060 12475 37368 12484
rect 37660 12238 37688 13790
rect 37832 13738 37884 13744
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37752 12918 37780 13126
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 37844 12434 37872 13738
rect 37936 13190 37964 14214
rect 38212 14074 38240 14758
rect 38304 14278 38332 15302
rect 38292 14272 38344 14278
rect 38292 14214 38344 14220
rect 38200 14068 38252 14074
rect 38200 14010 38252 14016
rect 38212 13938 38240 14010
rect 38200 13932 38252 13938
rect 38200 13874 38252 13880
rect 37924 13184 37976 13190
rect 37924 13126 37976 13132
rect 37844 12406 37964 12434
rect 37648 12232 37700 12238
rect 37648 12174 37700 12180
rect 36912 12096 36964 12102
rect 36912 12038 36964 12044
rect 36820 11620 36872 11626
rect 36820 11562 36872 11568
rect 36636 11552 36688 11558
rect 36636 11494 36688 11500
rect 36648 10810 36676 11494
rect 36832 11082 36860 11562
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36544 10600 36596 10606
rect 36544 10542 36596 10548
rect 36556 10266 36584 10542
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 35992 10124 36044 10130
rect 35992 10066 36044 10072
rect 36004 9722 36032 10066
rect 36084 9920 36136 9926
rect 36084 9862 36136 9868
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 35992 9716 36044 9722
rect 35992 9658 36044 9664
rect 36096 9586 36124 9862
rect 36084 9580 36136 9586
rect 36084 9522 36136 9528
rect 35992 9036 36044 9042
rect 35992 8978 36044 8984
rect 36004 8566 36032 8978
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36188 8090 36216 8502
rect 36176 8084 36228 8090
rect 36176 8026 36228 8032
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 36188 7342 36216 7686
rect 36280 7546 36308 9862
rect 36556 9178 36584 10202
rect 36648 10033 36676 10746
rect 36924 10146 36952 12038
rect 37060 11452 37368 11461
rect 37060 11450 37066 11452
rect 37122 11450 37146 11452
rect 37202 11450 37226 11452
rect 37282 11450 37306 11452
rect 37362 11450 37368 11452
rect 37122 11398 37124 11450
rect 37304 11398 37306 11450
rect 37060 11396 37066 11398
rect 37122 11396 37146 11398
rect 37202 11396 37226 11398
rect 37282 11396 37306 11398
rect 37362 11396 37368 11398
rect 37060 11387 37368 11396
rect 37660 11370 37688 12174
rect 37832 11688 37884 11694
rect 37832 11630 37884 11636
rect 37660 11342 37780 11370
rect 37844 11354 37872 11630
rect 37648 11280 37700 11286
rect 37648 11222 37700 11228
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 37568 10742 37596 11086
rect 37556 10736 37608 10742
rect 37556 10678 37608 10684
rect 37060 10364 37368 10373
rect 37060 10362 37066 10364
rect 37122 10362 37146 10364
rect 37202 10362 37226 10364
rect 37282 10362 37306 10364
rect 37362 10362 37368 10364
rect 37122 10310 37124 10362
rect 37304 10310 37306 10362
rect 37060 10308 37066 10310
rect 37122 10308 37146 10310
rect 37202 10308 37226 10310
rect 37282 10308 37306 10310
rect 37362 10308 37368 10310
rect 37060 10299 37368 10308
rect 36924 10118 37320 10146
rect 36924 10062 36952 10118
rect 36912 10056 36964 10062
rect 36634 10024 36690 10033
rect 37188 10056 37240 10062
rect 36912 9998 36964 10004
rect 37094 10024 37150 10033
rect 36634 9959 36690 9968
rect 37150 10004 37188 10010
rect 37150 9998 37240 10004
rect 37150 9982 37228 9998
rect 37094 9959 37150 9968
rect 37292 9450 37320 10118
rect 37372 10124 37424 10130
rect 37372 10066 37424 10072
rect 37280 9444 37332 9450
rect 37280 9386 37332 9392
rect 37384 9382 37412 10066
rect 37660 9586 37688 11222
rect 37752 11218 37780 11342
rect 37832 11348 37884 11354
rect 37832 11290 37884 11296
rect 37936 11234 37964 12406
rect 38304 12102 38332 14214
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 38108 11756 38160 11762
rect 38108 11698 38160 11704
rect 37740 11212 37792 11218
rect 37740 11154 37792 11160
rect 37844 11206 37964 11234
rect 37844 10130 37872 11206
rect 38120 11121 38148 11698
rect 38106 11112 38162 11121
rect 38396 11082 38424 17478
rect 38488 16436 38516 19314
rect 38672 18970 38700 19858
rect 38660 18964 38712 18970
rect 38660 18906 38712 18912
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38764 17678 38792 18022
rect 38752 17672 38804 17678
rect 38752 17614 38804 17620
rect 38568 17536 38620 17542
rect 38568 17478 38620 17484
rect 38580 16590 38608 17478
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38568 16584 38620 16590
rect 38568 16526 38620 16532
rect 38488 16408 38608 16436
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38488 12646 38516 14350
rect 38476 12640 38528 12646
rect 38476 12582 38528 12588
rect 38106 11047 38162 11056
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 38016 11008 38068 11014
rect 38016 10950 38068 10956
rect 37936 10198 37964 10950
rect 37924 10192 37976 10198
rect 37924 10134 37976 10140
rect 37832 10124 37884 10130
rect 37832 10066 37884 10072
rect 37648 9580 37700 9586
rect 37648 9522 37700 9528
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 37372 9376 37424 9382
rect 37372 9318 37424 9324
rect 37648 9376 37700 9382
rect 37648 9318 37700 9324
rect 36544 9172 36596 9178
rect 36544 9114 36596 9120
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 36372 8090 36400 8910
rect 36544 8832 36596 8838
rect 36544 8774 36596 8780
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36372 7546 36400 7754
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 36360 7540 36412 7546
rect 36360 7482 36412 7488
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 36188 6866 36216 7278
rect 36372 6866 36400 7482
rect 36464 6866 36492 8434
rect 36556 7818 36584 8774
rect 36544 7812 36596 7818
rect 36544 7754 36596 7760
rect 36740 6934 36768 9318
rect 37060 9276 37368 9285
rect 37060 9274 37066 9276
rect 37122 9274 37146 9276
rect 37202 9274 37226 9276
rect 37282 9274 37306 9276
rect 37362 9274 37368 9276
rect 37122 9222 37124 9274
rect 37304 9222 37306 9274
rect 37060 9220 37066 9222
rect 37122 9220 37146 9222
rect 37202 9220 37226 9222
rect 37282 9220 37306 9222
rect 37362 9220 37368 9222
rect 37060 9211 37368 9220
rect 36912 9036 36964 9042
rect 36912 8978 36964 8984
rect 36820 8968 36872 8974
rect 36820 8910 36872 8916
rect 36832 7274 36860 8910
rect 36924 8362 36952 8978
rect 37556 8900 37608 8906
rect 37556 8842 37608 8848
rect 37004 8492 37056 8498
rect 37004 8434 37056 8440
rect 37016 8362 37044 8434
rect 37568 8430 37596 8842
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 37556 8424 37608 8430
rect 37556 8366 37608 8372
rect 36912 8356 36964 8362
rect 36912 8298 36964 8304
rect 37004 8356 37056 8362
rect 37004 8298 37056 8304
rect 36820 7268 36872 7274
rect 36820 7210 36872 7216
rect 36728 6928 36780 6934
rect 36728 6870 36780 6876
rect 36924 6882 36952 8298
rect 37108 8294 37136 8366
rect 37096 8288 37148 8294
rect 37096 8230 37148 8236
rect 37060 8188 37368 8197
rect 37060 8186 37066 8188
rect 37122 8186 37146 8188
rect 37202 8186 37226 8188
rect 37282 8186 37306 8188
rect 37362 8186 37368 8188
rect 37122 8134 37124 8186
rect 37304 8134 37306 8186
rect 37060 8132 37066 8134
rect 37122 8132 37146 8134
rect 37202 8132 37226 8134
rect 37282 8132 37306 8134
rect 37362 8132 37368 8134
rect 37060 8123 37368 8132
rect 37060 7100 37368 7109
rect 37060 7098 37066 7100
rect 37122 7098 37146 7100
rect 37202 7098 37226 7100
rect 37282 7098 37306 7100
rect 37362 7098 37368 7100
rect 37122 7046 37124 7098
rect 37304 7046 37306 7098
rect 37060 7044 37066 7046
rect 37122 7044 37146 7046
rect 37202 7044 37226 7046
rect 37282 7044 37306 7046
rect 37362 7044 37368 7046
rect 37060 7035 37368 7044
rect 36924 6866 37044 6882
rect 37660 6866 37688 9318
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37844 7818 37872 8774
rect 37936 8430 37964 10134
rect 38028 10130 38056 10950
rect 38016 10124 38068 10130
rect 38016 10066 38068 10072
rect 38292 10124 38344 10130
rect 38292 10066 38344 10072
rect 38028 9722 38056 10066
rect 38304 9926 38332 10066
rect 38292 9920 38344 9926
rect 38292 9862 38344 9868
rect 38016 9716 38068 9722
rect 38016 9658 38068 9664
rect 38304 9654 38332 9862
rect 38292 9648 38344 9654
rect 38292 9590 38344 9596
rect 38304 9178 38332 9590
rect 38292 9172 38344 9178
rect 38292 9114 38344 9120
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 37832 7812 37884 7818
rect 37832 7754 37884 7760
rect 37936 7546 37964 8366
rect 37924 7540 37976 7546
rect 37924 7482 37976 7488
rect 37936 7426 37964 7482
rect 37844 7398 37964 7426
rect 36176 6860 36228 6866
rect 36176 6802 36228 6808
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 36452 6860 36504 6866
rect 36924 6860 37056 6866
rect 36924 6854 37004 6860
rect 36452 6802 36504 6808
rect 37004 6802 37056 6808
rect 37648 6860 37700 6866
rect 37648 6802 37700 6808
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 35900 5296 35952 5302
rect 35900 5238 35952 5244
rect 35912 4622 35940 5238
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35912 4282 35940 4558
rect 35900 4276 35952 4282
rect 35820 4236 35900 4264
rect 35820 3534 35848 4236
rect 35900 4218 35952 4224
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35900 3392 35952 3398
rect 35900 3334 35952 3340
rect 35716 3188 35768 3194
rect 35716 3130 35768 3136
rect 35624 2576 35676 2582
rect 35624 2518 35676 2524
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35820 1170 35848 2450
rect 35912 2446 35940 3334
rect 36004 2774 36032 6666
rect 36188 6458 36216 6802
rect 37188 6792 37240 6798
rect 37188 6734 37240 6740
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 37200 6322 37228 6734
rect 36728 6316 36780 6322
rect 36728 6258 36780 6264
rect 37188 6316 37240 6322
rect 37188 6258 37240 6264
rect 36740 5302 36768 6258
rect 37464 6112 37516 6118
rect 37464 6054 37516 6060
rect 37060 6012 37368 6021
rect 37060 6010 37066 6012
rect 37122 6010 37146 6012
rect 37202 6010 37226 6012
rect 37282 6010 37306 6012
rect 37362 6010 37368 6012
rect 37122 5958 37124 6010
rect 37304 5958 37306 6010
rect 37060 5956 37066 5958
rect 37122 5956 37146 5958
rect 37202 5956 37226 5958
rect 37282 5956 37306 5958
rect 37362 5956 37368 5958
rect 37060 5947 37368 5956
rect 37476 5914 37504 6054
rect 37464 5908 37516 5914
rect 37464 5850 37516 5856
rect 37660 5846 37688 6802
rect 37844 6458 37872 7398
rect 37924 7336 37976 7342
rect 37924 7278 37976 7284
rect 37936 7002 37964 7278
rect 37924 6996 37976 7002
rect 37924 6938 37976 6944
rect 37832 6452 37884 6458
rect 37832 6394 37884 6400
rect 38108 6316 38160 6322
rect 38108 6258 38160 6264
rect 38120 5914 38148 6258
rect 38292 6112 38344 6118
rect 38292 6054 38344 6060
rect 38108 5908 38160 5914
rect 38108 5850 38160 5856
rect 37648 5840 37700 5846
rect 37648 5782 37700 5788
rect 36820 5636 36872 5642
rect 36820 5578 36872 5584
rect 36832 5370 36860 5578
rect 38200 5568 38252 5574
rect 38200 5510 38252 5516
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 37556 5364 37608 5370
rect 37556 5306 37608 5312
rect 36728 5296 36780 5302
rect 36728 5238 36780 5244
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 36176 5092 36228 5098
rect 36176 5034 36228 5040
rect 36188 3398 36216 5034
rect 37060 4924 37368 4933
rect 37060 4922 37066 4924
rect 37122 4922 37146 4924
rect 37202 4922 37226 4924
rect 37282 4922 37306 4924
rect 37362 4922 37368 4924
rect 37122 4870 37124 4922
rect 37304 4870 37306 4922
rect 37060 4868 37066 4870
rect 37122 4868 37146 4870
rect 37202 4868 37226 4870
rect 37282 4868 37306 4870
rect 37362 4868 37368 4870
rect 37060 4859 37368 4868
rect 36268 4548 36320 4554
rect 36268 4490 36320 4496
rect 36452 4548 36504 4554
rect 36452 4490 36504 4496
rect 36280 4078 36308 4490
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36004 2746 36124 2774
rect 36096 2650 36124 2746
rect 36084 2644 36136 2650
rect 36084 2586 36136 2592
rect 36188 2446 36216 2858
rect 36372 2774 36400 4082
rect 36464 3942 36492 4490
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36556 3058 36584 4082
rect 36912 4072 36964 4078
rect 36912 4014 36964 4020
rect 36820 3936 36872 3942
rect 36820 3878 36872 3884
rect 36832 3466 36860 3878
rect 36820 3460 36872 3466
rect 36820 3402 36872 3408
rect 36544 3052 36596 3058
rect 36544 2994 36596 3000
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 36280 2746 36400 2774
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 35728 1142 35848 1170
rect 35728 800 35756 1142
rect 36280 800 36308 2746
rect 36832 2650 36860 2994
rect 36820 2644 36872 2650
rect 36820 2586 36872 2592
rect 36924 2446 36952 4014
rect 37060 3836 37368 3845
rect 37060 3834 37066 3836
rect 37122 3834 37146 3836
rect 37202 3834 37226 3836
rect 37282 3834 37306 3836
rect 37362 3834 37368 3836
rect 37122 3782 37124 3834
rect 37304 3782 37306 3834
rect 37060 3780 37066 3782
rect 37122 3780 37146 3782
rect 37202 3780 37226 3782
rect 37282 3780 37306 3782
rect 37362 3780 37368 3782
rect 37060 3771 37368 3780
rect 37476 3534 37504 5170
rect 37568 4826 37596 5306
rect 38212 5234 38240 5510
rect 38200 5228 38252 5234
rect 38200 5170 38252 5176
rect 37556 4820 37608 4826
rect 37556 4762 37608 4768
rect 37568 4049 37596 4762
rect 38304 4622 38332 6054
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 37648 4480 37700 4486
rect 37648 4422 37700 4428
rect 37660 4214 37688 4422
rect 38396 4214 38424 11018
rect 38488 9178 38516 12582
rect 38580 11898 38608 16408
rect 38672 14770 38700 16934
rect 38936 16788 38988 16794
rect 38936 16730 38988 16736
rect 38752 16584 38804 16590
rect 38752 16526 38804 16532
rect 38764 16454 38792 16526
rect 38752 16448 38804 16454
rect 38752 16390 38804 16396
rect 38764 16250 38792 16390
rect 38752 16244 38804 16250
rect 38752 16186 38804 16192
rect 38672 14742 38884 14770
rect 38752 14476 38804 14482
rect 38752 14418 38804 14424
rect 38660 14272 38712 14278
rect 38660 14214 38712 14220
rect 38672 13870 38700 14214
rect 38660 13864 38712 13870
rect 38660 13806 38712 13812
rect 38568 11892 38620 11898
rect 38568 11834 38620 11840
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38580 9722 38608 10610
rect 38568 9716 38620 9722
rect 38568 9658 38620 9664
rect 38476 9172 38528 9178
rect 38476 9114 38528 9120
rect 38764 7750 38792 14418
rect 38856 12434 38884 14742
rect 38948 14074 38976 16730
rect 39040 16726 39068 19858
rect 39132 19514 39160 19994
rect 39120 19508 39172 19514
rect 39120 19450 39172 19456
rect 39592 19446 39620 20742
rect 40052 19922 40080 22918
rect 40604 22642 40632 24006
rect 41156 23866 41184 24142
rect 41696 24064 41748 24070
rect 41696 24006 41748 24012
rect 41144 23860 41196 23866
rect 41144 23802 41196 23808
rect 41604 23656 41656 23662
rect 41604 23598 41656 23604
rect 41236 23520 41288 23526
rect 41236 23462 41288 23468
rect 41512 23520 41564 23526
rect 41512 23462 41564 23468
rect 40960 22976 41012 22982
rect 40960 22918 41012 22924
rect 40592 22636 40644 22642
rect 40592 22578 40644 22584
rect 40972 22094 41000 22918
rect 40696 22066 41000 22094
rect 41248 22094 41276 23462
rect 41524 23322 41552 23462
rect 41512 23316 41564 23322
rect 41512 23258 41564 23264
rect 41328 23044 41380 23050
rect 41512 23044 41564 23050
rect 41380 23004 41460 23032
rect 41328 22986 41380 22992
rect 41432 22710 41460 23004
rect 41512 22986 41564 22992
rect 41420 22704 41472 22710
rect 41420 22646 41472 22652
rect 41524 22166 41552 22986
rect 41616 22778 41644 23598
rect 41604 22772 41656 22778
rect 41604 22714 41656 22720
rect 41708 22642 41736 24006
rect 42260 22982 42288 24550
rect 42340 24200 42392 24206
rect 42340 24142 42392 24148
rect 42524 24200 42576 24206
rect 42524 24142 42576 24148
rect 42248 22976 42300 22982
rect 42248 22918 42300 22924
rect 42352 22778 42380 24142
rect 42536 23526 42564 24142
rect 42524 23520 42576 23526
rect 42524 23462 42576 23468
rect 42340 22772 42392 22778
rect 42340 22714 42392 22720
rect 42536 22710 42564 23462
rect 42628 23186 42656 24806
rect 42708 24754 42760 24760
rect 42892 24812 42944 24818
rect 42892 24754 42944 24760
rect 42708 24676 42760 24682
rect 42708 24618 42760 24624
rect 42720 24410 42748 24618
rect 42800 24608 42852 24614
rect 42800 24550 42852 24556
rect 42812 24410 42840 24550
rect 42708 24404 42760 24410
rect 42708 24346 42760 24352
rect 42800 24404 42852 24410
rect 42800 24346 42852 24352
rect 42720 23798 42748 24346
rect 42904 23798 42932 24754
rect 42984 24608 43036 24614
rect 42984 24550 43036 24556
rect 42996 24206 43024 24550
rect 42984 24200 43036 24206
rect 42984 24142 43036 24148
rect 43996 24200 44048 24206
rect 43996 24142 44048 24148
rect 42708 23792 42760 23798
rect 42708 23734 42760 23740
rect 42892 23792 42944 23798
rect 42892 23734 42944 23740
rect 42616 23180 42668 23186
rect 42616 23122 42668 23128
rect 42524 22704 42576 22710
rect 42524 22646 42576 22652
rect 41696 22636 41748 22642
rect 41696 22578 41748 22584
rect 42720 22556 42748 23734
rect 42904 22778 42932 23734
rect 43444 23180 43496 23186
rect 43444 23122 43496 23128
rect 43456 22982 43484 23122
rect 43628 23112 43680 23118
rect 43628 23054 43680 23060
rect 43720 23112 43772 23118
rect 43720 23054 43772 23060
rect 43076 22976 43128 22982
rect 43076 22918 43128 22924
rect 43444 22976 43496 22982
rect 43444 22918 43496 22924
rect 42892 22772 42944 22778
rect 42892 22714 42944 22720
rect 42536 22528 42748 22556
rect 42248 22432 42300 22438
rect 42248 22374 42300 22380
rect 41512 22160 41564 22166
rect 41512 22102 41564 22108
rect 41328 22094 41380 22098
rect 41248 22092 41380 22094
rect 41248 22066 41328 22092
rect 40500 20936 40552 20942
rect 40500 20878 40552 20884
rect 40224 20800 40276 20806
rect 40224 20742 40276 20748
rect 40408 20800 40460 20806
rect 40408 20742 40460 20748
rect 40236 20534 40264 20742
rect 40224 20528 40276 20534
rect 40224 20470 40276 20476
rect 40420 19922 40448 20742
rect 40040 19916 40092 19922
rect 40040 19858 40092 19864
rect 40408 19916 40460 19922
rect 40408 19858 40460 19864
rect 39856 19712 39908 19718
rect 39856 19654 39908 19660
rect 39580 19440 39632 19446
rect 39580 19382 39632 19388
rect 39868 18290 39896 19654
rect 40420 18630 40448 19858
rect 40512 19446 40540 20878
rect 40500 19440 40552 19446
rect 40500 19382 40552 19388
rect 40408 18624 40460 18630
rect 40408 18566 40460 18572
rect 39856 18284 39908 18290
rect 39856 18226 39908 18232
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40052 17814 40080 18022
rect 40040 17808 40092 17814
rect 40040 17750 40092 17756
rect 39672 17536 39724 17542
rect 39672 17478 39724 17484
rect 39856 17536 39908 17542
rect 39856 17478 39908 17484
rect 39684 17134 39712 17478
rect 39868 17338 39896 17478
rect 39856 17332 39908 17338
rect 39856 17274 39908 17280
rect 39212 17128 39264 17134
rect 39488 17128 39540 17134
rect 39212 17070 39264 17076
rect 39408 17076 39488 17082
rect 39408 17070 39540 17076
rect 39672 17128 39724 17134
rect 39672 17070 39724 17076
rect 39120 16992 39172 16998
rect 39120 16934 39172 16940
rect 39028 16720 39080 16726
rect 39028 16662 39080 16668
rect 39040 14618 39068 16662
rect 39028 14612 39080 14618
rect 39028 14554 39080 14560
rect 39132 14482 39160 16934
rect 39224 16794 39252 17070
rect 39408 17054 39528 17070
rect 39408 16998 39436 17054
rect 39396 16992 39448 16998
rect 39396 16934 39448 16940
rect 39488 16992 39540 16998
rect 39488 16934 39540 16940
rect 39212 16788 39264 16794
rect 39212 16730 39264 16736
rect 39224 16114 39252 16730
rect 39500 16658 39528 16934
rect 39488 16652 39540 16658
rect 39488 16594 39540 16600
rect 39212 16108 39264 16114
rect 39212 16050 39264 16056
rect 39396 14612 39448 14618
rect 39396 14554 39448 14560
rect 39120 14476 39172 14482
rect 39120 14418 39172 14424
rect 38936 14068 38988 14074
rect 38936 14010 38988 14016
rect 39408 13870 39436 14554
rect 39396 13864 39448 13870
rect 39224 13812 39396 13818
rect 39224 13806 39448 13812
rect 39224 13790 39436 13806
rect 38856 12406 39068 12434
rect 39040 11150 39068 12406
rect 39028 11144 39080 11150
rect 39028 11086 39080 11092
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38856 10266 38884 10406
rect 38844 10260 38896 10266
rect 38844 10202 38896 10208
rect 38936 9920 38988 9926
rect 38936 9862 38988 9868
rect 38948 9586 38976 9862
rect 38936 9580 38988 9586
rect 38936 9522 38988 9528
rect 38936 8424 38988 8430
rect 38936 8366 38988 8372
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38844 7268 38896 7274
rect 38844 7210 38896 7216
rect 38614 6860 38666 6866
rect 38488 6820 38614 6848
rect 38488 6458 38516 6820
rect 38614 6802 38666 6808
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 38856 6322 38884 7210
rect 38948 6866 38976 8366
rect 39132 8090 39160 8366
rect 39120 8084 39172 8090
rect 39120 8026 39172 8032
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39132 7546 39160 7822
rect 39120 7540 39172 7546
rect 39120 7482 39172 7488
rect 39224 7206 39252 13790
rect 39396 13252 39448 13258
rect 39396 13194 39448 13200
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39316 12306 39344 13126
rect 39304 12300 39356 12306
rect 39304 12242 39356 12248
rect 39408 12238 39436 13194
rect 39396 12232 39448 12238
rect 39396 12174 39448 12180
rect 39304 11008 39356 11014
rect 39304 10950 39356 10956
rect 39316 10810 39344 10950
rect 39304 10804 39356 10810
rect 39304 10746 39356 10752
rect 39684 8974 39712 17070
rect 39868 16726 39896 17274
rect 39856 16720 39908 16726
rect 39856 16662 39908 16668
rect 40052 14550 40080 17750
rect 40408 17672 40460 17678
rect 40408 17614 40460 17620
rect 40132 17604 40184 17610
rect 40132 17546 40184 17552
rect 40144 17338 40172 17546
rect 40132 17332 40184 17338
rect 40132 17274 40184 17280
rect 40420 16590 40448 17614
rect 40696 17542 40724 22066
rect 41328 22034 41380 22040
rect 42260 21554 42288 22374
rect 42248 21548 42300 21554
rect 42248 21490 42300 21496
rect 42536 21486 42564 22528
rect 42616 22432 42668 22438
rect 42616 22374 42668 22380
rect 42628 22166 42656 22374
rect 42616 22160 42668 22166
rect 42616 22102 42668 22108
rect 42524 21480 42576 21486
rect 42524 21422 42576 21428
rect 42156 21344 42208 21350
rect 42156 21286 42208 21292
rect 40868 20460 40920 20466
rect 40868 20402 40920 20408
rect 40880 19378 40908 20402
rect 41052 20256 41104 20262
rect 41052 20198 41104 20204
rect 41420 20256 41472 20262
rect 41420 20198 41472 20204
rect 41696 20256 41748 20262
rect 41696 20198 41748 20204
rect 41064 19854 41092 20198
rect 41052 19848 41104 19854
rect 41052 19790 41104 19796
rect 41236 19848 41288 19854
rect 41236 19790 41288 19796
rect 41064 19446 41092 19790
rect 41248 19514 41276 19790
rect 41236 19508 41288 19514
rect 41236 19450 41288 19456
rect 41052 19440 41104 19446
rect 41052 19382 41104 19388
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 40776 19304 40828 19310
rect 40776 19246 40828 19252
rect 40788 18970 40816 19246
rect 41432 19174 41460 20198
rect 41708 19854 41736 20198
rect 41696 19848 41748 19854
rect 41696 19790 41748 19796
rect 41420 19168 41472 19174
rect 41420 19110 41472 19116
rect 41788 19168 41840 19174
rect 41788 19110 41840 19116
rect 40776 18964 40828 18970
rect 40828 18924 41000 18952
rect 40776 18906 40828 18912
rect 40592 17536 40644 17542
rect 40592 17478 40644 17484
rect 40684 17536 40736 17542
rect 40684 17478 40736 17484
rect 40408 16584 40460 16590
rect 40408 16526 40460 16532
rect 40604 16182 40632 17478
rect 40696 17270 40724 17478
rect 40684 17264 40736 17270
rect 40684 17206 40736 17212
rect 40592 16176 40644 16182
rect 40592 16118 40644 16124
rect 40040 14544 40092 14550
rect 40040 14486 40092 14492
rect 40052 14006 40080 14486
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 40236 14074 40264 14350
rect 40776 14340 40828 14346
rect 40776 14282 40828 14288
rect 40224 14068 40276 14074
rect 40224 14010 40276 14016
rect 40040 14000 40092 14006
rect 40040 13942 40092 13948
rect 39764 13864 39816 13870
rect 39764 13806 39816 13812
rect 40500 13864 40552 13870
rect 40500 13806 40552 13812
rect 39776 13326 39804 13806
rect 39948 13728 40000 13734
rect 39948 13670 40000 13676
rect 40040 13728 40092 13734
rect 40040 13670 40092 13676
rect 39960 13569 39988 13670
rect 39946 13560 40002 13569
rect 39946 13495 40002 13504
rect 39764 13320 39816 13326
rect 39764 13262 39816 13268
rect 39856 13320 39908 13326
rect 39856 13262 39908 13268
rect 39776 12434 39804 13262
rect 39868 12986 39896 13262
rect 39856 12980 39908 12986
rect 39856 12922 39908 12928
rect 40052 12918 40080 13670
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 40316 12640 40368 12646
rect 40316 12582 40368 12588
rect 40408 12640 40460 12646
rect 40408 12582 40460 12588
rect 39776 12406 39896 12434
rect 39868 11218 39896 12406
rect 40040 11552 40092 11558
rect 40040 11494 40092 11500
rect 39856 11212 39908 11218
rect 39856 11154 39908 11160
rect 40052 10742 40080 11494
rect 40224 11076 40276 11082
rect 40224 11018 40276 11024
rect 40040 10736 40092 10742
rect 40040 10678 40092 10684
rect 40236 9654 40264 11018
rect 40328 10418 40356 12582
rect 40420 12306 40448 12582
rect 40512 12434 40540 13806
rect 40788 12918 40816 14282
rect 40868 14272 40920 14278
rect 40868 14214 40920 14220
rect 40880 14074 40908 14214
rect 40868 14068 40920 14074
rect 40868 14010 40920 14016
rect 40776 12912 40828 12918
rect 40776 12854 40828 12860
rect 40788 12442 40816 12854
rect 40972 12782 41000 18924
rect 41144 17672 41196 17678
rect 41144 17614 41196 17620
rect 41328 17672 41380 17678
rect 41328 17614 41380 17620
rect 41156 17338 41184 17614
rect 41144 17332 41196 17338
rect 41144 17274 41196 17280
rect 41340 16590 41368 17614
rect 41512 17128 41564 17134
rect 41512 17070 41564 17076
rect 41328 16584 41380 16590
rect 41328 16526 41380 16532
rect 41524 16250 41552 17070
rect 41604 16516 41656 16522
rect 41604 16458 41656 16464
rect 41616 16250 41644 16458
rect 41512 16244 41564 16250
rect 41512 16186 41564 16192
rect 41604 16244 41656 16250
rect 41604 16186 41656 16192
rect 41800 14822 41828 19110
rect 42168 15570 42196 21286
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 42352 16182 42380 20878
rect 42432 19304 42484 19310
rect 42432 19246 42484 19252
rect 42444 18766 42472 19246
rect 42432 18760 42484 18766
rect 42432 18702 42484 18708
rect 42444 17678 42472 18702
rect 42432 17672 42484 17678
rect 42432 17614 42484 17620
rect 42444 16794 42472 17614
rect 42536 17338 42564 21422
rect 42628 21350 42656 22102
rect 42904 21894 42932 22714
rect 43088 22098 43116 22918
rect 43168 22568 43220 22574
rect 43168 22510 43220 22516
rect 43076 22092 43128 22098
rect 43076 22034 43128 22040
rect 43180 21894 43208 22510
rect 43640 22166 43668 23054
rect 43732 22710 43760 23054
rect 44008 22778 44036 24142
rect 43996 22772 44048 22778
rect 43996 22714 44048 22720
rect 44192 22710 44220 26250
rect 44282 26140 44590 26149
rect 44282 26138 44288 26140
rect 44344 26138 44368 26140
rect 44424 26138 44448 26140
rect 44504 26138 44528 26140
rect 44584 26138 44590 26140
rect 44344 26086 44346 26138
rect 44526 26086 44528 26138
rect 44282 26084 44288 26086
rect 44344 26084 44368 26086
rect 44424 26084 44448 26086
rect 44504 26084 44528 26086
rect 44584 26084 44590 26086
rect 44282 26075 44590 26084
rect 45204 26042 45232 26862
rect 45468 26852 45520 26858
rect 45468 26794 45520 26800
rect 45376 26308 45428 26314
rect 45376 26250 45428 26256
rect 45192 26036 45244 26042
rect 45192 25978 45244 25984
rect 44916 25356 44968 25362
rect 44916 25298 44968 25304
rect 44282 25052 44590 25061
rect 44282 25050 44288 25052
rect 44344 25050 44368 25052
rect 44424 25050 44448 25052
rect 44504 25050 44528 25052
rect 44584 25050 44590 25052
rect 44344 24998 44346 25050
rect 44526 24998 44528 25050
rect 44282 24996 44288 24998
rect 44344 24996 44368 24998
rect 44424 24996 44448 24998
rect 44504 24996 44528 24998
rect 44584 24996 44590 24998
rect 44282 24987 44590 24996
rect 44640 24744 44692 24750
rect 44640 24686 44692 24692
rect 44652 24410 44680 24686
rect 44640 24404 44692 24410
rect 44640 24346 44692 24352
rect 44640 24064 44692 24070
rect 44640 24006 44692 24012
rect 44282 23964 44590 23973
rect 44282 23962 44288 23964
rect 44344 23962 44368 23964
rect 44424 23962 44448 23964
rect 44504 23962 44528 23964
rect 44584 23962 44590 23964
rect 44344 23910 44346 23962
rect 44526 23910 44528 23962
rect 44282 23908 44288 23910
rect 44344 23908 44368 23910
rect 44424 23908 44448 23910
rect 44504 23908 44528 23910
rect 44584 23908 44590 23910
rect 44282 23899 44590 23908
rect 44652 23730 44680 24006
rect 44272 23724 44324 23730
rect 44272 23666 44324 23672
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44284 23322 44312 23666
rect 44640 23520 44692 23526
rect 44640 23462 44692 23468
rect 44272 23316 44324 23322
rect 44272 23258 44324 23264
rect 44282 22876 44590 22885
rect 44282 22874 44288 22876
rect 44344 22874 44368 22876
rect 44424 22874 44448 22876
rect 44504 22874 44528 22876
rect 44584 22874 44590 22876
rect 44344 22822 44346 22874
rect 44526 22822 44528 22874
rect 44282 22820 44288 22822
rect 44344 22820 44368 22822
rect 44424 22820 44448 22822
rect 44504 22820 44528 22822
rect 44584 22820 44590 22822
rect 44282 22811 44590 22820
rect 43720 22704 43772 22710
rect 43720 22646 43772 22652
rect 44180 22704 44232 22710
rect 44180 22646 44232 22652
rect 43628 22160 43680 22166
rect 43628 22102 43680 22108
rect 42892 21888 42944 21894
rect 42892 21830 42944 21836
rect 43168 21888 43220 21894
rect 43168 21830 43220 21836
rect 42616 21344 42668 21350
rect 42616 21286 42668 21292
rect 42904 20806 42932 21830
rect 43180 20942 43208 21830
rect 43732 21690 43760 22646
rect 44652 22642 44680 23462
rect 44732 22976 44784 22982
rect 44732 22918 44784 22924
rect 44640 22636 44692 22642
rect 44640 22578 44692 22584
rect 44640 21888 44692 21894
rect 44640 21830 44692 21836
rect 44282 21788 44590 21797
rect 44282 21786 44288 21788
rect 44344 21786 44368 21788
rect 44424 21786 44448 21788
rect 44504 21786 44528 21788
rect 44584 21786 44590 21788
rect 44344 21734 44346 21786
rect 44526 21734 44528 21786
rect 44282 21732 44288 21734
rect 44344 21732 44368 21734
rect 44424 21732 44448 21734
rect 44504 21732 44528 21734
rect 44584 21732 44590 21734
rect 44282 21723 44590 21732
rect 43720 21684 43772 21690
rect 43720 21626 43772 21632
rect 43168 20936 43220 20942
rect 43168 20878 43220 20884
rect 44180 20936 44232 20942
rect 44180 20878 44232 20884
rect 43904 20868 43956 20874
rect 43904 20810 43956 20816
rect 42892 20800 42944 20806
rect 42892 20742 42944 20748
rect 43076 20800 43128 20806
rect 43076 20742 43128 20748
rect 42904 20602 42932 20742
rect 42892 20596 42944 20602
rect 42892 20538 42944 20544
rect 42984 20528 43036 20534
rect 42984 20470 43036 20476
rect 42996 19990 43024 20470
rect 42984 19984 43036 19990
rect 42984 19926 43036 19932
rect 43088 19378 43116 20742
rect 43720 20596 43772 20602
rect 43720 20538 43772 20544
rect 43260 20392 43312 20398
rect 43260 20334 43312 20340
rect 43272 20058 43300 20334
rect 43628 20324 43680 20330
rect 43628 20266 43680 20272
rect 43260 20052 43312 20058
rect 43260 19994 43312 20000
rect 43640 19922 43668 20266
rect 43628 19916 43680 19922
rect 43628 19858 43680 19864
rect 43732 19378 43760 20538
rect 43812 20460 43864 20466
rect 43812 20402 43864 20408
rect 43824 19922 43852 20402
rect 43916 19922 43944 20810
rect 43996 20324 44048 20330
rect 43996 20266 44048 20272
rect 43812 19916 43864 19922
rect 43812 19858 43864 19864
rect 43904 19916 43956 19922
rect 43904 19858 43956 19864
rect 43076 19372 43128 19378
rect 43076 19314 43128 19320
rect 43720 19372 43772 19378
rect 43720 19314 43772 19320
rect 43904 19304 43956 19310
rect 43904 19246 43956 19252
rect 43916 18086 43944 19246
rect 43168 18080 43220 18086
rect 43168 18022 43220 18028
rect 43904 18080 43956 18086
rect 43904 18022 43956 18028
rect 42524 17332 42576 17338
rect 42524 17274 42576 17280
rect 42432 16788 42484 16794
rect 42432 16730 42484 16736
rect 42340 16176 42392 16182
rect 42340 16118 42392 16124
rect 42352 15638 42380 16118
rect 42340 15632 42392 15638
rect 42340 15574 42392 15580
rect 42156 15564 42208 15570
rect 42156 15506 42208 15512
rect 41788 14816 41840 14822
rect 41788 14758 41840 14764
rect 42432 14816 42484 14822
rect 42432 14758 42484 14764
rect 42444 14482 42472 14758
rect 42432 14476 42484 14482
rect 42432 14418 42484 14424
rect 41144 14272 41196 14278
rect 41144 14214 41196 14220
rect 41156 14006 41184 14214
rect 41144 14000 41196 14006
rect 41144 13942 41196 13948
rect 41604 13728 41656 13734
rect 41604 13670 41656 13676
rect 41616 13394 41644 13670
rect 41604 13388 41656 13394
rect 41604 13330 41656 13336
rect 41616 12986 41644 13330
rect 42340 13252 42392 13258
rect 42340 13194 42392 13200
rect 41604 12980 41656 12986
rect 41604 12922 41656 12928
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 40776 12436 40828 12442
rect 40512 12406 40632 12434
rect 40408 12300 40460 12306
rect 40408 12242 40460 12248
rect 40328 10390 40448 10418
rect 40224 9648 40276 9654
rect 40224 9590 40276 9596
rect 40132 9376 40184 9382
rect 40132 9318 40184 9324
rect 39672 8968 39724 8974
rect 39672 8910 39724 8916
rect 39488 8900 39540 8906
rect 39488 8842 39540 8848
rect 39304 8288 39356 8294
rect 39304 8230 39356 8236
rect 39316 7886 39344 8230
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39396 7744 39448 7750
rect 39396 7686 39448 7692
rect 39212 7200 39264 7206
rect 39212 7142 39264 7148
rect 39304 7200 39356 7206
rect 39304 7142 39356 7148
rect 38936 6860 38988 6866
rect 38936 6802 38988 6808
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38844 6316 38896 6322
rect 38844 6258 38896 6264
rect 38660 5704 38712 5710
rect 38660 5646 38712 5652
rect 38672 4826 38700 5646
rect 38752 5024 38804 5030
rect 38752 4966 38804 4972
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 38660 4820 38712 4826
rect 38660 4762 38712 4768
rect 38764 4690 38792 4966
rect 38856 4690 38884 4966
rect 38752 4684 38804 4690
rect 38752 4626 38804 4632
rect 38844 4684 38896 4690
rect 38844 4626 38896 4632
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 38384 4208 38436 4214
rect 38384 4150 38436 4156
rect 38108 4140 38160 4146
rect 38108 4082 38160 4088
rect 38200 4140 38252 4146
rect 38200 4082 38252 4088
rect 38660 4140 38712 4146
rect 38856 4128 38884 4626
rect 38712 4100 38884 4128
rect 38660 4082 38712 4088
rect 37554 4040 37610 4049
rect 37554 3975 37610 3984
rect 37464 3528 37516 3534
rect 37002 3496 37058 3505
rect 37464 3470 37516 3476
rect 37002 3431 37058 3440
rect 37016 3194 37044 3431
rect 38120 3398 38148 4082
rect 38212 3738 38240 4082
rect 38200 3732 38252 3738
rect 38200 3674 38252 3680
rect 38568 3732 38620 3738
rect 38568 3674 38620 3680
rect 38108 3392 38160 3398
rect 38108 3334 38160 3340
rect 38212 3194 38240 3674
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37922 2952 37978 2961
rect 37060 2748 37368 2757
rect 37060 2746 37066 2748
rect 37122 2746 37146 2748
rect 37202 2746 37226 2748
rect 37282 2746 37306 2748
rect 37362 2746 37368 2748
rect 37122 2694 37124 2746
rect 37304 2694 37306 2746
rect 37060 2692 37066 2694
rect 37122 2692 37146 2694
rect 37202 2692 37226 2694
rect 37282 2692 37306 2694
rect 37362 2692 37368 2694
rect 37060 2683 37368 2692
rect 36820 2440 36872 2446
rect 36820 2382 36872 2388
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 36832 800 36860 2382
rect 37384 870 37504 898
rect 37384 800 37412 870
rect 34164 734 34468 762
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37476 762 37504 870
rect 37660 762 37688 2926
rect 37922 2887 37978 2896
rect 37936 800 37964 2887
rect 38580 2650 38608 3674
rect 38672 2854 38700 4082
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 38764 3466 38792 3878
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 38948 3194 38976 6666
rect 39316 5914 39344 7142
rect 39304 5908 39356 5914
rect 39304 5850 39356 5856
rect 39120 5568 39172 5574
rect 39120 5510 39172 5516
rect 39132 5234 39160 5510
rect 39120 5228 39172 5234
rect 39120 5170 39172 5176
rect 39132 4758 39160 5170
rect 39120 4752 39172 4758
rect 39120 4694 39172 4700
rect 39316 4282 39344 5850
rect 39408 4690 39436 7686
rect 39396 4684 39448 4690
rect 39396 4626 39448 4632
rect 39304 4276 39356 4282
rect 39304 4218 39356 4224
rect 38936 3188 38988 3194
rect 38936 3130 38988 3136
rect 39316 3126 39344 4218
rect 39500 3398 39528 8842
rect 40144 6730 40172 9318
rect 40420 8498 40448 10390
rect 40500 9920 40552 9926
rect 40500 9862 40552 9868
rect 40512 9586 40540 9862
rect 40500 9580 40552 9586
rect 40500 9522 40552 9528
rect 40604 9466 40632 12406
rect 40776 12378 40828 12384
rect 40868 11688 40920 11694
rect 40868 11630 40920 11636
rect 40880 10810 40908 11630
rect 40868 10804 40920 10810
rect 40868 10746 40920 10752
rect 40776 10464 40828 10470
rect 40776 10406 40828 10412
rect 40788 10130 40816 10406
rect 40776 10124 40828 10130
rect 40776 10066 40828 10072
rect 40972 9722 41000 12718
rect 41616 11898 41644 12922
rect 42352 12442 42380 13194
rect 42444 12646 42472 14418
rect 42536 13190 42564 17274
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 42812 15910 42840 17138
rect 43076 16448 43128 16454
rect 43076 16390 43128 16396
rect 42984 16108 43036 16114
rect 42984 16050 43036 16056
rect 42800 15904 42852 15910
rect 42800 15846 42852 15852
rect 42616 15564 42668 15570
rect 42616 15506 42668 15512
rect 42524 13184 42576 13190
rect 42524 13126 42576 13132
rect 42536 12918 42564 13126
rect 42524 12912 42576 12918
rect 42524 12854 42576 12860
rect 42628 12764 42656 15506
rect 42812 15366 42840 15846
rect 42800 15360 42852 15366
rect 42800 15302 42852 15308
rect 42708 14476 42760 14482
rect 42708 14418 42760 14424
rect 42720 13870 42748 14418
rect 42812 14346 42840 15302
rect 42996 15162 43024 16050
rect 42984 15156 43036 15162
rect 42984 15098 43036 15104
rect 43088 15026 43116 16390
rect 43076 15020 43128 15026
rect 43076 14962 43128 14968
rect 43180 14906 43208 18022
rect 43260 17604 43312 17610
rect 43260 17546 43312 17552
rect 43272 15638 43300 17546
rect 43812 16992 43864 16998
rect 43812 16934 43864 16940
rect 43824 16794 43852 16934
rect 43812 16788 43864 16794
rect 43812 16730 43864 16736
rect 43260 15632 43312 15638
rect 43260 15574 43312 15580
rect 43088 14878 43208 14906
rect 43352 14952 43404 14958
rect 43352 14894 43404 14900
rect 42800 14340 42852 14346
rect 42800 14282 42852 14288
rect 42892 14272 42944 14278
rect 42892 14214 42944 14220
rect 42708 13864 42760 13870
rect 42708 13806 42760 13812
rect 42536 12736 42656 12764
rect 42432 12640 42484 12646
rect 42432 12582 42484 12588
rect 42340 12436 42392 12442
rect 42536 12434 42564 12736
rect 42616 12640 42668 12646
rect 42616 12582 42668 12588
rect 42340 12378 42392 12384
rect 42444 12406 42564 12434
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 41604 11892 41656 11898
rect 41604 11834 41656 11840
rect 41616 11218 41644 11834
rect 41604 11212 41656 11218
rect 41604 11154 41656 11160
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 41340 10810 41368 11086
rect 41800 11082 41828 12038
rect 42156 11552 42208 11558
rect 42156 11494 42208 11500
rect 42064 11212 42116 11218
rect 42064 11154 42116 11160
rect 41788 11076 41840 11082
rect 41788 11018 41840 11024
rect 41328 10804 41380 10810
rect 41328 10746 41380 10752
rect 41328 10600 41380 10606
rect 41328 10542 41380 10548
rect 41340 9994 41368 10542
rect 41328 9988 41380 9994
rect 41328 9930 41380 9936
rect 41340 9722 41368 9930
rect 40960 9716 41012 9722
rect 40960 9658 41012 9664
rect 41328 9716 41380 9722
rect 41328 9658 41380 9664
rect 40512 9438 40632 9466
rect 40408 8492 40460 8498
rect 40408 8434 40460 8440
rect 40512 8362 40540 9438
rect 40224 8356 40276 8362
rect 40224 8298 40276 8304
rect 40500 8356 40552 8362
rect 40500 8298 40552 8304
rect 40132 6724 40184 6730
rect 40132 6666 40184 6672
rect 40040 6656 40092 6662
rect 40040 6598 40092 6604
rect 39672 6316 39724 6322
rect 39672 6258 39724 6264
rect 39948 6316 40000 6322
rect 39948 6258 40000 6264
rect 39684 5914 39712 6258
rect 39672 5908 39724 5914
rect 39672 5850 39724 5856
rect 39960 5166 39988 6258
rect 40052 5710 40080 6598
rect 40144 6390 40172 6666
rect 40132 6384 40184 6390
rect 40132 6326 40184 6332
rect 40144 5914 40172 6326
rect 40132 5908 40184 5914
rect 40132 5850 40184 5856
rect 40040 5704 40092 5710
rect 40040 5646 40092 5652
rect 39948 5160 40000 5166
rect 39948 5102 40000 5108
rect 39672 4616 39724 4622
rect 39672 4558 39724 4564
rect 39580 3936 39632 3942
rect 39578 3904 39580 3913
rect 39632 3904 39634 3913
rect 39578 3839 39634 3848
rect 39396 3392 39448 3398
rect 39396 3334 39448 3340
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39408 3194 39436 3334
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39304 3120 39356 3126
rect 39304 3062 39356 3068
rect 39212 3052 39264 3058
rect 39212 2994 39264 3000
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38568 2644 38620 2650
rect 38568 2586 38620 2592
rect 38672 2514 38700 2790
rect 39224 2650 39252 2994
rect 39684 2774 39712 4558
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 40144 4214 40172 4490
rect 40132 4208 40184 4214
rect 40132 4150 40184 4156
rect 39764 4140 39816 4146
rect 39764 4082 39816 4088
rect 39776 3738 39804 4082
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39764 3732 39816 3738
rect 39764 3674 39816 3680
rect 39960 3720 39988 4014
rect 40040 3732 40092 3738
rect 39960 3692 40040 3720
rect 39764 2848 39816 2854
rect 39764 2790 39816 2796
rect 39592 2746 39712 2774
rect 39212 2644 39264 2650
rect 39212 2586 39264 2592
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 39028 2508 39080 2514
rect 39028 2450 39080 2456
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38764 1442 38792 2382
rect 38488 1414 38792 1442
rect 38488 800 38516 1414
rect 39040 800 39068 2450
rect 39592 800 39620 2746
rect 39776 2632 39804 2790
rect 39684 2604 39804 2632
rect 39684 2446 39712 2604
rect 39960 2446 39988 3692
rect 40040 3674 40092 3680
rect 40132 3460 40184 3466
rect 40132 3402 40184 3408
rect 40144 2650 40172 3402
rect 40236 3058 40264 8298
rect 41340 8276 41368 9658
rect 41800 9654 41828 11018
rect 41972 11008 42024 11014
rect 41972 10950 42024 10956
rect 41984 10538 42012 10950
rect 42076 10674 42104 11154
rect 42064 10668 42116 10674
rect 42064 10610 42116 10616
rect 41972 10532 42024 10538
rect 41972 10474 42024 10480
rect 41984 10130 42012 10474
rect 42168 10266 42196 11494
rect 42444 10282 42472 12406
rect 42628 12170 42656 12582
rect 42616 12164 42668 12170
rect 42616 12106 42668 12112
rect 42628 10810 42656 12106
rect 42616 10804 42668 10810
rect 42616 10746 42668 10752
rect 42720 10470 42748 13806
rect 42904 12306 42932 14214
rect 42984 13864 43036 13870
rect 42984 13806 43036 13812
rect 42996 12986 43024 13806
rect 42984 12980 43036 12986
rect 42984 12922 43036 12928
rect 42996 12442 43024 12922
rect 43088 12782 43116 14878
rect 43364 13462 43392 14894
rect 43812 14816 43864 14822
rect 43812 14758 43864 14764
rect 43536 14408 43588 14414
rect 43536 14350 43588 14356
rect 43444 14272 43496 14278
rect 43444 14214 43496 14220
rect 43352 13456 43404 13462
rect 43352 13398 43404 13404
rect 43168 13184 43220 13190
rect 43168 13126 43220 13132
rect 43076 12776 43128 12782
rect 43076 12718 43128 12724
rect 42984 12436 43036 12442
rect 42984 12378 43036 12384
rect 42892 12300 42944 12306
rect 42892 12242 42944 12248
rect 43088 12102 43116 12718
rect 43180 12306 43208 13126
rect 43456 12986 43484 14214
rect 43548 14074 43576 14350
rect 43824 14346 43852 14758
rect 43904 14476 43956 14482
rect 43904 14418 43956 14424
rect 43812 14340 43864 14346
rect 43812 14282 43864 14288
rect 43536 14068 43588 14074
rect 43536 14010 43588 14016
rect 43628 14068 43680 14074
rect 43628 14010 43680 14016
rect 43640 13802 43668 14010
rect 43824 13938 43852 14282
rect 43916 13938 43944 14418
rect 43812 13932 43864 13938
rect 43812 13874 43864 13880
rect 43904 13932 43956 13938
rect 44008 13920 44036 20266
rect 44192 19514 44220 20878
rect 44652 20806 44680 21830
rect 44640 20800 44692 20806
rect 44640 20742 44692 20748
rect 44282 20700 44590 20709
rect 44282 20698 44288 20700
rect 44344 20698 44368 20700
rect 44424 20698 44448 20700
rect 44504 20698 44528 20700
rect 44584 20698 44590 20700
rect 44344 20646 44346 20698
rect 44526 20646 44528 20698
rect 44282 20644 44288 20646
rect 44344 20644 44368 20646
rect 44424 20644 44448 20646
rect 44504 20644 44528 20646
rect 44584 20644 44590 20646
rect 44282 20635 44590 20644
rect 44652 20398 44680 20742
rect 44744 20602 44772 22918
rect 44928 22574 44956 25298
rect 45008 25152 45060 25158
rect 45008 25094 45060 25100
rect 45020 24818 45048 25094
rect 45388 24818 45416 26250
rect 45480 25974 45508 26794
rect 45836 26784 45888 26790
rect 45836 26726 45888 26732
rect 45744 26240 45796 26246
rect 45744 26182 45796 26188
rect 45468 25968 45520 25974
rect 45468 25910 45520 25916
rect 45652 25900 45704 25906
rect 45652 25842 45704 25848
rect 45664 25226 45692 25842
rect 45756 25838 45784 26182
rect 45848 26042 45876 26726
rect 46308 26042 46336 26862
rect 46572 26376 46624 26382
rect 46572 26318 46624 26324
rect 46388 26240 46440 26246
rect 46388 26182 46440 26188
rect 45836 26036 45888 26042
rect 45836 25978 45888 25984
rect 46296 26036 46348 26042
rect 46296 25978 46348 25984
rect 45744 25832 45796 25838
rect 45744 25774 45796 25780
rect 45756 25537 45784 25774
rect 45742 25528 45798 25537
rect 45848 25498 45876 25978
rect 46020 25696 46072 25702
rect 46020 25638 46072 25644
rect 45742 25463 45798 25472
rect 45836 25492 45888 25498
rect 45836 25434 45888 25440
rect 46032 25430 46060 25638
rect 46020 25424 46072 25430
rect 46020 25366 46072 25372
rect 45928 25356 45980 25362
rect 45928 25298 45980 25304
rect 45652 25220 45704 25226
rect 45652 25162 45704 25168
rect 45008 24812 45060 24818
rect 45008 24754 45060 24760
rect 45376 24812 45428 24818
rect 45376 24754 45428 24760
rect 45664 23866 45692 25162
rect 45940 24954 45968 25298
rect 45928 24948 45980 24954
rect 45928 24890 45980 24896
rect 46400 24818 46428 26182
rect 46584 25974 46612 26318
rect 46676 26042 46704 26862
rect 47308 26784 47360 26790
rect 47308 26726 47360 26732
rect 47584 26784 47636 26790
rect 47584 26726 47636 26732
rect 47320 26382 47348 26726
rect 47308 26376 47360 26382
rect 47308 26318 47360 26324
rect 46848 26240 46900 26246
rect 46848 26182 46900 26188
rect 46860 26042 46888 26182
rect 47596 26042 47624 26726
rect 48148 26586 48176 26862
rect 48228 26852 48280 26858
rect 48228 26794 48280 26800
rect 48136 26580 48188 26586
rect 48136 26522 48188 26528
rect 48240 26382 48268 26794
rect 48780 26784 48832 26790
rect 48780 26726 48832 26732
rect 48792 26518 48820 26726
rect 48780 26512 48832 26518
rect 48780 26454 48832 26460
rect 48228 26376 48280 26382
rect 48228 26318 48280 26324
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 46664 26036 46716 26042
rect 46664 25978 46716 25984
rect 46848 26036 46900 26042
rect 46848 25978 46900 25984
rect 47584 26036 47636 26042
rect 47584 25978 47636 25984
rect 46572 25968 46624 25974
rect 46572 25910 46624 25916
rect 46860 25906 46888 25978
rect 46848 25900 46900 25906
rect 46848 25842 46900 25848
rect 46664 25832 46716 25838
rect 46664 25774 46716 25780
rect 46388 24812 46440 24818
rect 46388 24754 46440 24760
rect 46676 24682 46704 25774
rect 46768 25622 46980 25650
rect 46768 25294 46796 25622
rect 46952 25498 46980 25622
rect 46848 25492 46900 25498
rect 46848 25434 46900 25440
rect 46940 25492 46992 25498
rect 46940 25434 46992 25440
rect 46860 25294 46888 25434
rect 47596 25362 47624 25978
rect 48148 25906 48176 26250
rect 48136 25900 48188 25906
rect 48136 25842 48188 25848
rect 48240 25362 48268 26318
rect 48596 26240 48648 26246
rect 48596 26182 48648 26188
rect 48608 25906 48636 26182
rect 48596 25900 48648 25906
rect 48596 25842 48648 25848
rect 48792 25702 48820 26454
rect 49252 26042 49280 26862
rect 50252 26784 50304 26790
rect 50252 26726 50304 26732
rect 50712 26784 50764 26790
rect 50712 26726 50764 26732
rect 49884 26376 49936 26382
rect 49884 26318 49936 26324
rect 49240 26036 49292 26042
rect 49240 25978 49292 25984
rect 49896 25906 49924 26318
rect 50264 25974 50292 26726
rect 50724 26314 50752 26726
rect 50712 26308 50764 26314
rect 50712 26250 50764 26256
rect 50252 25968 50304 25974
rect 50252 25910 50304 25916
rect 49884 25900 49936 25906
rect 49884 25842 49936 25848
rect 48780 25696 48832 25702
rect 48780 25638 48832 25644
rect 47584 25356 47636 25362
rect 47584 25298 47636 25304
rect 48228 25356 48280 25362
rect 48228 25298 48280 25304
rect 46756 25288 46808 25294
rect 46756 25230 46808 25236
rect 46848 25288 46900 25294
rect 48792 25242 48820 25638
rect 49882 25528 49938 25537
rect 50816 25498 50844 26862
rect 51092 26042 51120 26862
rect 51368 26586 51396 27406
rect 51908 27328 51960 27334
rect 51908 27270 51960 27276
rect 51504 26684 51812 26693
rect 51504 26682 51510 26684
rect 51566 26682 51590 26684
rect 51646 26682 51670 26684
rect 51726 26682 51750 26684
rect 51806 26682 51812 26684
rect 51566 26630 51568 26682
rect 51748 26630 51750 26682
rect 51504 26628 51510 26630
rect 51566 26628 51590 26630
rect 51646 26628 51670 26630
rect 51726 26628 51750 26630
rect 51806 26628 51812 26630
rect 51504 26619 51812 26628
rect 51356 26580 51408 26586
rect 51356 26522 51408 26528
rect 51356 26240 51408 26246
rect 51356 26182 51408 26188
rect 51080 26036 51132 26042
rect 51080 25978 51132 25984
rect 50896 25900 50948 25906
rect 50896 25842 50948 25848
rect 50908 25498 50936 25842
rect 51368 25838 51396 26182
rect 51920 25906 51948 27270
rect 58726 27228 59034 27237
rect 58726 27226 58732 27228
rect 58788 27226 58812 27228
rect 58868 27226 58892 27228
rect 58948 27226 58972 27228
rect 59028 27226 59034 27228
rect 58788 27174 58790 27226
rect 58970 27174 58972 27226
rect 58726 27172 58732 27174
rect 58788 27172 58812 27174
rect 58868 27172 58892 27174
rect 58948 27172 58972 27174
rect 59028 27172 59034 27174
rect 58726 27163 59034 27172
rect 52000 26920 52052 26926
rect 54668 26920 54720 26926
rect 52000 26862 52052 26868
rect 54496 26880 54668 26908
rect 52012 26042 52040 26862
rect 52092 26784 52144 26790
rect 52092 26726 52144 26732
rect 53840 26784 53892 26790
rect 53840 26726 53892 26732
rect 52000 26036 52052 26042
rect 52000 25978 52052 25984
rect 51908 25900 51960 25906
rect 51908 25842 51960 25848
rect 51264 25832 51316 25838
rect 51264 25774 51316 25780
rect 51356 25832 51408 25838
rect 51356 25774 51408 25780
rect 52000 25832 52052 25838
rect 52000 25774 52052 25780
rect 49882 25463 49884 25472
rect 49936 25463 49938 25472
rect 50804 25492 50856 25498
rect 49884 25434 49936 25440
rect 50804 25434 50856 25440
rect 50896 25492 50948 25498
rect 50896 25434 50948 25440
rect 50908 25378 50936 25434
rect 46848 25230 46900 25236
rect 46664 24676 46716 24682
rect 46664 24618 46716 24624
rect 46676 24410 46704 24618
rect 46664 24404 46716 24410
rect 46664 24346 46716 24352
rect 46768 24290 46796 25230
rect 48700 25214 48820 25242
rect 50816 25350 50936 25378
rect 48044 25152 48096 25158
rect 48044 25094 48096 25100
rect 47492 24608 47544 24614
rect 47492 24550 47544 24556
rect 46768 24262 46888 24290
rect 46480 24200 46532 24206
rect 46480 24142 46532 24148
rect 46756 24200 46808 24206
rect 46756 24142 46808 24148
rect 45928 24064 45980 24070
rect 45928 24006 45980 24012
rect 45652 23860 45704 23866
rect 45652 23802 45704 23808
rect 45284 23656 45336 23662
rect 45284 23598 45336 23604
rect 45296 23526 45324 23598
rect 45100 23520 45152 23526
rect 45100 23462 45152 23468
rect 45284 23520 45336 23526
rect 45284 23462 45336 23468
rect 45008 23112 45060 23118
rect 45008 23054 45060 23060
rect 44916 22568 44968 22574
rect 44916 22510 44968 22516
rect 45020 22438 45048 23054
rect 45112 22710 45140 23462
rect 45296 23322 45324 23462
rect 45284 23316 45336 23322
rect 45336 23276 45416 23304
rect 45284 23258 45336 23264
rect 45100 22704 45152 22710
rect 45100 22646 45152 22652
rect 45008 22432 45060 22438
rect 45008 22374 45060 22380
rect 45020 22094 45048 22374
rect 44836 22066 45048 22094
rect 44836 21078 44864 22066
rect 44824 21072 44876 21078
rect 44824 21014 44876 21020
rect 44732 20596 44784 20602
rect 44732 20538 44784 20544
rect 44456 20392 44508 20398
rect 44456 20334 44508 20340
rect 44640 20392 44692 20398
rect 44640 20334 44692 20340
rect 44468 19718 44496 20334
rect 44836 20330 44864 21014
rect 45284 20392 45336 20398
rect 45284 20334 45336 20340
rect 44824 20324 44876 20330
rect 44824 20266 44876 20272
rect 45100 20256 45152 20262
rect 45100 20198 45152 20204
rect 44916 19916 44968 19922
rect 44916 19858 44968 19864
rect 44456 19712 44508 19718
rect 44456 19654 44508 19660
rect 44282 19612 44590 19621
rect 44282 19610 44288 19612
rect 44344 19610 44368 19612
rect 44424 19610 44448 19612
rect 44504 19610 44528 19612
rect 44584 19610 44590 19612
rect 44344 19558 44346 19610
rect 44526 19558 44528 19610
rect 44282 19556 44288 19558
rect 44344 19556 44368 19558
rect 44424 19556 44448 19558
rect 44504 19556 44528 19558
rect 44584 19556 44590 19558
rect 44282 19547 44590 19556
rect 44180 19508 44232 19514
rect 44180 19450 44232 19456
rect 44640 19168 44692 19174
rect 44640 19110 44692 19116
rect 44652 18834 44680 19110
rect 44928 18850 44956 19858
rect 45008 19848 45060 19854
rect 45008 19790 45060 19796
rect 45020 19310 45048 19790
rect 45112 19310 45140 20198
rect 45296 20058 45324 20334
rect 45284 20052 45336 20058
rect 45284 19994 45336 20000
rect 45008 19304 45060 19310
rect 45008 19246 45060 19252
rect 45100 19304 45152 19310
rect 45100 19246 45152 19252
rect 45020 18970 45048 19246
rect 45008 18964 45060 18970
rect 45008 18906 45060 18912
rect 44640 18828 44692 18834
rect 44928 18822 45048 18850
rect 44640 18770 44692 18776
rect 44282 18524 44590 18533
rect 44282 18522 44288 18524
rect 44344 18522 44368 18524
rect 44424 18522 44448 18524
rect 44504 18522 44528 18524
rect 44584 18522 44590 18524
rect 44344 18470 44346 18522
rect 44526 18470 44528 18522
rect 44282 18468 44288 18470
rect 44344 18468 44368 18470
rect 44424 18468 44448 18470
rect 44504 18468 44528 18470
rect 44584 18468 44590 18470
rect 44282 18459 44590 18468
rect 44640 18216 44692 18222
rect 44640 18158 44692 18164
rect 44088 18080 44140 18086
rect 44088 18022 44140 18028
rect 44180 18080 44232 18086
rect 44180 18022 44232 18028
rect 44100 16590 44128 18022
rect 44192 17542 44220 18022
rect 44180 17536 44232 17542
rect 44180 17478 44232 17484
rect 44192 17134 44220 17478
rect 44282 17436 44590 17445
rect 44282 17434 44288 17436
rect 44344 17434 44368 17436
rect 44424 17434 44448 17436
rect 44504 17434 44528 17436
rect 44584 17434 44590 17436
rect 44344 17382 44346 17434
rect 44526 17382 44528 17434
rect 44282 17380 44288 17382
rect 44344 17380 44368 17382
rect 44424 17380 44448 17382
rect 44504 17380 44528 17382
rect 44584 17380 44590 17382
rect 44282 17371 44590 17380
rect 44652 17338 44680 18158
rect 44824 17672 44876 17678
rect 44824 17614 44876 17620
rect 44732 17536 44784 17542
rect 44732 17478 44784 17484
rect 44640 17332 44692 17338
rect 44640 17274 44692 17280
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 44088 16584 44140 16590
rect 44088 16526 44140 16532
rect 44282 16348 44590 16357
rect 44282 16346 44288 16348
rect 44344 16346 44368 16348
rect 44424 16346 44448 16348
rect 44504 16346 44528 16348
rect 44584 16346 44590 16348
rect 44344 16294 44346 16346
rect 44526 16294 44528 16346
rect 44282 16292 44288 16294
rect 44344 16292 44368 16294
rect 44424 16292 44448 16294
rect 44504 16292 44528 16294
rect 44584 16292 44590 16294
rect 44282 16283 44590 16292
rect 44100 16114 44312 16130
rect 44100 16108 44324 16114
rect 44100 16102 44272 16108
rect 44100 15162 44128 16102
rect 44272 16050 44324 16056
rect 44180 16040 44232 16046
rect 44180 15982 44232 15988
rect 44640 16040 44692 16046
rect 44744 16028 44772 17478
rect 44836 16726 44864 17614
rect 44824 16720 44876 16726
rect 44824 16662 44876 16668
rect 44692 16000 44772 16028
rect 44640 15982 44692 15988
rect 44192 15570 44220 15982
rect 44180 15564 44232 15570
rect 44180 15506 44232 15512
rect 44652 15502 44680 15982
rect 44824 15972 44876 15978
rect 44824 15914 44876 15920
rect 44836 15638 44864 15914
rect 44824 15632 44876 15638
rect 44824 15574 44876 15580
rect 44640 15496 44692 15502
rect 44640 15438 44692 15444
rect 44282 15260 44590 15269
rect 44282 15258 44288 15260
rect 44344 15258 44368 15260
rect 44424 15258 44448 15260
rect 44504 15258 44528 15260
rect 44584 15258 44590 15260
rect 44344 15206 44346 15258
rect 44526 15206 44528 15258
rect 44282 15204 44288 15206
rect 44344 15204 44368 15206
rect 44424 15204 44448 15206
rect 44504 15204 44528 15206
rect 44584 15204 44590 15206
rect 44282 15195 44590 15204
rect 44088 15156 44140 15162
rect 44088 15098 44140 15104
rect 45020 14822 45048 18822
rect 45008 14816 45060 14822
rect 45008 14758 45060 14764
rect 44282 14172 44590 14181
rect 44282 14170 44288 14172
rect 44344 14170 44368 14172
rect 44424 14170 44448 14172
rect 44504 14170 44528 14172
rect 44584 14170 44590 14172
rect 44344 14118 44346 14170
rect 44526 14118 44528 14170
rect 44282 14116 44288 14118
rect 44344 14116 44368 14118
rect 44424 14116 44448 14118
rect 44504 14116 44528 14118
rect 44584 14116 44590 14118
rect 44282 14107 44590 14116
rect 45020 14074 45048 14758
rect 45008 14068 45060 14074
rect 45008 14010 45060 14016
rect 44088 13932 44140 13938
rect 44008 13892 44088 13920
rect 43904 13874 43956 13880
rect 44088 13874 44140 13880
rect 43628 13796 43680 13802
rect 43628 13738 43680 13744
rect 44100 13734 44128 13874
rect 45008 13864 45060 13870
rect 45008 13806 45060 13812
rect 44088 13728 44140 13734
rect 44088 13670 44140 13676
rect 44640 13320 44692 13326
rect 44640 13262 44692 13268
rect 44282 13084 44590 13093
rect 44282 13082 44288 13084
rect 44344 13082 44368 13084
rect 44424 13082 44448 13084
rect 44504 13082 44528 13084
rect 44584 13082 44590 13084
rect 44344 13030 44346 13082
rect 44526 13030 44528 13082
rect 44282 13028 44288 13030
rect 44344 13028 44368 13030
rect 44424 13028 44448 13030
rect 44504 13028 44528 13030
rect 44584 13028 44590 13030
rect 44282 13019 44590 13028
rect 43444 12980 43496 12986
rect 43444 12922 43496 12928
rect 43720 12912 43772 12918
rect 43720 12854 43772 12860
rect 43168 12300 43220 12306
rect 43168 12242 43220 12248
rect 43076 12096 43128 12102
rect 43076 12038 43128 12044
rect 42984 11688 43036 11694
rect 42984 11630 43036 11636
rect 42800 11552 42852 11558
rect 42800 11494 42852 11500
rect 42708 10464 42760 10470
rect 42708 10406 42760 10412
rect 42156 10260 42208 10266
rect 42156 10202 42208 10208
rect 42260 10254 42472 10282
rect 42168 10130 42196 10202
rect 41972 10124 42024 10130
rect 41972 10066 42024 10072
rect 42156 10124 42208 10130
rect 42156 10066 42208 10072
rect 41880 10056 41932 10062
rect 41880 9998 41932 10004
rect 41788 9648 41840 9654
rect 41788 9590 41840 9596
rect 41604 9376 41656 9382
rect 41892 9364 41920 9998
rect 42260 9674 42288 10254
rect 42432 10124 42484 10130
rect 42432 10066 42484 10072
rect 41656 9336 41920 9364
rect 41984 9646 42288 9674
rect 41604 9318 41656 9324
rect 41340 8248 41460 8276
rect 41052 7880 41104 7886
rect 41052 7822 41104 7828
rect 40960 7812 41012 7818
rect 40960 7754 41012 7760
rect 40500 7744 40552 7750
rect 40500 7686 40552 7692
rect 40512 7546 40540 7686
rect 40972 7546 41000 7754
rect 41064 7546 41092 7822
rect 41432 7546 41460 8248
rect 41512 7880 41564 7886
rect 41512 7822 41564 7828
rect 40500 7540 40552 7546
rect 40500 7482 40552 7488
rect 40960 7540 41012 7546
rect 40960 7482 41012 7488
rect 41052 7540 41104 7546
rect 41052 7482 41104 7488
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 41052 7336 41104 7342
rect 41052 7278 41104 7284
rect 41064 7002 41092 7278
rect 41052 6996 41104 7002
rect 41052 6938 41104 6944
rect 40408 6656 40460 6662
rect 40408 6598 40460 6604
rect 40420 6458 40448 6598
rect 40408 6452 40460 6458
rect 40408 6394 40460 6400
rect 41064 6186 41092 6938
rect 41432 6746 41460 7482
rect 41340 6730 41460 6746
rect 41328 6724 41460 6730
rect 41380 6718 41460 6724
rect 41328 6666 41380 6672
rect 41432 6186 41460 6718
rect 41052 6180 41104 6186
rect 41052 6122 41104 6128
rect 41420 6180 41472 6186
rect 41420 6122 41472 6128
rect 41524 5778 41552 7822
rect 41616 6746 41644 9318
rect 41788 7744 41840 7750
rect 41788 7686 41840 7692
rect 41800 7410 41828 7686
rect 41788 7404 41840 7410
rect 41788 7346 41840 7352
rect 41696 7336 41748 7342
rect 41696 7278 41748 7284
rect 41708 7206 41736 7278
rect 41696 7200 41748 7206
rect 41984 7188 42012 9646
rect 42444 9518 42472 10066
rect 42432 9512 42484 9518
rect 42432 9454 42484 9460
rect 42248 9036 42300 9042
rect 42248 8978 42300 8984
rect 42064 8288 42116 8294
rect 42064 8230 42116 8236
rect 42076 7478 42104 8230
rect 42260 7478 42288 8978
rect 42432 8288 42484 8294
rect 42432 8230 42484 8236
rect 42444 7818 42472 8230
rect 42432 7812 42484 7818
rect 42432 7754 42484 7760
rect 42340 7744 42392 7750
rect 42340 7686 42392 7692
rect 42064 7472 42116 7478
rect 42064 7414 42116 7420
rect 42248 7472 42300 7478
rect 42248 7414 42300 7420
rect 42064 7200 42116 7206
rect 41984 7160 42064 7188
rect 41696 7142 41748 7148
rect 42064 7142 42116 7148
rect 41972 6860 42024 6866
rect 41972 6802 42024 6808
rect 41880 6792 41932 6798
rect 41800 6752 41880 6780
rect 41800 6746 41828 6752
rect 41616 6718 41828 6746
rect 41880 6734 41932 6740
rect 41708 5846 41736 6718
rect 41984 6458 42012 6802
rect 42156 6792 42208 6798
rect 42352 6780 42380 7686
rect 42524 7472 42576 7478
rect 42524 7414 42576 7420
rect 42432 6860 42484 6866
rect 42432 6802 42484 6808
rect 42208 6752 42380 6780
rect 42156 6734 42208 6740
rect 41972 6452 42024 6458
rect 41972 6394 42024 6400
rect 42444 6390 42472 6802
rect 42536 6662 42564 7414
rect 42812 6882 42840 11494
rect 42996 11354 43024 11630
rect 43732 11558 43760 12854
rect 44088 12640 44140 12646
rect 44088 12582 44140 12588
rect 44100 12306 44128 12582
rect 44088 12300 44140 12306
rect 44088 12242 44140 12248
rect 44652 12238 44680 13262
rect 45020 13258 45048 13806
rect 44732 13252 44784 13258
rect 44732 13194 44784 13200
rect 45008 13252 45060 13258
rect 45008 13194 45060 13200
rect 44744 12442 44772 13194
rect 44732 12436 44784 12442
rect 44732 12378 44784 12384
rect 45112 12374 45140 19246
rect 45388 18086 45416 23276
rect 45468 23112 45520 23118
rect 45468 23054 45520 23060
rect 45480 22642 45508 23054
rect 45940 23050 45968 24006
rect 46492 23866 46520 24142
rect 46480 23860 46532 23866
rect 46480 23802 46532 23808
rect 46572 23724 46624 23730
rect 46572 23666 46624 23672
rect 45560 23044 45612 23050
rect 45560 22986 45612 22992
rect 45928 23044 45980 23050
rect 45928 22986 45980 22992
rect 45572 22710 45600 22986
rect 45560 22704 45612 22710
rect 45560 22646 45612 22652
rect 45468 22636 45520 22642
rect 45468 22578 45520 22584
rect 45572 20806 45600 22646
rect 46204 22636 46256 22642
rect 46204 22578 46256 22584
rect 46216 21690 46244 22578
rect 46388 22092 46440 22098
rect 46584 22094 46612 23666
rect 46664 23656 46716 23662
rect 46664 23598 46716 23604
rect 46676 23066 46704 23598
rect 46768 23322 46796 24142
rect 46756 23316 46808 23322
rect 46756 23258 46808 23264
rect 46860 23202 46888 24262
rect 47400 24064 47452 24070
rect 47400 24006 47452 24012
rect 46860 23174 46980 23202
rect 46676 23038 46796 23066
rect 46584 22066 46704 22094
rect 46388 22034 46440 22040
rect 46204 21684 46256 21690
rect 46204 21626 46256 21632
rect 46400 21146 46428 22034
rect 46676 21894 46704 22066
rect 46480 21888 46532 21894
rect 46480 21830 46532 21836
rect 46664 21888 46716 21894
rect 46664 21830 46716 21836
rect 46492 21554 46520 21830
rect 46480 21548 46532 21554
rect 46480 21490 46532 21496
rect 46768 21146 46796 23038
rect 46848 23044 46900 23050
rect 46848 22986 46900 22992
rect 46860 22098 46888 22986
rect 46952 22642 46980 23174
rect 47412 23118 47440 24006
rect 47504 23662 47532 24550
rect 47492 23656 47544 23662
rect 47492 23598 47544 23604
rect 47400 23112 47452 23118
rect 47400 23054 47452 23060
rect 46940 22636 46992 22642
rect 46940 22578 46992 22584
rect 47308 22432 47360 22438
rect 47308 22374 47360 22380
rect 46848 22092 46900 22098
rect 46848 22034 46900 22040
rect 46940 22024 46992 22030
rect 46940 21966 46992 21972
rect 46952 21690 46980 21966
rect 46940 21684 46992 21690
rect 46940 21626 46992 21632
rect 47320 21554 47348 22374
rect 47504 22094 47532 23598
rect 47584 22432 47636 22438
rect 47584 22374 47636 22380
rect 47412 22066 47532 22094
rect 47308 21548 47360 21554
rect 47308 21490 47360 21496
rect 46388 21140 46440 21146
rect 46388 21082 46440 21088
rect 46756 21140 46808 21146
rect 46756 21082 46808 21088
rect 45560 20800 45612 20806
rect 45560 20742 45612 20748
rect 45572 19854 45600 20742
rect 46768 20466 46796 21082
rect 46756 20460 46808 20466
rect 46756 20402 46808 20408
rect 45928 20256 45980 20262
rect 45928 20198 45980 20204
rect 46664 20256 46716 20262
rect 46664 20198 46716 20204
rect 47308 20256 47360 20262
rect 47308 20198 47360 20204
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45744 19848 45796 19854
rect 45744 19790 45796 19796
rect 45756 19378 45784 19790
rect 45940 19786 45968 20198
rect 45928 19780 45980 19786
rect 45928 19722 45980 19728
rect 45940 19514 45968 19722
rect 45928 19508 45980 19514
rect 45928 19450 45980 19456
rect 45468 19372 45520 19378
rect 45468 19314 45520 19320
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 46112 19372 46164 19378
rect 46112 19314 46164 19320
rect 45376 18080 45428 18086
rect 45376 18022 45428 18028
rect 45388 17746 45416 18022
rect 45376 17740 45428 17746
rect 45376 17682 45428 17688
rect 45284 17536 45336 17542
rect 45284 17478 45336 17484
rect 45296 17338 45324 17478
rect 45284 17332 45336 17338
rect 45284 17274 45336 17280
rect 45296 16114 45324 17274
rect 45388 17134 45416 17682
rect 45376 17128 45428 17134
rect 45376 17070 45428 17076
rect 45284 16108 45336 16114
rect 45284 16050 45336 16056
rect 45284 15904 45336 15910
rect 45284 15846 45336 15852
rect 45296 14482 45324 15846
rect 45376 14816 45428 14822
rect 45376 14758 45428 14764
rect 45284 14476 45336 14482
rect 45284 14418 45336 14424
rect 45388 13938 45416 14758
rect 45480 14362 45508 19314
rect 46124 18970 46152 19314
rect 46112 18964 46164 18970
rect 46112 18906 46164 18912
rect 46112 18828 46164 18834
rect 46112 18770 46164 18776
rect 46124 18154 46152 18770
rect 46676 18766 46704 20198
rect 47216 19916 47268 19922
rect 47216 19858 47268 19864
rect 47228 19378 47256 19858
rect 47216 19372 47268 19378
rect 47216 19314 47268 19320
rect 47320 19174 47348 20198
rect 47412 19242 47440 22066
rect 47596 22030 47624 22374
rect 48056 22098 48084 25094
rect 48136 24200 48188 24206
rect 48136 24142 48188 24148
rect 48148 23866 48176 24142
rect 48320 24064 48372 24070
rect 48320 24006 48372 24012
rect 48136 23860 48188 23866
rect 48136 23802 48188 23808
rect 48332 23594 48360 24006
rect 48504 23656 48556 23662
rect 48504 23598 48556 23604
rect 48320 23588 48372 23594
rect 48320 23530 48372 23536
rect 48332 22642 48360 23530
rect 48516 23322 48544 23598
rect 48700 23526 48728 25214
rect 50816 25158 50844 25350
rect 48780 25152 48832 25158
rect 48780 25094 48832 25100
rect 50804 25152 50856 25158
rect 50804 25094 50856 25100
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48504 23316 48556 23322
rect 48504 23258 48556 23264
rect 48792 22778 48820 25094
rect 50620 24812 50672 24818
rect 50620 24754 50672 24760
rect 50436 24064 50488 24070
rect 50436 24006 50488 24012
rect 49056 23792 49108 23798
rect 49056 23734 49108 23740
rect 48780 22772 48832 22778
rect 48780 22714 48832 22720
rect 48320 22636 48372 22642
rect 48320 22578 48372 22584
rect 48792 22506 48820 22714
rect 49068 22642 49096 23734
rect 50252 23656 50304 23662
rect 50252 23598 50304 23604
rect 50264 23526 50292 23598
rect 50252 23520 50304 23526
rect 50252 23462 50304 23468
rect 50264 23050 50292 23462
rect 50448 23050 50476 24006
rect 50252 23044 50304 23050
rect 50252 22986 50304 22992
rect 50436 23044 50488 23050
rect 50436 22986 50488 22992
rect 50632 22982 50660 24754
rect 50816 23730 50844 25094
rect 51172 24948 51224 24954
rect 51172 24890 51224 24896
rect 50988 24200 51040 24206
rect 50988 24142 51040 24148
rect 51000 23866 51028 24142
rect 50988 23860 51040 23866
rect 50988 23802 51040 23808
rect 50804 23724 50856 23730
rect 50804 23666 50856 23672
rect 50620 22976 50672 22982
rect 50620 22918 50672 22924
rect 50632 22778 50660 22918
rect 50620 22772 50672 22778
rect 50620 22714 50672 22720
rect 49056 22636 49108 22642
rect 49056 22578 49108 22584
rect 49240 22568 49292 22574
rect 49240 22510 49292 22516
rect 48780 22500 48832 22506
rect 48780 22442 48832 22448
rect 48228 22432 48280 22438
rect 48228 22374 48280 22380
rect 48044 22092 48096 22098
rect 48044 22034 48096 22040
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 48240 21690 48268 22374
rect 49252 22094 49280 22510
rect 49608 22500 49660 22506
rect 49608 22442 49660 22448
rect 49620 22137 49648 22442
rect 49068 22066 49280 22094
rect 49606 22128 49662 22137
rect 48320 21888 48372 21894
rect 48320 21830 48372 21836
rect 48964 21888 49016 21894
rect 48964 21830 49016 21836
rect 48228 21684 48280 21690
rect 48228 21626 48280 21632
rect 47492 20324 47544 20330
rect 47492 20266 47544 20272
rect 47504 19786 47532 20266
rect 47860 20256 47912 20262
rect 47860 20198 47912 20204
rect 47492 19780 47544 19786
rect 47492 19722 47544 19728
rect 47872 19378 47900 20198
rect 48332 19718 48360 21830
rect 48976 21554 49004 21830
rect 48964 21548 49016 21554
rect 48964 21490 49016 21496
rect 48596 21480 48648 21486
rect 48596 21422 48648 21428
rect 48412 21344 48464 21350
rect 48412 21286 48464 21292
rect 48424 20602 48452 21286
rect 48412 20596 48464 20602
rect 48412 20538 48464 20544
rect 48608 20058 48636 21422
rect 49068 21350 49096 22066
rect 49606 22063 49662 22072
rect 50160 22024 50212 22030
rect 50160 21966 50212 21972
rect 50068 21888 50120 21894
rect 50068 21830 50120 21836
rect 49056 21344 49108 21350
rect 49056 21286 49108 21292
rect 48596 20052 48648 20058
rect 48596 19994 48648 20000
rect 49068 19854 49096 21286
rect 49424 20528 49476 20534
rect 49424 20470 49476 20476
rect 49148 20392 49200 20398
rect 49148 20334 49200 20340
rect 49160 20058 49188 20334
rect 49148 20052 49200 20058
rect 49148 19994 49200 20000
rect 49056 19848 49108 19854
rect 49056 19790 49108 19796
rect 48320 19712 48372 19718
rect 48320 19654 48372 19660
rect 47860 19372 47912 19378
rect 47860 19314 47912 19320
rect 47400 19236 47452 19242
rect 47400 19178 47452 19184
rect 47216 19168 47268 19174
rect 47216 19110 47268 19116
rect 47308 19168 47360 19174
rect 47308 19110 47360 19116
rect 46664 18760 46716 18766
rect 46664 18702 46716 18708
rect 46480 18624 46532 18630
rect 46480 18566 46532 18572
rect 46112 18148 46164 18154
rect 46112 18090 46164 18096
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 45572 16114 45600 17138
rect 46020 16992 46072 16998
rect 46020 16934 46072 16940
rect 46032 16590 46060 16934
rect 46020 16584 46072 16590
rect 46020 16526 46072 16532
rect 45560 16108 45612 16114
rect 45560 16050 45612 16056
rect 45480 14334 45600 14362
rect 45468 14272 45520 14278
rect 45468 14214 45520 14220
rect 45480 14074 45508 14214
rect 45468 14068 45520 14074
rect 45468 14010 45520 14016
rect 45572 13954 45600 14334
rect 45744 14272 45796 14278
rect 45744 14214 45796 14220
rect 45756 14074 45784 14214
rect 45744 14068 45796 14074
rect 45744 14010 45796 14016
rect 45376 13932 45428 13938
rect 45376 13874 45428 13880
rect 45480 13926 45600 13954
rect 45836 13932 45888 13938
rect 45192 13388 45244 13394
rect 45192 13330 45244 13336
rect 45204 12850 45232 13330
rect 45388 13326 45416 13874
rect 45376 13320 45428 13326
rect 45376 13262 45428 13268
rect 45284 13184 45336 13190
rect 45284 13126 45336 13132
rect 45296 12986 45324 13126
rect 45388 12986 45416 13262
rect 45284 12980 45336 12986
rect 45284 12922 45336 12928
rect 45376 12980 45428 12986
rect 45376 12922 45428 12928
rect 45192 12844 45244 12850
rect 45192 12786 45244 12792
rect 45204 12442 45232 12786
rect 45192 12436 45244 12442
rect 45192 12378 45244 12384
rect 45100 12368 45152 12374
rect 45100 12310 45152 12316
rect 44640 12232 44692 12238
rect 44640 12174 44692 12180
rect 44282 11996 44590 12005
rect 44282 11994 44288 11996
rect 44344 11994 44368 11996
rect 44424 11994 44448 11996
rect 44504 11994 44528 11996
rect 44584 11994 44590 11996
rect 44344 11942 44346 11994
rect 44526 11942 44528 11994
rect 44282 11940 44288 11942
rect 44344 11940 44368 11942
rect 44424 11940 44448 11942
rect 44504 11940 44528 11942
rect 44584 11940 44590 11942
rect 44282 11931 44590 11940
rect 44456 11892 44508 11898
rect 44456 11834 44508 11840
rect 43720 11552 43772 11558
rect 43720 11494 43772 11500
rect 44468 11354 44496 11834
rect 44652 11354 44680 12174
rect 45100 11552 45152 11558
rect 45100 11494 45152 11500
rect 42984 11348 43036 11354
rect 42984 11290 43036 11296
rect 44456 11348 44508 11354
rect 44456 11290 44508 11296
rect 44640 11348 44692 11354
rect 44640 11290 44692 11296
rect 44180 11280 44232 11286
rect 44180 11222 44232 11228
rect 44088 11144 44140 11150
rect 44088 11086 44140 11092
rect 43904 11076 43956 11082
rect 43904 11018 43956 11024
rect 43536 11008 43588 11014
rect 43536 10950 43588 10956
rect 43548 10742 43576 10950
rect 43916 10810 43944 11018
rect 43904 10804 43956 10810
rect 43904 10746 43956 10752
rect 43536 10736 43588 10742
rect 43536 10678 43588 10684
rect 43812 10464 43864 10470
rect 43812 10406 43864 10412
rect 43260 10124 43312 10130
rect 43260 10066 43312 10072
rect 42892 9920 42944 9926
rect 42892 9862 42944 9868
rect 42904 7410 42932 9862
rect 43272 9382 43300 10066
rect 43352 10056 43404 10062
rect 43352 9998 43404 10004
rect 43364 9654 43392 9998
rect 43444 9920 43496 9926
rect 43444 9862 43496 9868
rect 43456 9722 43484 9862
rect 43444 9716 43496 9722
rect 43444 9658 43496 9664
rect 43352 9648 43404 9654
rect 43352 9590 43404 9596
rect 43824 9586 43852 10406
rect 43812 9580 43864 9586
rect 43812 9522 43864 9528
rect 44100 9450 44128 11086
rect 44192 10130 44220 11222
rect 44282 10908 44590 10917
rect 44282 10906 44288 10908
rect 44344 10906 44368 10908
rect 44424 10906 44448 10908
rect 44504 10906 44528 10908
rect 44584 10906 44590 10908
rect 44344 10854 44346 10906
rect 44526 10854 44528 10906
rect 44282 10852 44288 10854
rect 44344 10852 44368 10854
rect 44424 10852 44448 10854
rect 44504 10852 44528 10854
rect 44584 10852 44590 10854
rect 44282 10843 44590 10852
rect 44652 10674 44680 11290
rect 45112 10742 45140 11494
rect 45100 10736 45152 10742
rect 45100 10678 45152 10684
rect 44640 10668 44692 10674
rect 44640 10610 44692 10616
rect 44456 10600 44508 10606
rect 44456 10542 44508 10548
rect 44468 10266 44496 10542
rect 44456 10260 44508 10266
rect 44456 10202 44508 10208
rect 44652 10130 44680 10610
rect 44180 10124 44232 10130
rect 44180 10066 44232 10072
rect 44640 10124 44692 10130
rect 44640 10066 44692 10072
rect 45100 10124 45152 10130
rect 45100 10066 45152 10072
rect 44282 9820 44590 9829
rect 44282 9818 44288 9820
rect 44344 9818 44368 9820
rect 44424 9818 44448 9820
rect 44504 9818 44528 9820
rect 44584 9818 44590 9820
rect 44344 9766 44346 9818
rect 44526 9766 44528 9818
rect 44282 9764 44288 9766
rect 44344 9764 44368 9766
rect 44424 9764 44448 9766
rect 44504 9764 44528 9766
rect 44584 9764 44590 9766
rect 44282 9755 44590 9764
rect 45112 9722 45140 10066
rect 45100 9716 45152 9722
rect 45100 9658 45152 9664
rect 44088 9444 44140 9450
rect 44088 9386 44140 9392
rect 43260 9376 43312 9382
rect 43260 9318 43312 9324
rect 43272 9110 43300 9318
rect 43260 9104 43312 9110
rect 43260 9046 43312 9052
rect 44916 8832 44968 8838
rect 44916 8774 44968 8780
rect 44282 8732 44590 8741
rect 44282 8730 44288 8732
rect 44344 8730 44368 8732
rect 44424 8730 44448 8732
rect 44504 8730 44528 8732
rect 44584 8730 44590 8732
rect 44344 8678 44346 8730
rect 44526 8678 44528 8730
rect 44282 8676 44288 8678
rect 44344 8676 44368 8678
rect 44424 8676 44448 8678
rect 44504 8676 44528 8678
rect 44584 8676 44590 8678
rect 44282 8667 44590 8676
rect 44928 8566 44956 8774
rect 44916 8560 44968 8566
rect 44916 8502 44968 8508
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 42996 7954 43024 8434
rect 43076 8424 43128 8430
rect 43076 8366 43128 8372
rect 44732 8424 44784 8430
rect 44732 8366 44784 8372
rect 42984 7948 43036 7954
rect 42984 7890 43036 7896
rect 42984 7744 43036 7750
rect 42984 7686 43036 7692
rect 42996 7546 43024 7686
rect 43088 7546 43116 8366
rect 44180 8356 44232 8362
rect 44180 8298 44232 8304
rect 43904 8288 43956 8294
rect 43904 8230 43956 8236
rect 42984 7540 43036 7546
rect 42984 7482 43036 7488
rect 43076 7540 43128 7546
rect 43076 7482 43128 7488
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 42720 6854 42840 6882
rect 42996 6866 43024 7482
rect 43916 7342 43944 8230
rect 44192 7426 44220 8298
rect 44744 8090 44772 8366
rect 44732 8084 44784 8090
rect 44732 8026 44784 8032
rect 45296 8022 45324 12922
rect 45480 11694 45508 13926
rect 45836 13874 45888 13880
rect 45848 13530 45876 13874
rect 45836 13524 45888 13530
rect 45836 13466 45888 13472
rect 46124 13394 46152 18090
rect 46388 15972 46440 15978
rect 46388 15914 46440 15920
rect 46202 13560 46258 13569
rect 46202 13495 46258 13504
rect 46216 13462 46244 13495
rect 46204 13456 46256 13462
rect 46204 13398 46256 13404
rect 46112 13388 46164 13394
rect 46112 13330 46164 13336
rect 46124 12442 46152 13330
rect 46296 13184 46348 13190
rect 46296 13126 46348 13132
rect 45560 12436 45612 12442
rect 45560 12378 45612 12384
rect 46112 12436 46164 12442
rect 46112 12378 46164 12384
rect 45572 12170 45600 12378
rect 45560 12164 45612 12170
rect 45560 12106 45612 12112
rect 45468 11688 45520 11694
rect 45468 11630 45520 11636
rect 45652 11688 45704 11694
rect 45652 11630 45704 11636
rect 45928 11688 45980 11694
rect 45928 11630 45980 11636
rect 45560 11552 45612 11558
rect 45560 11494 45612 11500
rect 45572 11150 45600 11494
rect 45664 11354 45692 11630
rect 45652 11348 45704 11354
rect 45652 11290 45704 11296
rect 45560 11144 45612 11150
rect 45560 11086 45612 11092
rect 45652 11008 45704 11014
rect 45652 10950 45704 10956
rect 45664 10674 45692 10950
rect 45940 10810 45968 11630
rect 45928 10804 45980 10810
rect 45928 10746 45980 10752
rect 45652 10668 45704 10674
rect 45572 10628 45652 10656
rect 45376 8832 45428 8838
rect 45376 8774 45428 8780
rect 45388 8634 45416 8774
rect 45376 8628 45428 8634
rect 45376 8570 45428 8576
rect 45284 8016 45336 8022
rect 45284 7958 45336 7964
rect 45376 7880 45428 7886
rect 45374 7848 45376 7857
rect 45428 7848 45430 7857
rect 45374 7783 45430 7792
rect 45572 7750 45600 10628
rect 45652 10610 45704 10616
rect 46112 10464 46164 10470
rect 46112 10406 46164 10412
rect 45836 9988 45888 9994
rect 45836 9930 45888 9936
rect 45848 9722 45876 9930
rect 45836 9716 45888 9722
rect 45836 9658 45888 9664
rect 46124 9586 46152 10406
rect 46112 9580 46164 9586
rect 46112 9522 46164 9528
rect 46308 8974 46336 13126
rect 45652 8968 45704 8974
rect 45652 8910 45704 8916
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 44640 7744 44692 7750
rect 44640 7686 44692 7692
rect 45560 7744 45612 7750
rect 45560 7686 45612 7692
rect 44282 7644 44590 7653
rect 44282 7642 44288 7644
rect 44344 7642 44368 7644
rect 44424 7642 44448 7644
rect 44504 7642 44528 7644
rect 44584 7642 44590 7644
rect 44344 7590 44346 7642
rect 44526 7590 44528 7642
rect 44282 7588 44288 7590
rect 44344 7588 44368 7590
rect 44424 7588 44448 7590
rect 44504 7588 44528 7590
rect 44584 7588 44590 7590
rect 44282 7579 44590 7588
rect 44192 7410 44312 7426
rect 44192 7404 44324 7410
rect 44192 7398 44272 7404
rect 44272 7346 44324 7352
rect 43904 7336 43956 7342
rect 43904 7278 43956 7284
rect 43168 7200 43220 7206
rect 43168 7142 43220 7148
rect 43260 7200 43312 7206
rect 43260 7142 43312 7148
rect 42984 6860 43036 6866
rect 42524 6656 42576 6662
rect 42524 6598 42576 6604
rect 42616 6656 42668 6662
rect 42616 6598 42668 6604
rect 42432 6384 42484 6390
rect 42432 6326 42484 6332
rect 41788 6316 41840 6322
rect 41788 6258 41840 6264
rect 41696 5840 41748 5846
rect 41696 5782 41748 5788
rect 41512 5772 41564 5778
rect 41512 5714 41564 5720
rect 41524 5166 41552 5714
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41708 5302 41736 5510
rect 41696 5296 41748 5302
rect 41696 5238 41748 5244
rect 40868 5160 40920 5166
rect 40868 5102 40920 5108
rect 41512 5160 41564 5166
rect 41512 5102 41564 5108
rect 40684 5024 40736 5030
rect 40684 4966 40736 4972
rect 40696 4078 40724 4966
rect 40880 4690 40908 5102
rect 41512 5024 41564 5030
rect 41512 4966 41564 4972
rect 41604 5024 41656 5030
rect 41604 4966 41656 4972
rect 40868 4684 40920 4690
rect 40868 4626 40920 4632
rect 40684 4072 40736 4078
rect 40684 4014 40736 4020
rect 40696 3942 40724 4014
rect 40684 3936 40736 3942
rect 40684 3878 40736 3884
rect 40500 3392 40552 3398
rect 40500 3334 40552 3340
rect 40224 3052 40276 3058
rect 40224 2994 40276 3000
rect 40512 2650 40540 3334
rect 40696 3194 40724 3878
rect 40880 3602 40908 4626
rect 41524 4214 41552 4966
rect 41616 4622 41644 4966
rect 41604 4616 41656 4622
rect 41604 4558 41656 4564
rect 41512 4208 41564 4214
rect 41512 4150 41564 4156
rect 41420 4140 41472 4146
rect 41420 4082 41472 4088
rect 40868 3596 40920 3602
rect 40868 3538 40920 3544
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 41248 3194 41276 3334
rect 41432 3194 41460 4082
rect 41512 4004 41564 4010
rect 41512 3946 41564 3952
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 41420 3188 41472 3194
rect 41420 3130 41472 3136
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40132 2644 40184 2650
rect 40132 2586 40184 2592
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 40144 800 40172 2382
rect 40696 800 40724 2926
rect 41234 2816 41290 2825
rect 41234 2751 41290 2760
rect 41248 800 41276 2751
rect 41524 2650 41552 3946
rect 41800 3942 41828 6258
rect 42628 6254 42656 6598
rect 42616 6248 42668 6254
rect 42616 6190 42668 6196
rect 42628 5914 42656 6190
rect 42616 5908 42668 5914
rect 42616 5850 42668 5856
rect 42720 5574 42748 6854
rect 42984 6802 43036 6808
rect 43180 6746 43208 7142
rect 43272 6866 43300 7142
rect 43260 6860 43312 6866
rect 43260 6802 43312 6808
rect 44652 6798 44680 7686
rect 45572 7410 45600 7686
rect 45664 7546 45692 8910
rect 46296 8832 46348 8838
rect 46400 8786 46428 15914
rect 46492 12374 46520 18566
rect 47032 17128 47084 17134
rect 47032 17070 47084 17076
rect 47044 16590 47072 17070
rect 47032 16584 47084 16590
rect 47032 16526 47084 16532
rect 47228 16114 47256 19110
rect 47320 18834 47348 19110
rect 47308 18828 47360 18834
rect 47308 18770 47360 18776
rect 48412 18216 48464 18222
rect 48412 18158 48464 18164
rect 48780 18216 48832 18222
rect 48780 18158 48832 18164
rect 47860 18080 47912 18086
rect 47860 18022 47912 18028
rect 47768 17740 47820 17746
rect 47768 17682 47820 17688
rect 47676 17672 47728 17678
rect 47676 17614 47728 17620
rect 47688 17202 47716 17614
rect 47676 17196 47728 17202
rect 47676 17138 47728 17144
rect 47688 16794 47716 17138
rect 47676 16788 47728 16794
rect 47676 16730 47728 16736
rect 47216 16108 47268 16114
rect 47216 16050 47268 16056
rect 47124 15904 47176 15910
rect 47124 15846 47176 15852
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 46572 13728 46624 13734
rect 46572 13670 46624 13676
rect 46756 13728 46808 13734
rect 46756 13670 46808 13676
rect 46584 13394 46612 13670
rect 46572 13388 46624 13394
rect 46572 13330 46624 13336
rect 46768 13326 46796 13670
rect 46756 13320 46808 13326
rect 46756 13262 46808 13268
rect 46480 12368 46532 12374
rect 46532 12328 46612 12356
rect 46480 12310 46532 12316
rect 46478 12200 46534 12209
rect 46478 12135 46534 12144
rect 46492 12102 46520 12135
rect 46480 12096 46532 12102
rect 46480 12038 46532 12044
rect 46492 11354 46520 12038
rect 46480 11348 46532 11354
rect 46480 11290 46532 11296
rect 46478 11112 46534 11121
rect 46478 11047 46480 11056
rect 46532 11047 46534 11056
rect 46480 11018 46532 11024
rect 46584 11014 46612 12328
rect 46756 12232 46808 12238
rect 46756 12174 46808 12180
rect 46768 11898 46796 12174
rect 46756 11892 46808 11898
rect 46756 11834 46808 11840
rect 46940 11756 46992 11762
rect 46940 11698 46992 11704
rect 46572 11008 46624 11014
rect 46572 10950 46624 10956
rect 46664 8968 46716 8974
rect 46664 8910 46716 8916
rect 46676 8838 46704 8910
rect 46348 8780 46428 8786
rect 46296 8774 46428 8780
rect 46664 8832 46716 8838
rect 46664 8774 46716 8780
rect 46308 8758 46428 8774
rect 46308 8498 46336 8758
rect 46296 8492 46348 8498
rect 46296 8434 46348 8440
rect 46480 8288 46532 8294
rect 46480 8230 46532 8236
rect 46202 7848 46258 7857
rect 45836 7812 45888 7818
rect 46202 7783 46258 7792
rect 45836 7754 45888 7760
rect 45848 7546 45876 7754
rect 45652 7540 45704 7546
rect 45652 7482 45704 7488
rect 45836 7540 45888 7546
rect 45836 7482 45888 7488
rect 45928 7472 45980 7478
rect 45928 7414 45980 7420
rect 45560 7404 45612 7410
rect 45560 7346 45612 7352
rect 45560 7200 45612 7206
rect 45560 7142 45612 7148
rect 45572 6866 45600 7142
rect 45560 6860 45612 6866
rect 45560 6802 45612 6808
rect 44640 6792 44692 6798
rect 43180 6730 43300 6746
rect 44640 6734 44692 6740
rect 43180 6724 43312 6730
rect 43180 6718 43260 6724
rect 43260 6666 43312 6672
rect 43168 6656 43220 6662
rect 43168 6598 43220 6604
rect 42708 5568 42760 5574
rect 42708 5510 42760 5516
rect 42984 5568 43036 5574
rect 42984 5510 43036 5516
rect 42248 5024 42300 5030
rect 42248 4966 42300 4972
rect 42260 4486 42288 4966
rect 42720 4826 42748 5510
rect 42616 4820 42668 4826
rect 42616 4762 42668 4768
rect 42708 4820 42760 4826
rect 42708 4762 42760 4768
rect 42628 4706 42656 4762
rect 42628 4678 42748 4706
rect 42616 4548 42668 4554
rect 42616 4490 42668 4496
rect 42248 4480 42300 4486
rect 42248 4422 42300 4428
rect 42260 4214 42288 4422
rect 42248 4208 42300 4214
rect 42248 4150 42300 4156
rect 41972 4140 42024 4146
rect 41972 4082 42024 4088
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 41984 3398 42012 4082
rect 42628 3466 42656 4490
rect 42616 3460 42668 3466
rect 42616 3402 42668 3408
rect 42720 3398 42748 4678
rect 42996 4010 43024 5510
rect 43180 5370 43208 6598
rect 44282 6556 44590 6565
rect 44282 6554 44288 6556
rect 44344 6554 44368 6556
rect 44424 6554 44448 6556
rect 44504 6554 44528 6556
rect 44584 6554 44590 6556
rect 44344 6502 44346 6554
rect 44526 6502 44528 6554
rect 44282 6500 44288 6502
rect 44344 6500 44368 6502
rect 44424 6500 44448 6502
rect 44504 6500 44528 6502
rect 44584 6500 44590 6502
rect 44282 6491 44590 6500
rect 44548 6384 44600 6390
rect 44548 6326 44600 6332
rect 43260 6112 43312 6118
rect 43260 6054 43312 6060
rect 43272 5710 43300 6054
rect 44560 5914 44588 6326
rect 45940 6322 45968 7414
rect 46216 7002 46244 7783
rect 46388 7404 46440 7410
rect 46388 7346 46440 7352
rect 46296 7336 46348 7342
rect 46296 7278 46348 7284
rect 46204 6996 46256 7002
rect 46204 6938 46256 6944
rect 46308 6730 46336 7278
rect 46400 7002 46428 7346
rect 46492 7342 46520 8230
rect 46480 7336 46532 7342
rect 46480 7278 46532 7284
rect 46676 7188 46704 8774
rect 46756 7880 46808 7886
rect 46848 7880 46900 7886
rect 46756 7822 46808 7828
rect 46846 7848 46848 7857
rect 46900 7848 46902 7857
rect 46768 7410 46796 7822
rect 46846 7783 46902 7792
rect 46756 7404 46808 7410
rect 46756 7346 46808 7352
rect 46676 7160 46796 7188
rect 46388 6996 46440 7002
rect 46388 6938 46440 6944
rect 46296 6724 46348 6730
rect 46296 6666 46348 6672
rect 46388 6724 46440 6730
rect 46388 6666 46440 6672
rect 45928 6316 45980 6322
rect 45928 6258 45980 6264
rect 44548 5908 44600 5914
rect 44548 5850 44600 5856
rect 43260 5704 43312 5710
rect 43260 5646 43312 5652
rect 45468 5704 45520 5710
rect 45468 5646 45520 5652
rect 44180 5636 44232 5642
rect 44180 5578 44232 5584
rect 43168 5364 43220 5370
rect 43168 5306 43220 5312
rect 44192 5302 44220 5578
rect 44640 5568 44692 5574
rect 44640 5510 44692 5516
rect 44282 5468 44590 5477
rect 44282 5466 44288 5468
rect 44344 5466 44368 5468
rect 44424 5466 44448 5468
rect 44504 5466 44528 5468
rect 44584 5466 44590 5468
rect 44344 5414 44346 5466
rect 44526 5414 44528 5466
rect 44282 5412 44288 5414
rect 44344 5412 44368 5414
rect 44424 5412 44448 5414
rect 44504 5412 44528 5414
rect 44584 5412 44590 5414
rect 44282 5403 44590 5412
rect 43076 5296 43128 5302
rect 43076 5238 43128 5244
rect 44180 5296 44232 5302
rect 44180 5238 44232 5244
rect 43088 5030 43116 5238
rect 43076 5024 43128 5030
rect 43076 4966 43128 4972
rect 44652 4690 44680 5510
rect 44640 4684 44692 4690
rect 44640 4626 44692 4632
rect 43076 4616 43128 4622
rect 43076 4558 43128 4564
rect 43812 4616 43864 4622
rect 43812 4558 43864 4564
rect 44732 4616 44784 4622
rect 44732 4558 44784 4564
rect 45284 4616 45336 4622
rect 45284 4558 45336 4564
rect 43088 4078 43116 4558
rect 43536 4480 43588 4486
rect 43536 4422 43588 4428
rect 43628 4480 43680 4486
rect 43628 4422 43680 4428
rect 43720 4480 43772 4486
rect 43720 4422 43772 4428
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43442 4040 43498 4049
rect 42984 4004 43036 4010
rect 43442 3975 43498 3984
rect 42984 3946 43036 3952
rect 43456 3942 43484 3975
rect 43444 3936 43496 3942
rect 43444 3878 43496 3884
rect 43548 3534 43576 4422
rect 43168 3528 43220 3534
rect 43536 3528 43588 3534
rect 43168 3470 43220 3476
rect 43350 3496 43406 3505
rect 41972 3392 42024 3398
rect 41972 3334 42024 3340
rect 42340 3392 42392 3398
rect 42340 3334 42392 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 41788 2984 41840 2990
rect 41788 2926 41840 2932
rect 42246 2952 42302 2961
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 41800 800 41828 2926
rect 42246 2887 42302 2896
rect 42260 2446 42288 2887
rect 42352 2446 42380 3334
rect 43180 3194 43208 3470
rect 43536 3470 43588 3476
rect 43350 3431 43352 3440
rect 43404 3431 43406 3440
rect 43352 3402 43404 3408
rect 43168 3188 43220 3194
rect 43168 3130 43220 3136
rect 43640 3058 43668 4422
rect 43732 4214 43760 4422
rect 43720 4208 43772 4214
rect 43720 4150 43772 4156
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43444 2848 43496 2854
rect 43444 2790 43496 2796
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42248 2440 42300 2446
rect 42248 2382 42300 2388
rect 42340 2440 42392 2446
rect 42340 2382 42392 2388
rect 42352 870 42472 898
rect 42352 800 42380 870
rect 37476 734 37688 762
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42444 762 42472 870
rect 42628 762 42656 2450
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 42904 870 43024 898
rect 42904 800 42932 870
rect 42444 734 42656 762
rect 42890 0 42946 800
rect 42996 762 43024 870
rect 43180 762 43208 2382
rect 43456 800 43484 2790
rect 43824 2650 43852 4558
rect 44282 4380 44590 4389
rect 44282 4378 44288 4380
rect 44344 4378 44368 4380
rect 44424 4378 44448 4380
rect 44504 4378 44528 4380
rect 44584 4378 44590 4380
rect 44344 4326 44346 4378
rect 44526 4326 44528 4378
rect 44282 4324 44288 4326
rect 44344 4324 44368 4326
rect 44424 4324 44448 4326
rect 44504 4324 44528 4326
rect 44584 4324 44590 4326
rect 44282 4315 44590 4324
rect 44640 4276 44692 4282
rect 44640 4218 44692 4224
rect 44088 4004 44140 4010
rect 44088 3946 44140 3952
rect 43904 3936 43956 3942
rect 43904 3878 43956 3884
rect 43916 3641 43944 3878
rect 44100 3754 44128 3946
rect 44180 3936 44232 3942
rect 44178 3904 44180 3913
rect 44232 3904 44234 3913
rect 44652 3890 44680 4218
rect 44744 4078 44772 4558
rect 45100 4480 45152 4486
rect 45100 4422 45152 4428
rect 44824 4276 44876 4282
rect 44824 4218 44876 4224
rect 44732 4072 44784 4078
rect 44732 4014 44784 4020
rect 44652 3862 44772 3890
rect 44178 3839 44234 3848
rect 44100 3726 44220 3754
rect 43902 3632 43958 3641
rect 43902 3567 43958 3576
rect 43996 2984 44048 2990
rect 43996 2926 44048 2932
rect 43812 2644 43864 2650
rect 43812 2586 43864 2592
rect 44008 800 44036 2926
rect 44192 2650 44220 3726
rect 44640 3528 44692 3534
rect 44640 3470 44692 3476
rect 44282 3292 44590 3301
rect 44282 3290 44288 3292
rect 44344 3290 44368 3292
rect 44424 3290 44448 3292
rect 44504 3290 44528 3292
rect 44584 3290 44590 3292
rect 44344 3238 44346 3290
rect 44526 3238 44528 3290
rect 44282 3236 44288 3238
rect 44344 3236 44368 3238
rect 44424 3236 44448 3238
rect 44504 3236 44528 3238
rect 44584 3236 44590 3238
rect 44282 3227 44590 3236
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44282 2204 44590 2213
rect 44282 2202 44288 2204
rect 44344 2202 44368 2204
rect 44424 2202 44448 2204
rect 44504 2202 44528 2204
rect 44584 2202 44590 2204
rect 44344 2150 44346 2202
rect 44526 2150 44528 2202
rect 44282 2148 44288 2150
rect 44344 2148 44368 2150
rect 44424 2148 44448 2150
rect 44504 2148 44528 2150
rect 44584 2148 44590 2150
rect 44282 2139 44590 2148
rect 44652 1850 44680 3470
rect 44744 2582 44772 3862
rect 44836 3738 44864 4218
rect 45112 4214 45140 4422
rect 45100 4208 45152 4214
rect 45100 4150 45152 4156
rect 45296 4146 45324 4558
rect 45480 4486 45508 5646
rect 45560 5568 45612 5574
rect 45560 5510 45612 5516
rect 45572 5370 45600 5510
rect 45560 5364 45612 5370
rect 45560 5306 45612 5312
rect 45940 5234 45968 6258
rect 46308 5846 46336 6666
rect 46296 5840 46348 5846
rect 46296 5782 46348 5788
rect 46112 5704 46164 5710
rect 46112 5646 46164 5652
rect 46204 5704 46256 5710
rect 46204 5646 46256 5652
rect 46124 5370 46152 5646
rect 46112 5364 46164 5370
rect 46112 5306 46164 5312
rect 45928 5228 45980 5234
rect 45928 5170 45980 5176
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45468 4480 45520 4486
rect 45468 4422 45520 4428
rect 45480 4214 45508 4422
rect 45664 4282 45692 5102
rect 45744 4752 45796 4758
rect 45744 4694 45796 4700
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 45468 4208 45520 4214
rect 45468 4150 45520 4156
rect 45756 4146 45784 4694
rect 45940 4690 45968 5170
rect 45928 4684 45980 4690
rect 45928 4626 45980 4632
rect 45284 4140 45336 4146
rect 45284 4082 45336 4088
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45008 4072 45060 4078
rect 45008 4014 45060 4020
rect 44824 3732 44876 3738
rect 44824 3674 44876 3680
rect 44836 3058 44864 3674
rect 45020 3398 45048 4014
rect 45836 3936 45888 3942
rect 45836 3878 45888 3884
rect 45848 3534 45876 3878
rect 45940 3738 45968 4626
rect 46216 4622 46244 5646
rect 46296 5568 46348 5574
rect 46296 5510 46348 5516
rect 46308 5166 46336 5510
rect 46296 5160 46348 5166
rect 46296 5102 46348 5108
rect 46204 4616 46256 4622
rect 46204 4558 46256 4564
rect 45928 3732 45980 3738
rect 45928 3674 45980 3680
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 46216 3466 46244 4558
rect 46296 4208 46348 4214
rect 46296 4150 46348 4156
rect 46204 3460 46256 3466
rect 46204 3402 46256 3408
rect 45008 3392 45060 3398
rect 45008 3334 45060 3340
rect 46216 3194 46244 3402
rect 46204 3188 46256 3194
rect 46204 3130 46256 3136
rect 44824 3052 44876 3058
rect 44824 2994 44876 3000
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 44822 2816 44878 2825
rect 44822 2751 44878 2760
rect 44732 2576 44784 2582
rect 44732 2518 44784 2524
rect 44836 2446 44864 2751
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 44560 1822 44680 1850
rect 44560 800 44588 1822
rect 45112 800 45140 2926
rect 46308 2854 46336 4150
rect 46400 4049 46428 6666
rect 46480 5228 46532 5234
rect 46480 5170 46532 5176
rect 46492 4758 46520 5170
rect 46480 4752 46532 4758
rect 46480 4694 46532 4700
rect 46386 4040 46442 4049
rect 46386 3975 46442 3984
rect 46492 3942 46520 4694
rect 46664 4480 46716 4486
rect 46664 4422 46716 4428
rect 46676 4214 46704 4422
rect 46664 4208 46716 4214
rect 46664 4150 46716 4156
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46572 3392 46624 3398
rect 46572 3334 46624 3340
rect 46584 2990 46612 3334
rect 46676 3126 46704 4150
rect 46768 3126 46796 7160
rect 46848 6792 46900 6798
rect 46848 6734 46900 6740
rect 46860 6322 46888 6734
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46848 5024 46900 5030
rect 46848 4966 46900 4972
rect 46860 4622 46888 4966
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46952 3670 46980 11698
rect 47044 9042 47072 14010
rect 47136 12434 47164 15846
rect 47584 15564 47636 15570
rect 47584 15506 47636 15512
rect 47308 14272 47360 14278
rect 47308 14214 47360 14220
rect 47320 14006 47348 14214
rect 47308 14000 47360 14006
rect 47308 13942 47360 13948
rect 47216 13320 47268 13326
rect 47216 13262 47268 13268
rect 47228 12986 47256 13262
rect 47216 12980 47268 12986
rect 47216 12922 47268 12928
rect 47136 12406 47256 12434
rect 47228 12238 47256 12406
rect 47320 12306 47348 13942
rect 47400 13184 47452 13190
rect 47400 13126 47452 13132
rect 47412 12986 47440 13126
rect 47400 12980 47452 12986
rect 47400 12922 47452 12928
rect 47308 12300 47360 12306
rect 47308 12242 47360 12248
rect 47216 12232 47268 12238
rect 47216 12174 47268 12180
rect 47308 11552 47360 11558
rect 47308 11494 47360 11500
rect 47320 11150 47348 11494
rect 47283 11144 47348 11150
rect 47335 11104 47348 11144
rect 47400 11144 47452 11150
rect 47283 11086 47335 11092
rect 47400 11086 47452 11092
rect 47124 11008 47176 11014
rect 47124 10950 47176 10956
rect 47032 9036 47084 9042
rect 47032 8978 47084 8984
rect 47032 7880 47084 7886
rect 47032 7822 47084 7828
rect 47044 7478 47072 7822
rect 47032 7472 47084 7478
rect 47032 7414 47084 7420
rect 47032 6656 47084 6662
rect 47032 6598 47084 6604
rect 47044 5370 47072 6598
rect 47032 5364 47084 5370
rect 47032 5306 47084 5312
rect 47136 5250 47164 10950
rect 47412 10742 47440 11086
rect 47400 10736 47452 10742
rect 47400 10678 47452 10684
rect 47412 10266 47440 10678
rect 47400 10260 47452 10266
rect 47400 10202 47452 10208
rect 47596 9738 47624 15506
rect 47688 15026 47716 16730
rect 47780 16250 47808 17682
rect 47872 17270 47900 18022
rect 48424 17882 48452 18158
rect 48412 17876 48464 17882
rect 48412 17818 48464 17824
rect 48688 17808 48740 17814
rect 48688 17750 48740 17756
rect 48320 17536 48372 17542
rect 48320 17478 48372 17484
rect 47860 17264 47912 17270
rect 47860 17206 47912 17212
rect 48136 16584 48188 16590
rect 48136 16526 48188 16532
rect 47768 16244 47820 16250
rect 47768 16186 47820 16192
rect 48148 15638 48176 16526
rect 48332 15722 48360 17478
rect 48596 17264 48648 17270
rect 48596 17206 48648 17212
rect 48608 15910 48636 17206
rect 48700 16658 48728 17750
rect 48792 17338 48820 18158
rect 49332 18080 49384 18086
rect 49332 18022 49384 18028
rect 49240 17740 49292 17746
rect 49240 17682 49292 17688
rect 48964 17672 49016 17678
rect 49148 17672 49200 17678
rect 49016 17632 49148 17660
rect 48964 17614 49016 17620
rect 49148 17614 49200 17620
rect 48780 17332 48832 17338
rect 48780 17274 48832 17280
rect 49252 17270 49280 17682
rect 49344 17610 49372 18022
rect 49332 17604 49384 17610
rect 49332 17546 49384 17552
rect 49240 17264 49292 17270
rect 49240 17206 49292 17212
rect 49344 17134 49372 17546
rect 49332 17128 49384 17134
rect 49332 17070 49384 17076
rect 48780 16992 48832 16998
rect 48780 16934 48832 16940
rect 48792 16794 48820 16934
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 48688 16652 48740 16658
rect 48688 16594 48740 16600
rect 48688 16448 48740 16454
rect 48688 16390 48740 16396
rect 48700 16250 48728 16390
rect 48688 16244 48740 16250
rect 48688 16186 48740 16192
rect 48596 15904 48648 15910
rect 48596 15846 48648 15852
rect 48240 15694 48452 15722
rect 48136 15632 48188 15638
rect 48136 15574 48188 15580
rect 48044 15564 48096 15570
rect 48044 15506 48096 15512
rect 47676 15020 47728 15026
rect 47676 14962 47728 14968
rect 47768 12640 47820 12646
rect 47768 12582 47820 12588
rect 47676 11280 47728 11286
rect 47676 11222 47728 11228
rect 47228 9710 47624 9738
rect 47228 9382 47256 9710
rect 47216 9376 47268 9382
rect 47216 9318 47268 9324
rect 47228 8906 47256 9318
rect 47216 8900 47268 8906
rect 47216 8842 47268 8848
rect 47688 8566 47716 11222
rect 47780 11218 47808 12582
rect 47768 11212 47820 11218
rect 47768 11154 47820 11160
rect 47780 10810 47808 11154
rect 47768 10804 47820 10810
rect 47768 10746 47820 10752
rect 47952 10600 48004 10606
rect 47952 10542 48004 10548
rect 47964 10266 47992 10542
rect 48056 10470 48084 15506
rect 48240 15502 48268 15694
rect 48228 15496 48280 15502
rect 48228 15438 48280 15444
rect 48424 15026 48452 15694
rect 48608 15366 48636 15846
rect 48596 15360 48648 15366
rect 48596 15302 48648 15308
rect 48688 15360 48740 15366
rect 48688 15302 48740 15308
rect 48700 15094 48728 15302
rect 48688 15088 48740 15094
rect 48688 15030 48740 15036
rect 48412 15020 48464 15026
rect 48412 14962 48464 14968
rect 49332 15020 49384 15026
rect 49332 14962 49384 14968
rect 49344 14482 49372 14962
rect 49332 14476 49384 14482
rect 49332 14418 49384 14424
rect 48320 14340 48372 14346
rect 48320 14282 48372 14288
rect 48332 14074 48360 14282
rect 48780 14272 48832 14278
rect 48780 14214 48832 14220
rect 48872 14272 48924 14278
rect 48872 14214 48924 14220
rect 48320 14068 48372 14074
rect 48320 14010 48372 14016
rect 48792 13394 48820 14214
rect 48884 13938 48912 14214
rect 48872 13932 48924 13938
rect 48872 13874 48924 13880
rect 48136 13388 48188 13394
rect 48136 13330 48188 13336
rect 48780 13388 48832 13394
rect 48780 13330 48832 13336
rect 48148 11354 48176 13330
rect 48320 12776 48372 12782
rect 48320 12718 48372 12724
rect 48332 11898 48360 12718
rect 49056 12164 49108 12170
rect 49056 12106 49108 12112
rect 48596 12096 48648 12102
rect 48596 12038 48648 12044
rect 48780 12096 48832 12102
rect 48780 12038 48832 12044
rect 48320 11892 48372 11898
rect 48320 11834 48372 11840
rect 48320 11552 48372 11558
rect 48320 11494 48372 11500
rect 48136 11348 48188 11354
rect 48136 11290 48188 11296
rect 48148 10742 48176 11290
rect 48228 11280 48280 11286
rect 48228 11222 48280 11228
rect 48136 10736 48188 10742
rect 48136 10678 48188 10684
rect 48044 10464 48096 10470
rect 48044 10406 48096 10412
rect 48056 10266 48084 10406
rect 47952 10260 48004 10266
rect 47952 10202 48004 10208
rect 48044 10260 48096 10266
rect 48044 10202 48096 10208
rect 47860 9920 47912 9926
rect 47860 9862 47912 9868
rect 47872 9042 47900 9862
rect 47964 9518 47992 10202
rect 48148 9994 48176 10678
rect 48240 10674 48268 11222
rect 48228 10668 48280 10674
rect 48228 10610 48280 10616
rect 48136 9988 48188 9994
rect 48136 9930 48188 9936
rect 47952 9512 48004 9518
rect 47952 9454 48004 9460
rect 48136 9512 48188 9518
rect 48136 9454 48188 9460
rect 48044 9376 48096 9382
rect 48044 9318 48096 9324
rect 48056 9110 48084 9318
rect 48044 9104 48096 9110
rect 48044 9046 48096 9052
rect 47860 9036 47912 9042
rect 47860 8978 47912 8984
rect 47768 8832 47820 8838
rect 47768 8774 47820 8780
rect 47676 8560 47728 8566
rect 47676 8502 47728 8508
rect 47688 8022 47716 8502
rect 47676 8016 47728 8022
rect 47676 7958 47728 7964
rect 47780 7954 47808 8774
rect 47768 7948 47820 7954
rect 47768 7890 47820 7896
rect 47872 7546 47900 8978
rect 48148 8634 48176 9454
rect 48228 9376 48280 9382
rect 48228 9318 48280 9324
rect 48240 8838 48268 9318
rect 48228 8832 48280 8838
rect 48228 8774 48280 8780
rect 48136 8628 48188 8634
rect 48136 8570 48188 8576
rect 47952 7880 48004 7886
rect 47952 7822 48004 7828
rect 47216 7540 47268 7546
rect 47216 7482 47268 7488
rect 47860 7540 47912 7546
rect 47860 7482 47912 7488
rect 47044 5222 47164 5250
rect 47044 4282 47072 5222
rect 47124 4480 47176 4486
rect 47124 4422 47176 4428
rect 47032 4276 47084 4282
rect 47032 4218 47084 4224
rect 47136 4078 47164 4422
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 46940 3664 46992 3670
rect 47228 3618 47256 7482
rect 47308 6996 47360 7002
rect 47308 6938 47360 6944
rect 47320 6322 47348 6938
rect 47872 6934 47900 7482
rect 47860 6928 47912 6934
rect 47860 6870 47912 6876
rect 47400 6724 47452 6730
rect 47400 6666 47452 6672
rect 47412 6458 47440 6666
rect 47964 6662 47992 7822
rect 48044 7744 48096 7750
rect 48044 7686 48096 7692
rect 48056 6866 48084 7686
rect 48044 6860 48096 6866
rect 48044 6802 48096 6808
rect 47952 6656 48004 6662
rect 47952 6598 48004 6604
rect 47400 6452 47452 6458
rect 47400 6394 47452 6400
rect 47308 6316 47360 6322
rect 47964 6304 47992 6598
rect 48044 6316 48096 6322
rect 47964 6276 48044 6304
rect 47308 6258 47360 6264
rect 48044 6258 48096 6264
rect 47400 6248 47452 6254
rect 47400 6190 47452 6196
rect 47412 5914 47440 6190
rect 47400 5908 47452 5914
rect 47400 5850 47452 5856
rect 47860 5160 47912 5166
rect 47860 5102 47912 5108
rect 47768 4616 47820 4622
rect 47768 4558 47820 4564
rect 47780 4282 47808 4558
rect 47872 4486 47900 5102
rect 47860 4480 47912 4486
rect 47860 4422 47912 4428
rect 47952 4480 48004 4486
rect 47952 4422 48004 4428
rect 47768 4276 47820 4282
rect 47768 4218 47820 4224
rect 47492 4072 47544 4078
rect 47492 4014 47544 4020
rect 46940 3606 46992 3612
rect 47044 3590 47256 3618
rect 47044 3482 47072 3590
rect 46952 3454 47072 3482
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 47214 3496 47270 3505
rect 46952 3194 46980 3454
rect 47136 3194 47164 3470
rect 47270 3454 47348 3482
rect 47504 3466 47532 4014
rect 47780 3942 47808 4218
rect 47964 4146 47992 4422
rect 47952 4140 48004 4146
rect 47952 4082 48004 4088
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47214 3431 47270 3440
rect 46940 3188 46992 3194
rect 46940 3130 46992 3136
rect 47124 3188 47176 3194
rect 47124 3130 47176 3136
rect 46664 3120 46716 3126
rect 46664 3062 46716 3068
rect 46756 3120 46808 3126
rect 46756 3062 46808 3068
rect 46848 3120 46900 3126
rect 46848 3062 46900 3068
rect 46572 2984 46624 2990
rect 46676 2972 46704 3062
rect 46756 2984 46808 2990
rect 46676 2944 46756 2972
rect 46572 2926 46624 2932
rect 46756 2926 46808 2932
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 46296 2848 46348 2854
rect 46296 2790 46348 2796
rect 45572 2514 45600 2790
rect 45560 2508 45612 2514
rect 45560 2450 45612 2456
rect 46584 2446 46612 2926
rect 46860 2836 46888 3062
rect 46940 2916 46992 2922
rect 46940 2858 46992 2864
rect 46676 2808 46888 2836
rect 46572 2440 46624 2446
rect 46572 2382 46624 2388
rect 45652 2372 45704 2378
rect 45652 2314 45704 2320
rect 45664 800 45692 2314
rect 46216 870 46336 898
rect 46216 800 46244 870
rect 42996 734 43208 762
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46308 762 46336 870
rect 46676 762 46704 2808
rect 46952 2802 46980 2858
rect 46927 2774 46980 2802
rect 47320 2774 47348 3454
rect 47492 3460 47544 3466
rect 47492 3402 47544 3408
rect 46768 2746 46955 2774
rect 47228 2746 47348 2774
rect 46768 800 46796 2746
rect 47228 2650 47256 2746
rect 47216 2644 47268 2650
rect 47216 2586 47268 2592
rect 47676 2508 47728 2514
rect 47676 2450 47728 2456
rect 47320 870 47440 898
rect 47320 800 47348 870
rect 46308 734 46704 762
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47412 762 47440 870
rect 47688 762 47716 2450
rect 47964 2446 47992 4082
rect 48044 3936 48096 3942
rect 48044 3878 48096 3884
rect 48056 3534 48084 3878
rect 48044 3528 48096 3534
rect 48044 3470 48096 3476
rect 48332 3126 48360 11494
rect 48608 11218 48636 12038
rect 48792 11354 48820 12038
rect 49068 11898 49096 12106
rect 49056 11892 49108 11898
rect 49056 11834 49108 11840
rect 48872 11756 48924 11762
rect 48872 11698 48924 11704
rect 48884 11354 48912 11698
rect 49436 11558 49464 20470
rect 49792 19712 49844 19718
rect 49792 19654 49844 19660
rect 49700 19508 49752 19514
rect 49700 19450 49752 19456
rect 49516 17536 49568 17542
rect 49516 17478 49568 17484
rect 49528 17270 49556 17478
rect 49516 17264 49568 17270
rect 49516 17206 49568 17212
rect 49528 16046 49556 17206
rect 49712 16114 49740 19450
rect 49700 16108 49752 16114
rect 49700 16050 49752 16056
rect 49516 16040 49568 16046
rect 49516 15982 49568 15988
rect 49608 15428 49660 15434
rect 49608 15370 49660 15376
rect 49620 15162 49648 15370
rect 49608 15156 49660 15162
rect 49608 15098 49660 15104
rect 49620 14890 49648 15098
rect 49608 14884 49660 14890
rect 49608 14826 49660 14832
rect 49516 14816 49568 14822
rect 49516 14758 49568 14764
rect 49528 14482 49556 14758
rect 49516 14476 49568 14482
rect 49516 14418 49568 14424
rect 49700 14476 49752 14482
rect 49700 14418 49752 14424
rect 49528 14074 49556 14418
rect 49516 14068 49568 14074
rect 49516 14010 49568 14016
rect 49528 12209 49556 14010
rect 49712 13530 49740 14418
rect 49700 13524 49752 13530
rect 49700 13466 49752 13472
rect 49514 12200 49570 12209
rect 49514 12135 49570 12144
rect 49608 11688 49660 11694
rect 49608 11630 49660 11636
rect 49424 11552 49476 11558
rect 49424 11494 49476 11500
rect 49620 11354 49648 11630
rect 48780 11348 48832 11354
rect 48780 11290 48832 11296
rect 48872 11348 48924 11354
rect 48872 11290 48924 11296
rect 49608 11348 49660 11354
rect 49608 11290 49660 11296
rect 48596 11212 48648 11218
rect 48596 11154 48648 11160
rect 48410 11112 48466 11121
rect 48410 11047 48466 11056
rect 48424 7886 48452 11047
rect 48608 10742 48636 11154
rect 49700 11144 49752 11150
rect 49700 11086 49752 11092
rect 48688 11008 48740 11014
rect 48688 10950 48740 10956
rect 48700 10810 48728 10950
rect 48688 10804 48740 10810
rect 48688 10746 48740 10752
rect 48596 10736 48648 10742
rect 48596 10678 48648 10684
rect 48700 9042 48728 10746
rect 49712 10606 49740 11086
rect 49804 10810 49832 19654
rect 50080 17184 50108 21830
rect 50172 20534 50200 21966
rect 50252 21480 50304 21486
rect 50252 21422 50304 21428
rect 50264 21146 50292 21422
rect 50252 21140 50304 21146
rect 50252 21082 50304 21088
rect 50160 20528 50212 20534
rect 50160 20470 50212 20476
rect 50172 19922 50200 20470
rect 50160 19916 50212 19922
rect 50160 19858 50212 19864
rect 50172 19378 50200 19858
rect 50252 19780 50304 19786
rect 50252 19722 50304 19728
rect 50264 19514 50292 19722
rect 50252 19508 50304 19514
rect 50252 19450 50304 19456
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 50172 18290 50200 19314
rect 50160 18284 50212 18290
rect 50160 18226 50212 18232
rect 50160 17808 50212 17814
rect 50160 17750 50212 17756
rect 50172 17320 50200 17750
rect 50252 17536 50304 17542
rect 50632 17490 50660 22714
rect 50816 21486 50844 23666
rect 51184 22574 51212 24890
rect 51276 24614 51304 25774
rect 51504 25596 51812 25605
rect 51504 25594 51510 25596
rect 51566 25594 51590 25596
rect 51646 25594 51670 25596
rect 51726 25594 51750 25596
rect 51806 25594 51812 25596
rect 51566 25542 51568 25594
rect 51748 25542 51750 25594
rect 51504 25540 51510 25542
rect 51566 25540 51590 25542
rect 51646 25540 51670 25542
rect 51726 25540 51750 25542
rect 51806 25540 51812 25542
rect 51504 25531 51812 25540
rect 52012 25294 52040 25774
rect 52104 25362 52132 26726
rect 52368 26240 52420 26246
rect 52368 26182 52420 26188
rect 52276 25900 52328 25906
rect 52276 25842 52328 25848
rect 52288 25362 52316 25842
rect 52380 25770 52408 26182
rect 53852 25974 53880 26726
rect 54208 26376 54260 26382
rect 54208 26318 54260 26324
rect 54392 26376 54444 26382
rect 54392 26318 54444 26324
rect 53840 25968 53892 25974
rect 53840 25910 53892 25916
rect 52368 25764 52420 25770
rect 52368 25706 52420 25712
rect 54220 25498 54248 26318
rect 54404 25974 54432 26318
rect 54496 26042 54524 26880
rect 54668 26862 54720 26868
rect 54668 26512 54720 26518
rect 54668 26454 54720 26460
rect 54576 26240 54628 26246
rect 54576 26182 54628 26188
rect 54484 26036 54536 26042
rect 54484 25978 54536 25984
rect 54392 25968 54444 25974
rect 54392 25910 54444 25916
rect 54588 25906 54616 26182
rect 54576 25900 54628 25906
rect 54576 25842 54628 25848
rect 54208 25492 54260 25498
rect 54208 25434 54260 25440
rect 54588 25430 54616 25842
rect 54576 25424 54628 25430
rect 54576 25366 54628 25372
rect 54680 25362 54708 26454
rect 58726 26140 59034 26149
rect 58726 26138 58732 26140
rect 58788 26138 58812 26140
rect 58868 26138 58892 26140
rect 58948 26138 58972 26140
rect 59028 26138 59034 26140
rect 58788 26086 58790 26138
rect 58970 26086 58972 26138
rect 58726 26084 58732 26086
rect 58788 26084 58812 26086
rect 58868 26084 58892 26086
rect 58948 26084 58972 26086
rect 59028 26084 59034 26086
rect 58726 26075 59034 26084
rect 52092 25356 52144 25362
rect 52092 25298 52144 25304
rect 52276 25356 52328 25362
rect 52276 25298 52328 25304
rect 52552 25356 52604 25362
rect 52552 25298 52604 25304
rect 53380 25356 53432 25362
rect 53380 25298 53432 25304
rect 54668 25356 54720 25362
rect 54668 25298 54720 25304
rect 52000 25288 52052 25294
rect 52000 25230 52052 25236
rect 52012 24954 52040 25230
rect 52564 24954 52592 25298
rect 53196 25152 53248 25158
rect 53196 25094 53248 25100
rect 52000 24948 52052 24954
rect 52000 24890 52052 24896
rect 52552 24948 52604 24954
rect 52552 24890 52604 24896
rect 52552 24812 52604 24818
rect 52552 24754 52604 24760
rect 51264 24608 51316 24614
rect 51264 24550 51316 24556
rect 51276 23118 51304 24550
rect 51504 24508 51812 24517
rect 51504 24506 51510 24508
rect 51566 24506 51590 24508
rect 51646 24506 51670 24508
rect 51726 24506 51750 24508
rect 51806 24506 51812 24508
rect 51566 24454 51568 24506
rect 51748 24454 51750 24506
rect 51504 24452 51510 24454
rect 51566 24452 51590 24454
rect 51646 24452 51670 24454
rect 51726 24452 51750 24454
rect 51806 24452 51812 24454
rect 51504 24443 51812 24452
rect 51908 24200 51960 24206
rect 51908 24142 51960 24148
rect 51356 24064 51408 24070
rect 51356 24006 51408 24012
rect 51368 23662 51396 24006
rect 51356 23656 51408 23662
rect 51356 23598 51408 23604
rect 51368 23304 51396 23598
rect 51504 23420 51812 23429
rect 51504 23418 51510 23420
rect 51566 23418 51590 23420
rect 51646 23418 51670 23420
rect 51726 23418 51750 23420
rect 51806 23418 51812 23420
rect 51566 23366 51568 23418
rect 51748 23366 51750 23418
rect 51504 23364 51510 23366
rect 51566 23364 51590 23366
rect 51646 23364 51670 23366
rect 51726 23364 51750 23366
rect 51806 23364 51812 23366
rect 51504 23355 51812 23364
rect 51920 23322 51948 24142
rect 52460 24064 52512 24070
rect 52460 24006 52512 24012
rect 52000 23724 52052 23730
rect 52000 23666 52052 23672
rect 51908 23316 51960 23322
rect 51368 23276 51672 23304
rect 51264 23112 51316 23118
rect 51264 23054 51316 23060
rect 51644 22642 51672 23276
rect 51908 23258 51960 23264
rect 51816 22976 51868 22982
rect 51816 22918 51868 22924
rect 51632 22636 51684 22642
rect 51632 22578 51684 22584
rect 51172 22568 51224 22574
rect 51092 22516 51172 22522
rect 51448 22568 51500 22574
rect 51092 22510 51224 22516
rect 51368 22516 51448 22522
rect 51368 22510 51500 22516
rect 51092 22494 51212 22510
rect 51368 22494 51488 22510
rect 51828 22506 51856 22918
rect 52012 22778 52040 23666
rect 52472 23662 52500 24006
rect 52460 23656 52512 23662
rect 52460 23598 52512 23604
rect 52000 22772 52052 22778
rect 52000 22714 52052 22720
rect 52472 22642 52500 23598
rect 52460 22636 52512 22642
rect 52460 22578 52512 22584
rect 52368 22568 52420 22574
rect 52368 22510 52420 22516
rect 51816 22500 51868 22506
rect 50988 21956 51040 21962
rect 50988 21898 51040 21904
rect 51000 21690 51028 21898
rect 51092 21894 51120 22494
rect 51172 22432 51224 22438
rect 51172 22374 51224 22380
rect 51080 21888 51132 21894
rect 51080 21830 51132 21836
rect 51184 21690 51212 22374
rect 51368 22098 51396 22494
rect 51816 22442 51868 22448
rect 51504 22332 51812 22341
rect 51504 22330 51510 22332
rect 51566 22330 51590 22332
rect 51646 22330 51670 22332
rect 51726 22330 51750 22332
rect 51806 22330 51812 22332
rect 51566 22278 51568 22330
rect 51748 22278 51750 22330
rect 51504 22276 51510 22278
rect 51566 22276 51590 22278
rect 51646 22276 51670 22278
rect 51726 22276 51750 22278
rect 51806 22276 51812 22278
rect 51504 22267 51812 22276
rect 51356 22092 51408 22098
rect 51356 22034 51408 22040
rect 50988 21684 51040 21690
rect 50988 21626 51040 21632
rect 51172 21684 51224 21690
rect 51172 21626 51224 21632
rect 51368 21622 51396 22034
rect 51356 21616 51408 21622
rect 51356 21558 51408 21564
rect 50804 21480 50856 21486
rect 50804 21422 50856 21428
rect 51264 21480 51316 21486
rect 51264 21422 51316 21428
rect 51276 19718 51304 21422
rect 51356 21344 51408 21350
rect 51356 21286 51408 21292
rect 51264 19712 51316 19718
rect 51264 19654 51316 19660
rect 51368 19514 51396 21286
rect 51504 21244 51812 21253
rect 51504 21242 51510 21244
rect 51566 21242 51590 21244
rect 51646 21242 51670 21244
rect 51726 21242 51750 21244
rect 51806 21242 51812 21244
rect 51566 21190 51568 21242
rect 51748 21190 51750 21242
rect 51504 21188 51510 21190
rect 51566 21188 51590 21190
rect 51646 21188 51670 21190
rect 51726 21188 51750 21190
rect 51806 21188 51812 21190
rect 51504 21179 51812 21188
rect 52380 21146 52408 22510
rect 52092 21140 52144 21146
rect 52092 21082 52144 21088
rect 52368 21140 52420 21146
rect 52368 21082 52420 21088
rect 51504 20156 51812 20165
rect 51504 20154 51510 20156
rect 51566 20154 51590 20156
rect 51646 20154 51670 20156
rect 51726 20154 51750 20156
rect 51806 20154 51812 20156
rect 51566 20102 51568 20154
rect 51748 20102 51750 20154
rect 51504 20100 51510 20102
rect 51566 20100 51590 20102
rect 51646 20100 51670 20102
rect 51726 20100 51750 20102
rect 51806 20100 51812 20102
rect 51504 20091 51812 20100
rect 52000 19984 52052 19990
rect 52000 19926 52052 19932
rect 51816 19916 51868 19922
rect 51816 19858 51868 19864
rect 51828 19514 51856 19858
rect 51356 19508 51408 19514
rect 51356 19450 51408 19456
rect 51816 19508 51868 19514
rect 51816 19450 51868 19456
rect 51264 19440 51316 19446
rect 51264 19382 51316 19388
rect 50988 19372 51040 19378
rect 50988 19314 51040 19320
rect 50304 17484 50660 17490
rect 50252 17478 50660 17484
rect 50264 17462 50660 17478
rect 50172 17292 50384 17320
rect 50160 17196 50212 17202
rect 50080 17156 50160 17184
rect 50080 16726 50108 17156
rect 50160 17138 50212 17144
rect 50356 17184 50384 17292
rect 50436 17196 50488 17202
rect 50356 17156 50436 17184
rect 50252 16992 50304 16998
rect 50252 16934 50304 16940
rect 50068 16720 50120 16726
rect 50068 16662 50120 16668
rect 50264 15502 50292 16934
rect 50356 16250 50384 17156
rect 50436 17138 50488 17144
rect 50632 17134 50660 17462
rect 50620 17128 50672 17134
rect 50620 17070 50672 17076
rect 50712 16652 50764 16658
rect 50712 16594 50764 16600
rect 50344 16244 50396 16250
rect 50344 16186 50396 16192
rect 50620 16040 50672 16046
rect 50620 15982 50672 15988
rect 50344 15904 50396 15910
rect 50344 15846 50396 15852
rect 50436 15904 50488 15910
rect 50436 15846 50488 15852
rect 50252 15496 50304 15502
rect 50252 15438 50304 15444
rect 50068 15428 50120 15434
rect 50068 15370 50120 15376
rect 49884 15360 49936 15366
rect 49884 15302 49936 15308
rect 49896 14414 49924 15302
rect 50080 14958 50108 15370
rect 50068 14952 50120 14958
rect 50068 14894 50120 14900
rect 49884 14408 49936 14414
rect 49884 14350 49936 14356
rect 49976 14272 50028 14278
rect 49976 14214 50028 14220
rect 49988 14006 50016 14214
rect 49976 14000 50028 14006
rect 49976 13942 50028 13948
rect 49988 12986 50016 13942
rect 49976 12980 50028 12986
rect 49976 12922 50028 12928
rect 49988 11762 50016 12922
rect 50080 12714 50108 14894
rect 50068 12708 50120 12714
rect 50068 12650 50120 12656
rect 49976 11756 50028 11762
rect 50356 11744 50384 15846
rect 50448 14006 50476 15846
rect 50632 15162 50660 15982
rect 50724 15162 50752 16594
rect 50620 15156 50672 15162
rect 50620 15098 50672 15104
rect 50712 15156 50764 15162
rect 50712 15098 50764 15104
rect 50896 14952 50948 14958
rect 50896 14894 50948 14900
rect 50804 14408 50856 14414
rect 50804 14350 50856 14356
rect 50436 14000 50488 14006
rect 50436 13942 50488 13948
rect 50436 13728 50488 13734
rect 50436 13670 50488 13676
rect 50448 13190 50476 13670
rect 50816 13326 50844 14350
rect 50908 14074 50936 14894
rect 50896 14068 50948 14074
rect 50896 14010 50948 14016
rect 50804 13320 50856 13326
rect 50804 13262 50856 13268
rect 50436 13184 50488 13190
rect 50436 13126 50488 13132
rect 50448 11914 50476 13126
rect 50528 12844 50580 12850
rect 50528 12786 50580 12792
rect 50540 12442 50568 12786
rect 50528 12436 50580 12442
rect 50528 12378 50580 12384
rect 50448 11886 50568 11914
rect 50436 11756 50488 11762
rect 50356 11716 50436 11744
rect 49976 11698 50028 11704
rect 50436 11698 50488 11704
rect 50540 11354 50568 11886
rect 51000 11558 51028 19314
rect 51172 18624 51224 18630
rect 51172 18566 51224 18572
rect 51184 17202 51212 18566
rect 51172 17196 51224 17202
rect 51172 17138 51224 17144
rect 51276 16250 51304 19382
rect 51504 19068 51812 19077
rect 51504 19066 51510 19068
rect 51566 19066 51590 19068
rect 51646 19066 51670 19068
rect 51726 19066 51750 19068
rect 51806 19066 51812 19068
rect 51566 19014 51568 19066
rect 51748 19014 51750 19066
rect 51504 19012 51510 19014
rect 51566 19012 51590 19014
rect 51646 19012 51670 19014
rect 51726 19012 51750 19014
rect 51806 19012 51812 19014
rect 51504 19003 51812 19012
rect 51816 18760 51868 18766
rect 51816 18702 51868 18708
rect 51828 18426 51856 18702
rect 51908 18624 51960 18630
rect 51908 18566 51960 18572
rect 51920 18426 51948 18566
rect 51816 18420 51868 18426
rect 51816 18362 51868 18368
rect 51908 18420 51960 18426
rect 51908 18362 51960 18368
rect 51908 18080 51960 18086
rect 51908 18022 51960 18028
rect 51504 17980 51812 17989
rect 51504 17978 51510 17980
rect 51566 17978 51590 17980
rect 51646 17978 51670 17980
rect 51726 17978 51750 17980
rect 51806 17978 51812 17980
rect 51566 17926 51568 17978
rect 51748 17926 51750 17978
rect 51504 17924 51510 17926
rect 51566 17924 51590 17926
rect 51646 17924 51670 17926
rect 51726 17924 51750 17926
rect 51806 17924 51812 17926
rect 51504 17915 51812 17924
rect 51920 17678 51948 18022
rect 51908 17672 51960 17678
rect 51908 17614 51960 17620
rect 51908 17536 51960 17542
rect 51908 17478 51960 17484
rect 51920 17134 51948 17478
rect 51908 17128 51960 17134
rect 51908 17070 51960 17076
rect 51356 17060 51408 17066
rect 51356 17002 51408 17008
rect 51368 16794 51396 17002
rect 51504 16892 51812 16901
rect 51504 16890 51510 16892
rect 51566 16890 51590 16892
rect 51646 16890 51670 16892
rect 51726 16890 51750 16892
rect 51806 16890 51812 16892
rect 51566 16838 51568 16890
rect 51748 16838 51750 16890
rect 51504 16836 51510 16838
rect 51566 16836 51590 16838
rect 51646 16836 51670 16838
rect 51726 16836 51750 16838
rect 51806 16836 51812 16838
rect 51504 16827 51812 16836
rect 51356 16788 51408 16794
rect 51356 16730 51408 16736
rect 51264 16244 51316 16250
rect 51264 16186 51316 16192
rect 51276 15570 51304 16186
rect 52012 16114 52040 19926
rect 52104 19854 52132 21082
rect 52184 20936 52236 20942
rect 52184 20878 52236 20884
rect 52196 20602 52224 20878
rect 52184 20596 52236 20602
rect 52184 20538 52236 20544
rect 52368 20256 52420 20262
rect 52368 20198 52420 20204
rect 52380 20058 52408 20198
rect 52368 20052 52420 20058
rect 52368 19994 52420 20000
rect 52092 19848 52144 19854
rect 52092 19790 52144 19796
rect 52276 19712 52328 19718
rect 52276 19654 52328 19660
rect 52092 17536 52144 17542
rect 52092 17478 52144 17484
rect 52104 17338 52132 17478
rect 52092 17332 52144 17338
rect 52092 17274 52144 17280
rect 52184 17128 52236 17134
rect 52184 17070 52236 17076
rect 52092 16448 52144 16454
rect 52092 16390 52144 16396
rect 52000 16108 52052 16114
rect 52000 16050 52052 16056
rect 51356 15904 51408 15910
rect 51356 15846 51408 15852
rect 51264 15564 51316 15570
rect 51264 15506 51316 15512
rect 51264 15360 51316 15366
rect 51264 15302 51316 15308
rect 51080 14884 51132 14890
rect 51080 14826 51132 14832
rect 51092 14482 51120 14826
rect 51276 14618 51304 15302
rect 51264 14612 51316 14618
rect 51264 14554 51316 14560
rect 51080 14476 51132 14482
rect 51080 14418 51132 14424
rect 51264 14476 51316 14482
rect 51264 14418 51316 14424
rect 51080 13864 51132 13870
rect 51080 13806 51132 13812
rect 51092 12238 51120 13806
rect 51276 13734 51304 14418
rect 51264 13728 51316 13734
rect 51264 13670 51316 13676
rect 51368 12434 51396 15846
rect 51504 15804 51812 15813
rect 51504 15802 51510 15804
rect 51566 15802 51590 15804
rect 51646 15802 51670 15804
rect 51726 15802 51750 15804
rect 51806 15802 51812 15804
rect 51566 15750 51568 15802
rect 51748 15750 51750 15802
rect 51504 15748 51510 15750
rect 51566 15748 51590 15750
rect 51646 15748 51670 15750
rect 51726 15748 51750 15750
rect 51806 15748 51812 15750
rect 51504 15739 51812 15748
rect 51908 15564 51960 15570
rect 51908 15506 51960 15512
rect 51816 15360 51868 15366
rect 51816 15302 51868 15308
rect 51828 14906 51856 15302
rect 51920 15042 51948 15506
rect 52104 15502 52132 16390
rect 52092 15496 52144 15502
rect 52092 15438 52144 15444
rect 51920 15014 52040 15042
rect 51828 14878 51948 14906
rect 51504 14716 51812 14725
rect 51504 14714 51510 14716
rect 51566 14714 51590 14716
rect 51646 14714 51670 14716
rect 51726 14714 51750 14716
rect 51806 14714 51812 14716
rect 51566 14662 51568 14714
rect 51748 14662 51750 14714
rect 51504 14660 51510 14662
rect 51566 14660 51590 14662
rect 51646 14660 51670 14662
rect 51726 14660 51750 14662
rect 51806 14660 51812 14662
rect 51504 14651 51812 14660
rect 51920 13938 51948 14878
rect 52012 14498 52040 15014
rect 52104 14890 52132 15438
rect 52196 15366 52224 17070
rect 52184 15360 52236 15366
rect 52184 15302 52236 15308
rect 52196 15162 52224 15302
rect 52184 15156 52236 15162
rect 52184 15098 52236 15104
rect 52092 14884 52144 14890
rect 52092 14826 52144 14832
rect 52012 14470 52132 14498
rect 52000 14408 52052 14414
rect 52000 14350 52052 14356
rect 52012 14074 52040 14350
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 51908 13932 51960 13938
rect 51908 13874 51960 13880
rect 52000 13864 52052 13870
rect 52000 13806 52052 13812
rect 51504 13628 51812 13637
rect 51504 13626 51510 13628
rect 51566 13626 51590 13628
rect 51646 13626 51670 13628
rect 51726 13626 51750 13628
rect 51806 13626 51812 13628
rect 51566 13574 51568 13626
rect 51748 13574 51750 13626
rect 51504 13572 51510 13574
rect 51566 13572 51590 13574
rect 51646 13572 51670 13574
rect 51726 13572 51750 13574
rect 51806 13572 51812 13574
rect 51504 13563 51812 13572
rect 51504 12540 51812 12549
rect 51504 12538 51510 12540
rect 51566 12538 51590 12540
rect 51646 12538 51670 12540
rect 51726 12538 51750 12540
rect 51806 12538 51812 12540
rect 51566 12486 51568 12538
rect 51748 12486 51750 12538
rect 51504 12484 51510 12486
rect 51566 12484 51590 12486
rect 51646 12484 51670 12486
rect 51726 12484 51750 12486
rect 51806 12484 51812 12486
rect 51504 12475 51812 12484
rect 52012 12442 52040 13806
rect 51184 12406 51396 12434
rect 52000 12436 52052 12442
rect 51080 12232 51132 12238
rect 51080 12174 51132 12180
rect 51184 11762 51212 12406
rect 52000 12378 52052 12384
rect 52104 12322 52132 14470
rect 52012 12294 52132 12322
rect 51262 12200 51318 12209
rect 51262 12135 51318 12144
rect 51172 11756 51224 11762
rect 51172 11698 51224 11704
rect 50712 11552 50764 11558
rect 50712 11494 50764 11500
rect 50988 11552 51040 11558
rect 50988 11494 51040 11500
rect 50528 11348 50580 11354
rect 50528 11290 50580 11296
rect 49792 10804 49844 10810
rect 49792 10746 49844 10752
rect 50540 10674 50568 11290
rect 49884 10668 49936 10674
rect 50528 10668 50580 10674
rect 49936 10628 50016 10656
rect 49884 10610 49936 10616
rect 49700 10600 49752 10606
rect 49700 10542 49752 10548
rect 49700 10056 49752 10062
rect 49700 9998 49752 10004
rect 49712 9722 49740 9998
rect 49700 9716 49752 9722
rect 49700 9658 49752 9664
rect 48688 9036 48740 9042
rect 48688 8978 48740 8984
rect 49148 8832 49200 8838
rect 49148 8774 49200 8780
rect 49160 8634 49188 8774
rect 49148 8628 49200 8634
rect 49148 8570 49200 8576
rect 49884 8288 49936 8294
rect 49884 8230 49936 8236
rect 49792 8016 49844 8022
rect 49792 7958 49844 7964
rect 48412 7880 48464 7886
rect 48412 7822 48464 7828
rect 48596 7744 48648 7750
rect 48596 7686 48648 7692
rect 48608 7410 48636 7686
rect 48596 7404 48648 7410
rect 48596 7346 48648 7352
rect 49804 7002 49832 7958
rect 49896 7478 49924 8230
rect 49884 7472 49936 7478
rect 49884 7414 49936 7420
rect 49792 6996 49844 7002
rect 49792 6938 49844 6944
rect 48412 6792 48464 6798
rect 48412 6734 48464 6740
rect 48424 6458 48452 6734
rect 48412 6452 48464 6458
rect 48412 6394 48464 6400
rect 49332 6316 49384 6322
rect 49332 6258 49384 6264
rect 49344 5914 49372 6258
rect 49332 5908 49384 5914
rect 49332 5850 49384 5856
rect 49700 5840 49752 5846
rect 49700 5782 49752 5788
rect 49712 5370 49740 5782
rect 49700 5364 49752 5370
rect 49700 5306 49752 5312
rect 49332 5024 49384 5030
rect 49332 4966 49384 4972
rect 49700 5024 49752 5030
rect 49700 4966 49752 4972
rect 49344 4826 49372 4966
rect 49332 4820 49384 4826
rect 49332 4762 49384 4768
rect 49712 4486 49740 4966
rect 49884 4616 49936 4622
rect 49884 4558 49936 4564
rect 48688 4480 48740 4486
rect 48688 4422 48740 4428
rect 49700 4480 49752 4486
rect 49700 4422 49752 4428
rect 48700 4282 48728 4422
rect 49896 4282 49924 4558
rect 48688 4276 48740 4282
rect 48688 4218 48740 4224
rect 49884 4276 49936 4282
rect 49884 4218 49936 4224
rect 48596 3392 48648 3398
rect 48596 3334 48648 3340
rect 48608 3126 48636 3334
rect 48700 3194 48728 4218
rect 49240 4140 49292 4146
rect 49240 4082 49292 4088
rect 49424 4140 49476 4146
rect 49424 4082 49476 4088
rect 48964 4072 49016 4078
rect 48964 4014 49016 4020
rect 48976 3466 49004 4014
rect 49252 3670 49280 4082
rect 49240 3664 49292 3670
rect 49240 3606 49292 3612
rect 49056 3528 49108 3534
rect 49056 3470 49108 3476
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 3194 49004 3402
rect 48688 3188 48740 3194
rect 48688 3130 48740 3136
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48320 3120 48372 3126
rect 48320 3062 48372 3068
rect 48596 3120 48648 3126
rect 48596 3062 48648 3068
rect 49068 3058 49096 3470
rect 49148 3392 49200 3398
rect 49148 3334 49200 3340
rect 49160 3058 49188 3334
rect 49056 3052 49108 3058
rect 49056 2994 49108 3000
rect 49148 3052 49200 3058
rect 49148 2994 49200 3000
rect 48964 2984 49016 2990
rect 48964 2926 49016 2932
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 47860 2372 47912 2378
rect 47860 2314 47912 2320
rect 47872 800 47900 2314
rect 48424 800 48452 2382
rect 48976 800 49004 2926
rect 49436 2922 49464 4082
rect 49792 4072 49844 4078
rect 49792 4014 49844 4020
rect 49424 2916 49476 2922
rect 49424 2858 49476 2864
rect 49804 2650 49832 4014
rect 49988 3380 50016 10628
rect 50528 10610 50580 10616
rect 50252 10600 50304 10606
rect 50252 10542 50304 10548
rect 50264 10266 50292 10542
rect 50252 10260 50304 10266
rect 50252 10202 50304 10208
rect 50620 10056 50672 10062
rect 50620 9998 50672 10004
rect 50632 9722 50660 9998
rect 50620 9716 50672 9722
rect 50620 9658 50672 9664
rect 50160 9376 50212 9382
rect 50160 9318 50212 9324
rect 50068 9104 50120 9110
rect 50068 9046 50120 9052
rect 50080 8294 50108 9046
rect 50172 9042 50200 9318
rect 50160 9036 50212 9042
rect 50160 8978 50212 8984
rect 50172 8430 50200 8978
rect 50160 8424 50212 8430
rect 50160 8366 50212 8372
rect 50436 8424 50488 8430
rect 50436 8366 50488 8372
rect 50068 8288 50120 8294
rect 50068 8230 50120 8236
rect 50172 7206 50200 8366
rect 50448 8090 50476 8366
rect 50436 8084 50488 8090
rect 50436 8026 50488 8032
rect 50620 7744 50672 7750
rect 50620 7686 50672 7692
rect 50160 7200 50212 7206
rect 50160 7142 50212 7148
rect 50172 6322 50200 7142
rect 50160 6316 50212 6322
rect 50160 6258 50212 6264
rect 50436 6112 50488 6118
rect 50436 6054 50488 6060
rect 50448 5234 50476 6054
rect 50632 5778 50660 7686
rect 50620 5772 50672 5778
rect 50620 5714 50672 5720
rect 50436 5228 50488 5234
rect 50436 5170 50488 5176
rect 50252 5092 50304 5098
rect 50252 5034 50304 5040
rect 50160 4752 50212 4758
rect 50160 4694 50212 4700
rect 50172 4622 50200 4694
rect 50160 4616 50212 4622
rect 50160 4558 50212 4564
rect 50068 4480 50120 4486
rect 50068 4422 50120 4428
rect 50080 3534 50108 4422
rect 50172 3738 50200 4558
rect 50264 3942 50292 5034
rect 50724 4146 50752 11494
rect 51172 11008 51224 11014
rect 51172 10950 51224 10956
rect 51184 10674 51212 10950
rect 51172 10668 51224 10674
rect 51172 10610 51224 10616
rect 50804 10464 50856 10470
rect 50804 10406 50856 10412
rect 50816 9654 50844 10406
rect 51184 10146 51212 10610
rect 51092 10118 51212 10146
rect 50804 9648 50856 9654
rect 50804 9590 50856 9596
rect 51092 9518 51120 10118
rect 51172 9988 51224 9994
rect 51172 9930 51224 9936
rect 51080 9512 51132 9518
rect 51080 9454 51132 9460
rect 51184 9450 51212 9930
rect 51276 9518 51304 12135
rect 51356 12096 51408 12102
rect 51356 12038 51408 12044
rect 51264 9512 51316 9518
rect 51264 9454 51316 9460
rect 51172 9444 51224 9450
rect 51172 9386 51224 9392
rect 51276 8634 51304 9454
rect 51264 8628 51316 8634
rect 51264 8570 51316 8576
rect 51368 8090 51396 12038
rect 51908 11552 51960 11558
rect 51908 11494 51960 11500
rect 51504 11452 51812 11461
rect 51504 11450 51510 11452
rect 51566 11450 51590 11452
rect 51646 11450 51670 11452
rect 51726 11450 51750 11452
rect 51806 11450 51812 11452
rect 51566 11398 51568 11450
rect 51748 11398 51750 11450
rect 51504 11396 51510 11398
rect 51566 11396 51590 11398
rect 51646 11396 51670 11398
rect 51726 11396 51750 11398
rect 51806 11396 51812 11398
rect 51504 11387 51812 11396
rect 51920 11082 51948 11494
rect 51908 11076 51960 11082
rect 51908 11018 51960 11024
rect 52012 10810 52040 12294
rect 52092 12164 52144 12170
rect 52092 12106 52144 12112
rect 52000 10804 52052 10810
rect 52000 10746 52052 10752
rect 51504 10364 51812 10373
rect 51504 10362 51510 10364
rect 51566 10362 51590 10364
rect 51646 10362 51670 10364
rect 51726 10362 51750 10364
rect 51806 10362 51812 10364
rect 51566 10310 51568 10362
rect 51748 10310 51750 10362
rect 51504 10308 51510 10310
rect 51566 10308 51590 10310
rect 51646 10308 51670 10310
rect 51726 10308 51750 10310
rect 51806 10308 51812 10310
rect 51504 10299 51812 10308
rect 51724 10056 51776 10062
rect 51724 9998 51776 10004
rect 51908 10056 51960 10062
rect 51908 9998 51960 10004
rect 51736 9586 51764 9998
rect 51920 9654 51948 9998
rect 52000 9920 52052 9926
rect 52000 9862 52052 9868
rect 51908 9648 51960 9654
rect 51908 9590 51960 9596
rect 51724 9580 51776 9586
rect 51724 9522 51776 9528
rect 51736 9450 51764 9522
rect 51724 9444 51776 9450
rect 51724 9386 51776 9392
rect 51908 9376 51960 9382
rect 51908 9318 51960 9324
rect 51504 9276 51812 9285
rect 51504 9274 51510 9276
rect 51566 9274 51590 9276
rect 51646 9274 51670 9276
rect 51726 9274 51750 9276
rect 51806 9274 51812 9276
rect 51566 9222 51568 9274
rect 51748 9222 51750 9274
rect 51504 9220 51510 9222
rect 51566 9220 51590 9222
rect 51646 9220 51670 9222
rect 51726 9220 51750 9222
rect 51806 9220 51812 9222
rect 51504 9211 51812 9220
rect 51920 9042 51948 9318
rect 51908 9036 51960 9042
rect 51908 8978 51960 8984
rect 51908 8492 51960 8498
rect 51908 8434 51960 8440
rect 51504 8188 51812 8197
rect 51504 8186 51510 8188
rect 51566 8186 51590 8188
rect 51646 8186 51670 8188
rect 51726 8186 51750 8188
rect 51806 8186 51812 8188
rect 51566 8134 51568 8186
rect 51748 8134 51750 8186
rect 51504 8132 51510 8134
rect 51566 8132 51590 8134
rect 51646 8132 51670 8134
rect 51726 8132 51750 8134
rect 51806 8132 51812 8134
rect 51504 8123 51812 8132
rect 51080 8084 51132 8090
rect 51080 8026 51132 8032
rect 51356 8084 51408 8090
rect 51356 8026 51408 8032
rect 50988 7880 51040 7886
rect 50988 7822 51040 7828
rect 51000 7546 51028 7822
rect 50988 7540 51040 7546
rect 50988 7482 51040 7488
rect 50896 7200 50948 7206
rect 50896 7142 50948 7148
rect 50908 6390 50936 7142
rect 50896 6384 50948 6390
rect 50896 6326 50948 6332
rect 50804 6112 50856 6118
rect 50804 6054 50856 6060
rect 50816 5846 50844 6054
rect 50804 5840 50856 5846
rect 50804 5782 50856 5788
rect 50988 5024 51040 5030
rect 50988 4966 51040 4972
rect 51000 4214 51028 4966
rect 50988 4208 51040 4214
rect 50988 4150 51040 4156
rect 50436 4140 50488 4146
rect 50436 4082 50488 4088
rect 50712 4140 50764 4146
rect 50712 4082 50764 4088
rect 50448 4049 50476 4082
rect 50434 4040 50490 4049
rect 50434 3975 50490 3984
rect 50252 3936 50304 3942
rect 50252 3878 50304 3884
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 50068 3528 50120 3534
rect 50068 3470 50120 3476
rect 49988 3352 50200 3380
rect 50068 2984 50120 2990
rect 50068 2926 50120 2932
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49712 1442 49740 2382
rect 49528 1414 49740 1442
rect 49528 800 49556 1414
rect 50080 800 50108 2926
rect 50172 2650 50200 3352
rect 51000 2922 51028 4150
rect 51092 3126 51120 8026
rect 51356 7812 51408 7818
rect 51356 7754 51408 7760
rect 51264 7336 51316 7342
rect 51264 7278 51316 7284
rect 51276 5914 51304 7278
rect 51368 6882 51396 7754
rect 51504 7100 51812 7109
rect 51504 7098 51510 7100
rect 51566 7098 51590 7100
rect 51646 7098 51670 7100
rect 51726 7098 51750 7100
rect 51806 7098 51812 7100
rect 51566 7046 51568 7098
rect 51748 7046 51750 7098
rect 51504 7044 51510 7046
rect 51566 7044 51590 7046
rect 51646 7044 51670 7046
rect 51726 7044 51750 7046
rect 51806 7044 51812 7046
rect 51504 7035 51812 7044
rect 51368 6866 51488 6882
rect 51368 6860 51500 6866
rect 51368 6854 51448 6860
rect 51448 6802 51500 6808
rect 51632 6792 51684 6798
rect 51632 6734 51684 6740
rect 51644 6100 51672 6734
rect 51368 6072 51672 6100
rect 51264 5908 51316 5914
rect 51264 5850 51316 5856
rect 51368 5710 51396 6072
rect 51504 6012 51812 6021
rect 51504 6010 51510 6012
rect 51566 6010 51590 6012
rect 51646 6010 51670 6012
rect 51726 6010 51750 6012
rect 51806 6010 51812 6012
rect 51566 5958 51568 6010
rect 51748 5958 51750 6010
rect 51504 5956 51510 5958
rect 51566 5956 51590 5958
rect 51646 5956 51670 5958
rect 51726 5956 51750 5958
rect 51806 5956 51812 5958
rect 51504 5947 51812 5956
rect 51632 5772 51684 5778
rect 51632 5714 51684 5720
rect 51356 5704 51408 5710
rect 51356 5646 51408 5652
rect 51368 5370 51396 5646
rect 51644 5370 51672 5714
rect 51356 5364 51408 5370
rect 51356 5306 51408 5312
rect 51632 5364 51684 5370
rect 51632 5306 51684 5312
rect 51264 5228 51316 5234
rect 51264 5170 51316 5176
rect 51172 4140 51224 4146
rect 51172 4082 51224 4088
rect 51184 3466 51212 4082
rect 51172 3460 51224 3466
rect 51172 3402 51224 3408
rect 51080 3120 51132 3126
rect 51080 3062 51132 3068
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 51172 2848 51224 2854
rect 51172 2790 51224 2796
rect 51184 2650 51212 2790
rect 50160 2644 50212 2650
rect 50160 2586 50212 2592
rect 51172 2644 51224 2650
rect 51172 2586 51224 2592
rect 51276 2530 51304 5170
rect 51356 5024 51408 5030
rect 51356 4966 51408 4972
rect 51368 4826 51396 4966
rect 51504 4924 51812 4933
rect 51504 4922 51510 4924
rect 51566 4922 51590 4924
rect 51646 4922 51670 4924
rect 51726 4922 51750 4924
rect 51806 4922 51812 4924
rect 51566 4870 51568 4922
rect 51748 4870 51750 4922
rect 51504 4868 51510 4870
rect 51566 4868 51590 4870
rect 51646 4868 51670 4870
rect 51726 4868 51750 4870
rect 51806 4868 51812 4870
rect 51504 4859 51812 4868
rect 51356 4820 51408 4826
rect 51356 4762 51408 4768
rect 51816 4820 51868 4826
rect 51816 4762 51868 4768
rect 51828 4554 51856 4762
rect 51816 4548 51868 4554
rect 51816 4490 51868 4496
rect 51356 4004 51408 4010
rect 51356 3946 51408 3952
rect 51368 3058 51396 3946
rect 51504 3836 51812 3845
rect 51504 3834 51510 3836
rect 51566 3834 51590 3836
rect 51646 3834 51670 3836
rect 51726 3834 51750 3836
rect 51806 3834 51812 3836
rect 51566 3782 51568 3834
rect 51748 3782 51750 3834
rect 51504 3780 51510 3782
rect 51566 3780 51590 3782
rect 51646 3780 51670 3782
rect 51726 3780 51750 3782
rect 51806 3780 51812 3782
rect 51504 3771 51812 3780
rect 51920 3194 51948 8434
rect 52012 7546 52040 9862
rect 52000 7540 52052 7546
rect 52000 7482 52052 7488
rect 52000 7336 52052 7342
rect 52000 7278 52052 7284
rect 52012 6662 52040 7278
rect 52000 6656 52052 6662
rect 52000 6598 52052 6604
rect 52000 6316 52052 6322
rect 52000 6258 52052 6264
rect 52012 5778 52040 6258
rect 52000 5772 52052 5778
rect 52000 5714 52052 5720
rect 52000 5568 52052 5574
rect 52000 5510 52052 5516
rect 52012 5302 52040 5510
rect 52000 5296 52052 5302
rect 52000 5238 52052 5244
rect 52000 4140 52052 4146
rect 52000 4082 52052 4088
rect 51908 3188 51960 3194
rect 51908 3130 51960 3136
rect 52012 3058 52040 4082
rect 51356 3052 51408 3058
rect 51356 2994 51408 3000
rect 52000 3052 52052 3058
rect 52000 2994 52052 3000
rect 51724 2984 51776 2990
rect 52104 2938 52132 12106
rect 52196 8634 52224 15098
rect 52288 13870 52316 19654
rect 52564 18766 52592 24754
rect 52644 24200 52696 24206
rect 52644 24142 52696 24148
rect 52656 23322 52684 24142
rect 52736 24064 52788 24070
rect 52736 24006 52788 24012
rect 52644 23316 52696 23322
rect 52644 23258 52696 23264
rect 52748 23050 52776 24006
rect 53104 23520 53156 23526
rect 53104 23462 53156 23468
rect 52736 23044 52788 23050
rect 52736 22986 52788 22992
rect 53116 22778 53144 23462
rect 53208 22778 53236 25094
rect 53392 24954 53420 25298
rect 58726 25052 59034 25061
rect 58726 25050 58732 25052
rect 58788 25050 58812 25052
rect 58868 25050 58892 25052
rect 58948 25050 58972 25052
rect 59028 25050 59034 25052
rect 58788 24998 58790 25050
rect 58970 24998 58972 25050
rect 58726 24996 58732 24998
rect 58788 24996 58812 24998
rect 58868 24996 58892 24998
rect 58948 24996 58972 24998
rect 59028 24996 59034 24998
rect 58726 24987 59034 24996
rect 53380 24948 53432 24954
rect 53380 24890 53432 24896
rect 53288 24200 53340 24206
rect 53288 24142 53340 24148
rect 54392 24200 54444 24206
rect 54392 24142 54444 24148
rect 55312 24200 55364 24206
rect 55312 24142 55364 24148
rect 56876 24200 56928 24206
rect 56876 24142 56928 24148
rect 57244 24200 57296 24206
rect 57244 24142 57296 24148
rect 53300 23866 53328 24142
rect 53656 24064 53708 24070
rect 53656 24006 53708 24012
rect 53840 24064 53892 24070
rect 53840 24006 53892 24012
rect 53288 23860 53340 23866
rect 53288 23802 53340 23808
rect 53668 23662 53696 24006
rect 53656 23656 53708 23662
rect 53656 23598 53708 23604
rect 53564 22976 53616 22982
rect 53564 22918 53616 22924
rect 53104 22772 53156 22778
rect 53104 22714 53156 22720
rect 53196 22772 53248 22778
rect 53196 22714 53248 22720
rect 53576 22710 53604 22918
rect 53564 22704 53616 22710
rect 53564 22646 53616 22652
rect 52644 22568 52696 22574
rect 52644 22510 52696 22516
rect 52656 22098 52684 22510
rect 52736 22432 52788 22438
rect 52736 22374 52788 22380
rect 52644 22092 52696 22098
rect 52644 22034 52696 22040
rect 52748 21554 52776 22374
rect 52826 22128 52882 22137
rect 52826 22063 52882 22072
rect 52840 21622 52868 22063
rect 52828 21616 52880 21622
rect 52828 21558 52880 21564
rect 52736 21548 52788 21554
rect 52736 21490 52788 21496
rect 53564 20936 53616 20942
rect 53564 20878 53616 20884
rect 53196 20800 53248 20806
rect 53196 20742 53248 20748
rect 52736 20460 52788 20466
rect 52736 20402 52788 20408
rect 52748 20058 52776 20402
rect 52736 20052 52788 20058
rect 52736 19994 52788 20000
rect 52748 19514 52776 19994
rect 52736 19508 52788 19514
rect 52736 19450 52788 19456
rect 53208 19378 53236 20742
rect 53576 20602 53604 20878
rect 53564 20596 53616 20602
rect 53564 20538 53616 20544
rect 53196 19372 53248 19378
rect 53196 19314 53248 19320
rect 52460 18760 52512 18766
rect 52460 18702 52512 18708
rect 52552 18760 52604 18766
rect 52552 18702 52604 18708
rect 52472 17338 52500 18702
rect 52564 18426 52592 18702
rect 52552 18420 52604 18426
rect 52552 18362 52604 18368
rect 52552 18216 52604 18222
rect 52552 18158 52604 18164
rect 52564 17882 52592 18158
rect 53380 18080 53432 18086
rect 53380 18022 53432 18028
rect 52552 17876 52604 17882
rect 52552 17818 52604 17824
rect 52552 17740 52604 17746
rect 52552 17682 52604 17688
rect 52460 17332 52512 17338
rect 52460 17274 52512 17280
rect 52564 16998 52592 17682
rect 53392 17202 53420 18022
rect 53380 17196 53432 17202
rect 53380 17138 53432 17144
rect 52552 16992 52604 16998
rect 52552 16934 52604 16940
rect 52368 16652 52420 16658
rect 52368 16594 52420 16600
rect 52380 15026 52408 16594
rect 53472 15496 53524 15502
rect 53472 15438 53524 15444
rect 52460 15360 52512 15366
rect 52460 15302 52512 15308
rect 53380 15360 53432 15366
rect 53380 15302 53432 15308
rect 52472 15094 52500 15302
rect 52460 15088 52512 15094
rect 52460 15030 52512 15036
rect 52368 15020 52420 15026
rect 52368 14962 52420 14968
rect 52368 14884 52420 14890
rect 52368 14826 52420 14832
rect 52380 14482 52408 14826
rect 52368 14476 52420 14482
rect 52368 14418 52420 14424
rect 53392 14414 53420 15302
rect 53380 14408 53432 14414
rect 53380 14350 53432 14356
rect 53012 14272 53064 14278
rect 53012 14214 53064 14220
rect 53024 13870 53052 14214
rect 52276 13864 52328 13870
rect 52276 13806 52328 13812
rect 53012 13864 53064 13870
rect 53012 13806 53064 13812
rect 52276 12640 52328 12646
rect 52276 12582 52328 12588
rect 52184 8628 52236 8634
rect 52184 8570 52236 8576
rect 52288 7954 52316 12582
rect 52368 12232 52420 12238
rect 52368 12174 52420 12180
rect 52380 11354 52408 12174
rect 52920 12096 52972 12102
rect 52920 12038 52972 12044
rect 52460 11688 52512 11694
rect 52460 11630 52512 11636
rect 52472 11354 52500 11630
rect 52736 11552 52788 11558
rect 52736 11494 52788 11500
rect 52368 11348 52420 11354
rect 52368 11290 52420 11296
rect 52460 11348 52512 11354
rect 52460 11290 52512 11296
rect 52748 10742 52776 11494
rect 52932 11218 52960 12038
rect 53288 11688 53340 11694
rect 53288 11630 53340 11636
rect 52920 11212 52972 11218
rect 52920 11154 52972 11160
rect 52828 11008 52880 11014
rect 52828 10950 52880 10956
rect 52736 10736 52788 10742
rect 52736 10678 52788 10684
rect 52736 10600 52788 10606
rect 52840 10554 52868 10950
rect 52788 10548 52868 10554
rect 52736 10542 52868 10548
rect 52748 10526 52868 10542
rect 52748 9518 52776 10526
rect 52932 10062 52960 11154
rect 53104 10668 53156 10674
rect 53104 10610 53156 10616
rect 53116 10198 53144 10610
rect 53300 10470 53328 11630
rect 53484 11354 53512 15438
rect 53472 11348 53524 11354
rect 53472 11290 53524 11296
rect 53380 10804 53432 10810
rect 53380 10746 53432 10752
rect 53392 10606 53420 10746
rect 53380 10600 53432 10606
rect 53380 10542 53432 10548
rect 53288 10464 53340 10470
rect 53288 10406 53340 10412
rect 53392 10198 53420 10542
rect 53104 10192 53156 10198
rect 53104 10134 53156 10140
rect 53380 10192 53432 10198
rect 53380 10134 53432 10140
rect 52920 10056 52972 10062
rect 52920 9998 52972 10004
rect 52736 9512 52788 9518
rect 52736 9454 52788 9460
rect 53288 9512 53340 9518
rect 53288 9454 53340 9460
rect 52644 8288 52696 8294
rect 52644 8230 52696 8236
rect 52656 7954 52684 8230
rect 52276 7948 52328 7954
rect 52276 7890 52328 7896
rect 52644 7948 52696 7954
rect 52644 7890 52696 7896
rect 52748 7750 52776 9454
rect 53300 9178 53328 9454
rect 53288 9172 53340 9178
rect 53288 9114 53340 9120
rect 53196 8832 53248 8838
rect 53196 8774 53248 8780
rect 52828 8288 52880 8294
rect 52828 8230 52880 8236
rect 52840 7886 52868 8230
rect 52828 7880 52880 7886
rect 52828 7822 52880 7828
rect 52736 7744 52788 7750
rect 52736 7686 52788 7692
rect 52276 7200 52328 7206
rect 52276 7142 52328 7148
rect 52184 6656 52236 6662
rect 52184 6598 52236 6604
rect 52196 5846 52224 6598
rect 52288 6390 52316 7142
rect 52644 6792 52696 6798
rect 52644 6734 52696 6740
rect 52748 6746 52776 7686
rect 52840 6866 52868 7822
rect 52828 6860 52880 6866
rect 52828 6802 52880 6808
rect 52656 6458 52684 6734
rect 52748 6718 52868 6746
rect 52644 6452 52696 6458
rect 52644 6394 52696 6400
rect 52276 6384 52328 6390
rect 52276 6326 52328 6332
rect 52184 5840 52236 5846
rect 52184 5782 52236 5788
rect 52736 5704 52788 5710
rect 52736 5646 52788 5652
rect 52644 5568 52696 5574
rect 52644 5510 52696 5516
rect 52368 5296 52420 5302
rect 52368 5238 52420 5244
rect 52380 4162 52408 5238
rect 52656 4554 52684 5510
rect 52748 5370 52776 5646
rect 52840 5574 52868 6718
rect 52828 5568 52880 5574
rect 52828 5510 52880 5516
rect 52736 5364 52788 5370
rect 52736 5306 52788 5312
rect 52644 4548 52696 4554
rect 52644 4490 52696 4496
rect 52380 4146 52500 4162
rect 52840 4146 52868 5510
rect 53012 4616 53064 4622
rect 53012 4558 53064 4564
rect 52380 4140 52512 4146
rect 52380 4134 52460 4140
rect 52460 4082 52512 4088
rect 52828 4140 52880 4146
rect 52828 4082 52880 4088
rect 52368 3936 52420 3942
rect 52368 3878 52420 3884
rect 52380 3534 52408 3878
rect 53024 3534 53052 4558
rect 53208 4486 53236 8774
rect 53668 8498 53696 23598
rect 53852 23050 53880 24006
rect 54404 23866 54432 24142
rect 54576 24064 54628 24070
rect 54576 24006 54628 24012
rect 55220 24064 55272 24070
rect 55220 24006 55272 24012
rect 54392 23860 54444 23866
rect 54392 23802 54444 23808
rect 54588 23662 54616 24006
rect 55232 23798 55260 24006
rect 55220 23792 55272 23798
rect 55220 23734 55272 23740
rect 54576 23656 54628 23662
rect 54576 23598 54628 23604
rect 53840 23044 53892 23050
rect 53840 22986 53892 22992
rect 54300 20936 54352 20942
rect 54300 20878 54352 20884
rect 53840 20868 53892 20874
rect 53840 20810 53892 20816
rect 53852 19938 53880 20810
rect 54024 20800 54076 20806
rect 54024 20742 54076 20748
rect 54036 20602 54064 20742
rect 54024 20596 54076 20602
rect 54024 20538 54076 20544
rect 54024 20392 54076 20398
rect 54024 20334 54076 20340
rect 53852 19922 53972 19938
rect 53852 19916 53984 19922
rect 53852 19910 53932 19916
rect 53932 19858 53984 19864
rect 53840 18216 53892 18222
rect 53840 18158 53892 18164
rect 53852 17882 53880 18158
rect 53840 17876 53892 17882
rect 53840 17818 53892 17824
rect 54036 15706 54064 20334
rect 54116 19848 54168 19854
rect 54116 19790 54168 19796
rect 54128 19446 54156 19790
rect 54208 19712 54260 19718
rect 54208 19654 54260 19660
rect 54116 19440 54168 19446
rect 54116 19382 54168 19388
rect 54128 18970 54156 19382
rect 54220 19378 54248 19654
rect 54312 19514 54340 20878
rect 54484 20256 54536 20262
rect 54484 20198 54536 20204
rect 54392 19780 54444 19786
rect 54392 19722 54444 19728
rect 54404 19514 54432 19722
rect 54496 19718 54524 20198
rect 54484 19712 54536 19718
rect 54484 19654 54536 19660
rect 54300 19508 54352 19514
rect 54300 19450 54352 19456
rect 54392 19508 54444 19514
rect 54392 19450 54444 19456
rect 54208 19372 54260 19378
rect 54208 19314 54260 19320
rect 54116 18964 54168 18970
rect 54116 18906 54168 18912
rect 54128 17202 54156 18906
rect 54484 17672 54536 17678
rect 54484 17614 54536 17620
rect 54208 17536 54260 17542
rect 54208 17478 54260 17484
rect 54116 17196 54168 17202
rect 54116 17138 54168 17144
rect 54128 16794 54156 17138
rect 54116 16788 54168 16794
rect 54116 16730 54168 16736
rect 54220 16046 54248 17478
rect 54496 17338 54524 17614
rect 54484 17332 54536 17338
rect 54484 17274 54536 17280
rect 54208 16040 54260 16046
rect 54208 15982 54260 15988
rect 54024 15700 54076 15706
rect 54024 15642 54076 15648
rect 54116 15496 54168 15502
rect 54116 15438 54168 15444
rect 54128 15162 54156 15438
rect 54116 15156 54168 15162
rect 54116 15098 54168 15104
rect 54220 15094 54248 15982
rect 54300 15360 54352 15366
rect 54300 15302 54352 15308
rect 54208 15088 54260 15094
rect 54208 15030 54260 15036
rect 54208 14952 54260 14958
rect 54208 14894 54260 14900
rect 54220 14822 54248 14894
rect 53840 14816 53892 14822
rect 53840 14758 53892 14764
rect 54208 14816 54260 14822
rect 54208 14758 54260 14764
rect 53852 12442 53880 14758
rect 54312 13938 54340 15302
rect 54300 13932 54352 13938
rect 54300 13874 54352 13880
rect 54116 12640 54168 12646
rect 54116 12582 54168 12588
rect 53840 12436 53892 12442
rect 53840 12378 53892 12384
rect 54128 11830 54156 12582
rect 54588 12434 54616 23598
rect 55324 23322 55352 24142
rect 56048 24064 56100 24070
rect 56048 24006 56100 24012
rect 56600 24064 56652 24070
rect 56600 24006 56652 24012
rect 55772 23724 55824 23730
rect 55772 23666 55824 23672
rect 55496 23520 55548 23526
rect 55496 23462 55548 23468
rect 55312 23316 55364 23322
rect 55312 23258 55364 23264
rect 55508 22642 55536 23462
rect 55784 23322 55812 23666
rect 55772 23316 55824 23322
rect 55772 23258 55824 23264
rect 55784 22778 55812 23258
rect 56060 23186 56088 24006
rect 56612 23798 56640 24006
rect 56600 23792 56652 23798
rect 56600 23734 56652 23740
rect 56324 23656 56376 23662
rect 56324 23598 56376 23604
rect 56048 23180 56100 23186
rect 56048 23122 56100 23128
rect 55956 23112 56008 23118
rect 55956 23054 56008 23060
rect 55772 22772 55824 22778
rect 55772 22714 55824 22720
rect 55496 22636 55548 22642
rect 55496 22578 55548 22584
rect 55968 22166 55996 23054
rect 56336 22642 56364 23598
rect 56508 23180 56560 23186
rect 56508 23122 56560 23128
rect 56324 22636 56376 22642
rect 56324 22578 56376 22584
rect 56520 22166 56548 23122
rect 56692 22976 56744 22982
rect 56692 22918 56744 22924
rect 55956 22160 56008 22166
rect 55956 22102 56008 22108
rect 56508 22160 56560 22166
rect 56508 22102 56560 22108
rect 55220 21888 55272 21894
rect 55220 21830 55272 21836
rect 55864 21888 55916 21894
rect 55864 21830 55916 21836
rect 55232 21622 55260 21830
rect 55404 21684 55456 21690
rect 55404 21626 55456 21632
rect 55220 21616 55272 21622
rect 55220 21558 55272 21564
rect 54852 20800 54904 20806
rect 54852 20742 54904 20748
rect 54864 20330 54892 20742
rect 54852 20324 54904 20330
rect 54852 20266 54904 20272
rect 55036 20052 55088 20058
rect 55036 19994 55088 20000
rect 55048 19378 55076 19994
rect 55036 19372 55088 19378
rect 55036 19314 55088 19320
rect 55232 17542 55260 21558
rect 55416 20466 55444 21626
rect 55772 21548 55824 21554
rect 55772 21490 55824 21496
rect 55680 20936 55732 20942
rect 55680 20878 55732 20884
rect 55404 20460 55456 20466
rect 55404 20402 55456 20408
rect 55220 17536 55272 17542
rect 55220 17478 55272 17484
rect 55232 17270 55260 17478
rect 54944 17264 54996 17270
rect 54944 17206 54996 17212
rect 55220 17264 55272 17270
rect 55220 17206 55272 17212
rect 55416 17218 55444 20402
rect 55588 20392 55640 20398
rect 55588 20334 55640 20340
rect 55600 19786 55628 20334
rect 55692 19854 55720 20878
rect 55784 20602 55812 21490
rect 55772 20596 55824 20602
rect 55772 20538 55824 20544
rect 55680 19848 55732 19854
rect 55680 19790 55732 19796
rect 55588 19780 55640 19786
rect 55588 19722 55640 19728
rect 55600 19514 55628 19722
rect 55588 19508 55640 19514
rect 55588 19450 55640 19456
rect 55692 19378 55720 19790
rect 55680 19372 55732 19378
rect 55680 19314 55732 19320
rect 54760 16448 54812 16454
rect 54760 16390 54812 16396
rect 54772 16182 54800 16390
rect 54760 16176 54812 16182
rect 54760 16118 54812 16124
rect 54852 15496 54904 15502
rect 54852 15438 54904 15444
rect 54864 15162 54892 15438
rect 54852 15156 54904 15162
rect 54852 15098 54904 15104
rect 54956 14550 54984 17206
rect 55416 17190 55536 17218
rect 55508 17134 55536 17190
rect 55496 17128 55548 17134
rect 55496 17070 55548 17076
rect 55876 17082 55904 21830
rect 55968 21690 55996 22102
rect 56048 22092 56100 22098
rect 56048 22034 56100 22040
rect 55956 21684 56008 21690
rect 55956 21626 56008 21632
rect 56060 20398 56088 22034
rect 56704 21690 56732 22918
rect 56888 21894 56916 24142
rect 57256 23322 57284 24142
rect 57336 24064 57388 24070
rect 57336 24006 57388 24012
rect 57244 23316 57296 23322
rect 57244 23258 57296 23264
rect 56968 23112 57020 23118
rect 56968 23054 57020 23060
rect 56980 22438 57008 23054
rect 57060 22976 57112 22982
rect 57060 22918 57112 22924
rect 56968 22432 57020 22438
rect 56968 22374 57020 22380
rect 56980 22030 57008 22374
rect 57072 22234 57100 22918
rect 57348 22710 57376 24006
rect 58726 23964 59034 23973
rect 58726 23962 58732 23964
rect 58788 23962 58812 23964
rect 58868 23962 58892 23964
rect 58948 23962 58972 23964
rect 59028 23962 59034 23964
rect 58788 23910 58790 23962
rect 58970 23910 58972 23962
rect 58726 23908 58732 23910
rect 58788 23908 58812 23910
rect 58868 23908 58892 23910
rect 58948 23908 58972 23910
rect 59028 23908 59034 23910
rect 58726 23899 59034 23908
rect 57612 23656 57664 23662
rect 57612 23598 57664 23604
rect 57624 22778 57652 23598
rect 58072 23588 58124 23594
rect 58072 23530 58124 23536
rect 57796 23520 57848 23526
rect 57796 23462 57848 23468
rect 57888 23520 57940 23526
rect 57888 23462 57940 23468
rect 57808 22982 57836 23462
rect 57900 23186 57928 23462
rect 57888 23180 57940 23186
rect 57888 23122 57940 23128
rect 57796 22976 57848 22982
rect 57796 22918 57848 22924
rect 57612 22772 57664 22778
rect 57612 22714 57664 22720
rect 57336 22704 57388 22710
rect 57336 22646 57388 22652
rect 57060 22228 57112 22234
rect 57060 22170 57112 22176
rect 57808 22030 57836 22918
rect 58084 22642 58112 23530
rect 58726 22876 59034 22885
rect 58726 22874 58732 22876
rect 58788 22874 58812 22876
rect 58868 22874 58892 22876
rect 58948 22874 58972 22876
rect 59028 22874 59034 22876
rect 58788 22822 58790 22874
rect 58970 22822 58972 22874
rect 58726 22820 58732 22822
rect 58788 22820 58812 22822
rect 58868 22820 58892 22822
rect 58948 22820 58972 22822
rect 59028 22820 59034 22822
rect 58726 22811 59034 22820
rect 58072 22636 58124 22642
rect 58072 22578 58124 22584
rect 56968 22024 57020 22030
rect 56968 21966 57020 21972
rect 57796 22024 57848 22030
rect 57796 21966 57848 21972
rect 57980 22024 58032 22030
rect 57980 21966 58032 21972
rect 56876 21888 56928 21894
rect 56876 21830 56928 21836
rect 57428 21888 57480 21894
rect 57428 21830 57480 21836
rect 56692 21684 56744 21690
rect 56692 21626 56744 21632
rect 56784 21344 56836 21350
rect 56784 21286 56836 21292
rect 56796 20874 56824 21286
rect 56784 20868 56836 20874
rect 56784 20810 56836 20816
rect 56324 20800 56376 20806
rect 56324 20742 56376 20748
rect 56336 20398 56364 20742
rect 56048 20392 56100 20398
rect 56048 20334 56100 20340
rect 56324 20392 56376 20398
rect 56324 20334 56376 20340
rect 56232 19372 56284 19378
rect 56232 19314 56284 19320
rect 56244 17746 56272 19314
rect 56232 17740 56284 17746
rect 56232 17682 56284 17688
rect 56244 17626 56272 17682
rect 55956 17604 56008 17610
rect 55956 17546 56008 17552
rect 56152 17598 56272 17626
rect 55968 17202 55996 17546
rect 55956 17196 56008 17202
rect 55956 17138 56008 17144
rect 55404 17060 55456 17066
rect 55404 17002 55456 17008
rect 55220 15496 55272 15502
rect 55220 15438 55272 15444
rect 55036 15428 55088 15434
rect 55036 15370 55088 15376
rect 55128 15428 55180 15434
rect 55128 15370 55180 15376
rect 55048 15162 55076 15370
rect 55036 15156 55088 15162
rect 55036 15098 55088 15104
rect 55140 15026 55168 15370
rect 55128 15020 55180 15026
rect 55128 14962 55180 14968
rect 55036 14952 55088 14958
rect 55036 14894 55088 14900
rect 54944 14544 54996 14550
rect 54944 14486 54996 14492
rect 54956 13938 54984 14486
rect 55048 14278 55076 14894
rect 55036 14272 55088 14278
rect 55036 14214 55088 14220
rect 54944 13932 54996 13938
rect 54944 13874 54996 13880
rect 54956 12986 54984 13874
rect 54944 12980 54996 12986
rect 54944 12922 54996 12928
rect 54668 12776 54720 12782
rect 54668 12718 54720 12724
rect 54680 12442 54708 12718
rect 54496 12406 54616 12434
rect 54668 12436 54720 12442
rect 54116 11824 54168 11830
rect 54116 11766 54168 11772
rect 53748 11688 53800 11694
rect 53748 11630 53800 11636
rect 53760 11218 53788 11630
rect 53748 11212 53800 11218
rect 53748 11154 53800 11160
rect 54300 10600 54352 10606
rect 54300 10542 54352 10548
rect 54312 10266 54340 10542
rect 54300 10260 54352 10266
rect 54300 10202 54352 10208
rect 53840 9376 53892 9382
rect 53840 9318 53892 9324
rect 53656 8492 53708 8498
rect 53656 8434 53708 8440
rect 53380 8424 53432 8430
rect 53380 8366 53432 8372
rect 53392 7546 53420 8366
rect 53852 7970 53880 9318
rect 54300 8900 54352 8906
rect 54300 8842 54352 8848
rect 54312 8498 54340 8842
rect 54300 8492 54352 8498
rect 54300 8434 54352 8440
rect 53760 7942 53880 7970
rect 53760 7818 53788 7942
rect 54312 7886 54340 8434
rect 54300 7880 54352 7886
rect 54300 7822 54352 7828
rect 53748 7812 53800 7818
rect 53748 7754 53800 7760
rect 54208 7812 54260 7818
rect 54208 7754 54260 7760
rect 53380 7540 53432 7546
rect 53380 7482 53432 7488
rect 54116 7404 54168 7410
rect 54116 7346 54168 7352
rect 53932 7200 53984 7206
rect 53932 7142 53984 7148
rect 53944 6866 53972 7142
rect 53932 6860 53984 6866
rect 53932 6802 53984 6808
rect 53380 6656 53432 6662
rect 53380 6598 53432 6604
rect 53392 5370 53420 6598
rect 54128 6254 54156 7346
rect 54220 7002 54248 7754
rect 54312 7546 54340 7822
rect 54300 7540 54352 7546
rect 54300 7482 54352 7488
rect 54300 7200 54352 7206
rect 54300 7142 54352 7148
rect 54208 6996 54260 7002
rect 54208 6938 54260 6944
rect 54312 6866 54340 7142
rect 54496 6905 54524 12406
rect 54668 12378 54720 12384
rect 54668 12096 54720 12102
rect 54668 12038 54720 12044
rect 54680 10674 54708 12038
rect 54668 10668 54720 10674
rect 54668 10610 54720 10616
rect 54680 9722 54708 10610
rect 55048 10606 55076 14214
rect 55232 14074 55260 15438
rect 55312 14952 55364 14958
rect 55312 14894 55364 14900
rect 55324 14618 55352 14894
rect 55312 14612 55364 14618
rect 55312 14554 55364 14560
rect 55220 14068 55272 14074
rect 55220 14010 55272 14016
rect 55128 12980 55180 12986
rect 55128 12922 55180 12928
rect 55140 12434 55168 12922
rect 55312 12436 55364 12442
rect 55140 12406 55312 12434
rect 55312 12378 55364 12384
rect 55312 12232 55364 12238
rect 55312 12174 55364 12180
rect 55324 11898 55352 12174
rect 55312 11892 55364 11898
rect 55312 11834 55364 11840
rect 55128 11008 55180 11014
rect 55128 10950 55180 10956
rect 55140 10606 55168 10950
rect 55036 10600 55088 10606
rect 55036 10542 55088 10548
rect 55128 10600 55180 10606
rect 55128 10542 55180 10548
rect 55416 10266 55444 17002
rect 55508 16794 55536 17070
rect 55876 17054 55996 17082
rect 55496 16788 55548 16794
rect 55496 16730 55548 16736
rect 55508 14498 55536 16730
rect 55864 16584 55916 16590
rect 55864 16526 55916 16532
rect 55876 16046 55904 16526
rect 55864 16040 55916 16046
rect 55864 15982 55916 15988
rect 55680 15904 55732 15910
rect 55680 15846 55732 15852
rect 55508 14482 55628 14498
rect 55508 14476 55640 14482
rect 55508 14470 55588 14476
rect 55588 14418 55640 14424
rect 55496 13864 55548 13870
rect 55496 13806 55548 13812
rect 55508 13530 55536 13806
rect 55600 13530 55628 14418
rect 55496 13524 55548 13530
rect 55496 13466 55548 13472
rect 55588 13524 55640 13530
rect 55588 13466 55640 13472
rect 55600 12986 55628 13466
rect 55588 12980 55640 12986
rect 55588 12922 55640 12928
rect 55600 11626 55628 12922
rect 55692 12434 55720 15846
rect 55692 12406 55812 12434
rect 55588 11620 55640 11626
rect 55588 11562 55640 11568
rect 55404 10260 55456 10266
rect 55404 10202 55456 10208
rect 55312 9988 55364 9994
rect 55312 9930 55364 9936
rect 54668 9716 54720 9722
rect 54668 9658 54720 9664
rect 54680 7546 54708 9658
rect 54760 9376 54812 9382
rect 54760 9318 54812 9324
rect 54772 8634 54800 9318
rect 54760 8628 54812 8634
rect 54760 8570 54812 8576
rect 55324 8362 55352 9930
rect 55312 8356 55364 8362
rect 55312 8298 55364 8304
rect 55036 7812 55088 7818
rect 55036 7754 55088 7760
rect 55048 7546 55076 7754
rect 55128 7744 55180 7750
rect 55128 7686 55180 7692
rect 55140 7546 55168 7686
rect 54668 7540 54720 7546
rect 54668 7482 54720 7488
rect 55036 7540 55088 7546
rect 55036 7482 55088 7488
rect 55128 7540 55180 7546
rect 55128 7482 55180 7488
rect 54852 7336 54904 7342
rect 54852 7278 54904 7284
rect 54482 6896 54538 6905
rect 54300 6860 54352 6866
rect 54482 6831 54538 6840
rect 54300 6802 54352 6808
rect 54116 6248 54168 6254
rect 54116 6190 54168 6196
rect 54864 6118 54892 7278
rect 55128 6792 55180 6798
rect 55128 6734 55180 6740
rect 54852 6112 54904 6118
rect 54852 6054 54904 6060
rect 54944 6112 54996 6118
rect 54944 6054 54996 6060
rect 54668 5568 54720 5574
rect 54668 5510 54720 5516
rect 53380 5364 53432 5370
rect 53380 5306 53432 5312
rect 53564 5228 53616 5234
rect 53564 5170 53616 5176
rect 53932 5228 53984 5234
rect 53932 5170 53984 5176
rect 53196 4480 53248 4486
rect 53196 4422 53248 4428
rect 53576 4282 53604 5170
rect 53840 4820 53892 4826
rect 53840 4762 53892 4768
rect 53656 4752 53708 4758
rect 53656 4694 53708 4700
rect 53564 4276 53616 4282
rect 53564 4218 53616 4224
rect 53380 4140 53432 4146
rect 53380 4082 53432 4088
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 52184 3460 52236 3466
rect 52184 3402 52236 3408
rect 51776 2932 51948 2938
rect 51724 2926 51948 2932
rect 51736 2910 51948 2926
rect 51504 2748 51812 2757
rect 51504 2746 51510 2748
rect 51566 2746 51590 2748
rect 51646 2746 51670 2748
rect 51726 2746 51750 2748
rect 51806 2746 51812 2748
rect 51566 2694 51568 2746
rect 51748 2694 51750 2746
rect 51504 2692 51510 2694
rect 51566 2692 51590 2694
rect 51646 2692 51670 2694
rect 51726 2692 51750 2694
rect 51806 2692 51812 2694
rect 51504 2683 51812 2692
rect 51184 2502 51304 2530
rect 50632 2378 50844 2394
rect 50632 2372 50856 2378
rect 50632 2366 50804 2372
rect 50632 800 50660 2366
rect 50804 2314 50856 2320
rect 51184 800 51212 2502
rect 51920 1578 51948 2910
rect 52012 2910 52132 2938
rect 52012 2650 52040 2910
rect 52196 2774 52224 3402
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 53104 3392 53156 3398
rect 53104 3334 53156 3340
rect 52564 3126 52592 3334
rect 53116 3126 53144 3334
rect 52552 3120 52604 3126
rect 52552 3062 52604 3068
rect 53104 3120 53156 3126
rect 53104 3062 53156 3068
rect 52104 2746 52224 2774
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52104 2446 52132 2746
rect 52460 2508 52512 2514
rect 52460 2450 52512 2456
rect 52092 2440 52144 2446
rect 52092 2382 52144 2388
rect 51736 1550 51948 1578
rect 51736 800 51764 1550
rect 52472 1442 52500 2450
rect 52564 2446 52592 3062
rect 53392 2650 53420 4082
rect 53576 3126 53604 4218
rect 53668 3126 53696 4694
rect 53748 4616 53800 4622
rect 53748 4558 53800 4564
rect 53564 3120 53616 3126
rect 53564 3062 53616 3068
rect 53656 3120 53708 3126
rect 53656 3062 53708 3068
rect 53760 2990 53788 4558
rect 53852 3738 53880 4762
rect 53944 4282 53972 5170
rect 54680 5030 54708 5510
rect 54668 5024 54720 5030
rect 54668 4966 54720 4972
rect 54852 5024 54904 5030
rect 54852 4966 54904 4972
rect 54680 4826 54708 4966
rect 54668 4820 54720 4826
rect 54668 4762 54720 4768
rect 54864 4622 54892 4966
rect 54852 4616 54904 4622
rect 54852 4558 54904 4564
rect 54116 4480 54168 4486
rect 54116 4422 54168 4428
rect 54300 4480 54352 4486
rect 54300 4422 54352 4428
rect 53932 4276 53984 4282
rect 53932 4218 53984 4224
rect 53840 3732 53892 3738
rect 53840 3674 53892 3680
rect 53944 3074 53972 4218
rect 54128 4146 54156 4422
rect 54312 4146 54340 4422
rect 54496 4146 54616 4162
rect 54116 4140 54168 4146
rect 54116 4082 54168 4088
rect 54300 4140 54352 4146
rect 54300 4082 54352 4088
rect 54496 4140 54628 4146
rect 54496 4134 54576 4140
rect 54300 3936 54352 3942
rect 54300 3878 54352 3884
rect 54312 3466 54340 3878
rect 54300 3460 54352 3466
rect 54300 3402 54352 3408
rect 53852 3058 53972 3074
rect 53840 3052 53972 3058
rect 53892 3046 53972 3052
rect 53840 2994 53892 3000
rect 53748 2984 53800 2990
rect 53748 2926 53800 2932
rect 54208 2984 54260 2990
rect 54208 2926 54260 2932
rect 53380 2644 53432 2650
rect 53380 2586 53432 2592
rect 52552 2440 52604 2446
rect 52552 2382 52604 2388
rect 53380 2440 53432 2446
rect 53380 2382 53432 2388
rect 52920 2372 52972 2378
rect 52920 2314 52972 2320
rect 52288 1414 52500 1442
rect 52288 800 52316 1414
rect 52932 1306 52960 2314
rect 52840 1278 52960 1306
rect 52840 800 52868 1278
rect 53392 800 53420 2382
rect 53944 870 54064 898
rect 53944 800 53972 870
rect 47412 734 47716 762
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54036 762 54064 870
rect 54220 762 54248 2926
rect 54496 800 54524 4134
rect 54576 4082 54628 4088
rect 54864 4078 54892 4558
rect 54852 4072 54904 4078
rect 54574 4040 54630 4049
rect 54852 4014 54904 4020
rect 54574 3975 54630 3984
rect 54588 3942 54616 3975
rect 54576 3936 54628 3942
rect 54576 3878 54628 3884
rect 54956 3398 54984 6054
rect 55140 5914 55168 6734
rect 55416 6458 55444 10202
rect 55600 9654 55628 11562
rect 55588 9648 55640 9654
rect 55588 9590 55640 9596
rect 55496 9512 55548 9518
rect 55496 9454 55548 9460
rect 55508 8634 55536 9454
rect 55600 9178 55628 9590
rect 55588 9172 55640 9178
rect 55588 9114 55640 9120
rect 55496 8628 55548 8634
rect 55496 8570 55548 8576
rect 55600 8514 55628 9114
rect 55600 8486 55720 8514
rect 55692 8430 55720 8486
rect 55680 8424 55732 8430
rect 55680 8366 55732 8372
rect 55588 6656 55640 6662
rect 55588 6598 55640 6604
rect 55404 6452 55456 6458
rect 55404 6394 55456 6400
rect 55496 6248 55548 6254
rect 55496 6190 55548 6196
rect 55404 6112 55456 6118
rect 55404 6054 55456 6060
rect 55128 5908 55180 5914
rect 55128 5850 55180 5856
rect 55140 5234 55168 5850
rect 55416 5234 55444 6054
rect 55508 5370 55536 6190
rect 55600 5370 55628 6598
rect 55784 6225 55812 12406
rect 55864 11144 55916 11150
rect 55864 11086 55916 11092
rect 55876 10810 55904 11086
rect 55864 10804 55916 10810
rect 55864 10746 55916 10752
rect 55968 8974 55996 17054
rect 56152 16658 56180 17598
rect 56336 17490 56364 20334
rect 56692 20256 56744 20262
rect 56692 20198 56744 20204
rect 56508 19780 56560 19786
rect 56508 19722 56560 19728
rect 56520 18970 56548 19722
rect 56704 19514 56732 20198
rect 56692 19508 56744 19514
rect 56692 19450 56744 19456
rect 56796 19394 56824 20810
rect 57440 20602 57468 21830
rect 57612 21480 57664 21486
rect 57612 21422 57664 21428
rect 57624 21146 57652 21422
rect 57612 21140 57664 21146
rect 57612 21082 57664 21088
rect 57808 20890 57836 21966
rect 57992 21690 58020 21966
rect 58726 21788 59034 21797
rect 58726 21786 58732 21788
rect 58788 21786 58812 21788
rect 58868 21786 58892 21788
rect 58948 21786 58972 21788
rect 59028 21786 59034 21788
rect 58788 21734 58790 21786
rect 58970 21734 58972 21786
rect 58726 21732 58732 21734
rect 58788 21732 58812 21734
rect 58868 21732 58892 21734
rect 58948 21732 58972 21734
rect 59028 21732 59034 21734
rect 58726 21723 59034 21732
rect 57980 21684 58032 21690
rect 57980 21626 58032 21632
rect 57888 21344 57940 21350
rect 57888 21286 57940 21292
rect 57900 21146 57928 21286
rect 57888 21140 57940 21146
rect 57888 21082 57940 21088
rect 57808 20862 58020 20890
rect 57992 20806 58020 20862
rect 57520 20800 57572 20806
rect 57520 20742 57572 20748
rect 57980 20800 58032 20806
rect 57980 20742 58032 20748
rect 58072 20800 58124 20806
rect 58072 20742 58124 20748
rect 57428 20596 57480 20602
rect 57428 20538 57480 20544
rect 57532 20466 57560 20742
rect 57520 20460 57572 20466
rect 57520 20402 57572 20408
rect 56968 20392 57020 20398
rect 56968 20334 57020 20340
rect 56980 19854 57008 20334
rect 57428 20324 57480 20330
rect 57428 20266 57480 20272
rect 56968 19848 57020 19854
rect 56968 19790 57020 19796
rect 56980 19514 57008 19790
rect 56968 19508 57020 19514
rect 56968 19450 57020 19456
rect 56704 19366 56824 19394
rect 56508 18964 56560 18970
rect 56508 18906 56560 18912
rect 56600 18624 56652 18630
rect 56600 18566 56652 18572
rect 56508 18148 56560 18154
rect 56508 18090 56560 18096
rect 56244 17462 56364 17490
rect 56140 16652 56192 16658
rect 56140 16594 56192 16600
rect 56152 15026 56180 16594
rect 56244 16130 56272 17462
rect 56520 17338 56548 18090
rect 56612 17678 56640 18566
rect 56600 17672 56652 17678
rect 56600 17614 56652 17620
rect 56600 17536 56652 17542
rect 56600 17478 56652 17484
rect 56508 17332 56560 17338
rect 56508 17274 56560 17280
rect 56612 17218 56640 17478
rect 56520 17190 56640 17218
rect 56520 17134 56548 17190
rect 56324 17128 56376 17134
rect 56324 17070 56376 17076
rect 56508 17128 56560 17134
rect 56508 17070 56560 17076
rect 56336 16250 56364 17070
rect 56508 16992 56560 16998
rect 56508 16934 56560 16940
rect 56324 16244 56376 16250
rect 56324 16186 56376 16192
rect 56244 16102 56364 16130
rect 56232 15360 56284 15366
rect 56232 15302 56284 15308
rect 56244 15094 56272 15302
rect 56232 15088 56284 15094
rect 56232 15030 56284 15036
rect 56140 15020 56192 15026
rect 56140 14962 56192 14968
rect 56048 14884 56100 14890
rect 56048 14826 56100 14832
rect 56060 14482 56088 14826
rect 56244 14482 56272 15030
rect 56336 14498 56364 16102
rect 56520 14618 56548 16934
rect 56508 14612 56560 14618
rect 56508 14554 56560 14560
rect 56048 14476 56100 14482
rect 56048 14418 56100 14424
rect 56232 14476 56284 14482
rect 56336 14470 56548 14498
rect 56232 14418 56284 14424
rect 56140 13864 56192 13870
rect 56140 13806 56192 13812
rect 56152 13530 56180 13806
rect 56140 13524 56192 13530
rect 56140 13466 56192 13472
rect 56520 12434 56548 14470
rect 56704 13394 56732 19366
rect 57152 18760 57204 18766
rect 57152 18702 57204 18708
rect 57164 18426 57192 18702
rect 57152 18420 57204 18426
rect 57152 18362 57204 18368
rect 56968 18284 57020 18290
rect 56968 18226 57020 18232
rect 56876 18216 56928 18222
rect 56876 18158 56928 18164
rect 56888 16114 56916 18158
rect 56980 17202 57008 18226
rect 56968 17196 57020 17202
rect 56968 17138 57020 17144
rect 57060 17128 57112 17134
rect 57060 17070 57112 17076
rect 56876 16108 56928 16114
rect 56876 16050 56928 16056
rect 56888 15366 56916 16050
rect 57072 16046 57100 17070
rect 57152 16652 57204 16658
rect 57152 16594 57204 16600
rect 57164 16250 57192 16594
rect 57152 16244 57204 16250
rect 57152 16186 57204 16192
rect 57060 16040 57112 16046
rect 57060 15982 57112 15988
rect 57152 15564 57204 15570
rect 57152 15506 57204 15512
rect 56784 15360 56836 15366
rect 56784 15302 56836 15308
rect 56876 15360 56928 15366
rect 56876 15302 56928 15308
rect 56796 14482 56824 15302
rect 56784 14476 56836 14482
rect 56784 14418 56836 14424
rect 56692 13388 56744 13394
rect 56692 13330 56744 13336
rect 56784 13388 56836 13394
rect 56784 13330 56836 13336
rect 56692 12640 56744 12646
rect 56692 12582 56744 12588
rect 56428 12406 56548 12434
rect 56600 12436 56652 12442
rect 56232 12232 56284 12238
rect 56232 12174 56284 12180
rect 56140 12164 56192 12170
rect 56140 12106 56192 12112
rect 56152 11762 56180 12106
rect 56244 11898 56272 12174
rect 56232 11892 56284 11898
rect 56232 11834 56284 11840
rect 56140 11756 56192 11762
rect 56140 11698 56192 11704
rect 56244 11218 56272 11834
rect 56232 11212 56284 11218
rect 56232 11154 56284 11160
rect 56324 10260 56376 10266
rect 56324 10202 56376 10208
rect 56140 9580 56192 9586
rect 56140 9522 56192 9528
rect 55956 8968 56008 8974
rect 55956 8910 56008 8916
rect 56152 8498 56180 9522
rect 56336 9518 56364 10202
rect 56324 9512 56376 9518
rect 56324 9454 56376 9460
rect 56232 9376 56284 9382
rect 56232 9318 56284 9324
rect 56244 9178 56272 9318
rect 56232 9172 56284 9178
rect 56232 9114 56284 9120
rect 56232 8968 56284 8974
rect 56232 8910 56284 8916
rect 56140 8492 56192 8498
rect 56140 8434 56192 8440
rect 56244 7886 56272 8910
rect 56232 7880 56284 7886
rect 56232 7822 56284 7828
rect 55770 6216 55826 6225
rect 55770 6151 55826 6160
rect 56140 6112 56192 6118
rect 56140 6054 56192 6060
rect 56152 5642 56180 6054
rect 56244 5692 56272 7822
rect 56324 7200 56376 7206
rect 56324 7142 56376 7148
rect 56336 6866 56364 7142
rect 56324 6860 56376 6866
rect 56324 6802 56376 6808
rect 56428 6361 56456 12406
rect 56600 12378 56652 12384
rect 56508 11688 56560 11694
rect 56508 11630 56560 11636
rect 56520 10810 56548 11630
rect 56612 11626 56640 12378
rect 56704 12238 56732 12582
rect 56692 12232 56744 12238
rect 56692 12174 56744 12180
rect 56600 11620 56652 11626
rect 56600 11562 56652 11568
rect 56692 11552 56744 11558
rect 56692 11494 56744 11500
rect 56508 10804 56560 10810
rect 56508 10746 56560 10752
rect 56600 9172 56652 9178
rect 56600 9114 56652 9120
rect 56508 8424 56560 8430
rect 56508 8366 56560 8372
rect 56520 7546 56548 8366
rect 56612 7886 56640 9114
rect 56600 7880 56652 7886
rect 56600 7822 56652 7828
rect 56704 7546 56732 11494
rect 56796 10606 56824 13330
rect 56888 13190 56916 15302
rect 56968 14408 57020 14414
rect 56968 14350 57020 14356
rect 56980 13326 57008 14350
rect 56968 13320 57020 13326
rect 56968 13262 57020 13268
rect 56876 13184 56928 13190
rect 56876 13126 56928 13132
rect 56968 12844 57020 12850
rect 56968 12786 57020 12792
rect 56876 11620 56928 11626
rect 56876 11562 56928 11568
rect 56784 10600 56836 10606
rect 56784 10542 56836 10548
rect 56784 8628 56836 8634
rect 56784 8570 56836 8576
rect 56796 7546 56824 8570
rect 56888 8362 56916 11562
rect 56980 10674 57008 12786
rect 57164 12782 57192 15506
rect 57336 15360 57388 15366
rect 57336 15302 57388 15308
rect 57348 15094 57376 15302
rect 57336 15088 57388 15094
rect 57336 15030 57388 15036
rect 57244 14272 57296 14278
rect 57244 14214 57296 14220
rect 57060 12776 57112 12782
rect 57060 12718 57112 12724
rect 57152 12776 57204 12782
rect 57152 12718 57204 12724
rect 57072 12102 57100 12718
rect 57060 12096 57112 12102
rect 57060 12038 57112 12044
rect 57072 11898 57100 12038
rect 57060 11892 57112 11898
rect 57060 11834 57112 11840
rect 57060 11688 57112 11694
rect 57060 11630 57112 11636
rect 57072 10810 57100 11630
rect 57060 10804 57112 10810
rect 57060 10746 57112 10752
rect 56968 10668 57020 10674
rect 56968 10610 57020 10616
rect 56980 10010 57008 10610
rect 57256 10130 57284 14214
rect 57440 11558 57468 20266
rect 57992 19938 58020 20742
rect 58084 20534 58112 20742
rect 58726 20700 59034 20709
rect 58726 20698 58732 20700
rect 58788 20698 58812 20700
rect 58868 20698 58892 20700
rect 58948 20698 58972 20700
rect 59028 20698 59034 20700
rect 58788 20646 58790 20698
rect 58970 20646 58972 20698
rect 58726 20644 58732 20646
rect 58788 20644 58812 20646
rect 58868 20644 58892 20646
rect 58948 20644 58972 20646
rect 59028 20644 59034 20646
rect 58726 20635 59034 20644
rect 58072 20528 58124 20534
rect 58072 20470 58124 20476
rect 58164 20052 58216 20058
rect 58164 19994 58216 20000
rect 57992 19910 58112 19938
rect 58084 19718 58112 19910
rect 58072 19712 58124 19718
rect 58072 19654 58124 19660
rect 57612 19168 57664 19174
rect 57612 19110 57664 19116
rect 57520 16448 57572 16454
rect 57520 16390 57572 16396
rect 57532 16250 57560 16390
rect 57520 16244 57572 16250
rect 57520 16186 57572 16192
rect 57624 15026 57652 19110
rect 57704 18216 57756 18222
rect 57704 18158 57756 18164
rect 57716 17882 57744 18158
rect 57704 17876 57756 17882
rect 57704 17818 57756 17824
rect 57796 15156 57848 15162
rect 57796 15098 57848 15104
rect 57612 15020 57664 15026
rect 57612 14962 57664 14968
rect 57704 14816 57756 14822
rect 57704 14758 57756 14764
rect 57716 14006 57744 14758
rect 57808 14482 57836 15098
rect 57796 14476 57848 14482
rect 57796 14418 57848 14424
rect 57704 14000 57756 14006
rect 57704 13942 57756 13948
rect 57520 13184 57572 13190
rect 57520 13126 57572 13132
rect 57428 11552 57480 11558
rect 57428 11494 57480 11500
rect 57336 11144 57388 11150
rect 57336 11086 57388 11092
rect 57348 10810 57376 11086
rect 57336 10804 57388 10810
rect 57336 10746 57388 10752
rect 57440 10690 57468 11494
rect 57348 10662 57468 10690
rect 57244 10124 57296 10130
rect 57244 10066 57296 10072
rect 56980 9982 57100 10010
rect 56968 9920 57020 9926
rect 56968 9862 57020 9868
rect 56876 8356 56928 8362
rect 56876 8298 56928 8304
rect 56508 7540 56560 7546
rect 56508 7482 56560 7488
rect 56692 7540 56744 7546
rect 56692 7482 56744 7488
rect 56784 7540 56836 7546
rect 56784 7482 56836 7488
rect 56600 6792 56652 6798
rect 56600 6734 56652 6740
rect 56414 6352 56470 6361
rect 56414 6287 56470 6296
rect 56324 5704 56376 5710
rect 56244 5664 56324 5692
rect 56324 5646 56376 5652
rect 56140 5636 56192 5642
rect 56140 5578 56192 5584
rect 55496 5364 55548 5370
rect 55496 5306 55548 5312
rect 55588 5364 55640 5370
rect 55588 5306 55640 5312
rect 56336 5234 56364 5646
rect 55128 5228 55180 5234
rect 55128 5170 55180 5176
rect 55404 5228 55456 5234
rect 55404 5170 55456 5176
rect 56324 5228 56376 5234
rect 56324 5170 56376 5176
rect 56416 5228 56468 5234
rect 56416 5170 56468 5176
rect 56324 5092 56376 5098
rect 56324 5034 56376 5040
rect 56336 4690 56364 5034
rect 56428 4826 56456 5170
rect 56416 4820 56468 4826
rect 56416 4762 56468 4768
rect 56324 4684 56376 4690
rect 56324 4626 56376 4632
rect 55220 4480 55272 4486
rect 55220 4422 55272 4428
rect 55232 3534 55260 4422
rect 56336 4282 56364 4626
rect 56612 4282 56640 6734
rect 56876 6724 56928 6730
rect 56876 6666 56928 6672
rect 56692 5568 56744 5574
rect 56692 5510 56744 5516
rect 56704 4690 56732 5510
rect 56888 4706 56916 6666
rect 56980 6458 57008 9862
rect 57072 9722 57100 9982
rect 57060 9716 57112 9722
rect 57060 9658 57112 9664
rect 57072 7750 57100 9658
rect 57152 9444 57204 9450
rect 57152 9386 57204 9392
rect 57164 8974 57192 9386
rect 57152 8968 57204 8974
rect 57152 8910 57204 8916
rect 57164 8634 57192 8910
rect 57244 8900 57296 8906
rect 57244 8842 57296 8848
rect 57256 8634 57284 8842
rect 57152 8628 57204 8634
rect 57152 8570 57204 8576
rect 57244 8628 57296 8634
rect 57244 8570 57296 8576
rect 57060 7744 57112 7750
rect 57060 7686 57112 7692
rect 57072 7002 57100 7686
rect 57060 6996 57112 7002
rect 57060 6938 57112 6944
rect 57244 6656 57296 6662
rect 57244 6598 57296 6604
rect 56968 6452 57020 6458
rect 56968 6394 57020 6400
rect 57060 6112 57112 6118
rect 57060 6054 57112 6060
rect 57072 5710 57100 6054
rect 57060 5704 57112 5710
rect 57060 5646 57112 5652
rect 57256 5574 57284 6598
rect 57244 5568 57296 5574
rect 57244 5510 57296 5516
rect 56968 5024 57020 5030
rect 56968 4966 57020 4972
rect 56692 4684 56744 4690
rect 56692 4626 56744 4632
rect 56796 4678 56916 4706
rect 56324 4276 56376 4282
rect 56324 4218 56376 4224
rect 56600 4276 56652 4282
rect 56600 4218 56652 4224
rect 55404 3936 55456 3942
rect 55404 3878 55456 3884
rect 55128 3528 55180 3534
rect 55128 3470 55180 3476
rect 55220 3528 55272 3534
rect 55220 3470 55272 3476
rect 54944 3392 54996 3398
rect 54944 3334 54996 3340
rect 54956 3097 54984 3334
rect 54942 3088 54998 3097
rect 54942 3023 54998 3032
rect 55036 2984 55088 2990
rect 55036 2926 55088 2932
rect 55048 800 55076 2926
rect 55140 2650 55168 3470
rect 55416 3466 55444 3878
rect 56600 3732 56652 3738
rect 56600 3674 56652 3680
rect 55404 3460 55456 3466
rect 55404 3402 55456 3408
rect 56612 2650 56640 3674
rect 56796 2650 56824 4678
rect 56980 4146 57008 4966
rect 57152 4616 57204 4622
rect 57152 4558 57204 4564
rect 57164 4282 57192 4558
rect 57152 4276 57204 4282
rect 57152 4218 57204 4224
rect 56968 4140 57020 4146
rect 56968 4082 57020 4088
rect 56876 4072 56928 4078
rect 56876 4014 56928 4020
rect 56888 3398 56916 4014
rect 57164 3738 57192 4218
rect 57256 4214 57284 5510
rect 57348 4214 57376 10662
rect 57532 9568 57560 13126
rect 57808 12434 57836 14418
rect 57888 14408 57940 14414
rect 57888 14350 57940 14356
rect 57900 14006 57928 14350
rect 57888 14000 57940 14006
rect 57888 13942 57940 13948
rect 58084 12918 58112 19654
rect 58176 18834 58204 19994
rect 58440 19984 58492 19990
rect 58440 19926 58492 19932
rect 58452 19378 58480 19926
rect 58726 19612 59034 19621
rect 58726 19610 58732 19612
rect 58788 19610 58812 19612
rect 58868 19610 58892 19612
rect 58948 19610 58972 19612
rect 59028 19610 59034 19612
rect 58788 19558 58790 19610
rect 58970 19558 58972 19610
rect 58726 19556 58732 19558
rect 58788 19556 58812 19558
rect 58868 19556 58892 19558
rect 58948 19556 58972 19558
rect 59028 19556 59034 19558
rect 58726 19547 59034 19556
rect 58440 19372 58492 19378
rect 58440 19314 58492 19320
rect 58164 18828 58216 18834
rect 58164 18770 58216 18776
rect 58726 18524 59034 18533
rect 58726 18522 58732 18524
rect 58788 18522 58812 18524
rect 58868 18522 58892 18524
rect 58948 18522 58972 18524
rect 59028 18522 59034 18524
rect 58788 18470 58790 18522
rect 58970 18470 58972 18522
rect 58726 18468 58732 18470
rect 58788 18468 58812 18470
rect 58868 18468 58892 18470
rect 58948 18468 58972 18470
rect 59028 18468 59034 18470
rect 58726 18459 59034 18468
rect 58726 17436 59034 17445
rect 58726 17434 58732 17436
rect 58788 17434 58812 17436
rect 58868 17434 58892 17436
rect 58948 17434 58972 17436
rect 59028 17434 59034 17436
rect 58788 17382 58790 17434
rect 58970 17382 58972 17434
rect 58726 17380 58732 17382
rect 58788 17380 58812 17382
rect 58868 17380 58892 17382
rect 58948 17380 58972 17382
rect 59028 17380 59034 17382
rect 58726 17371 59034 17380
rect 58726 16348 59034 16357
rect 58726 16346 58732 16348
rect 58788 16346 58812 16348
rect 58868 16346 58892 16348
rect 58948 16346 58972 16348
rect 59028 16346 59034 16348
rect 58788 16294 58790 16346
rect 58970 16294 58972 16346
rect 58726 16292 58732 16294
rect 58788 16292 58812 16294
rect 58868 16292 58892 16294
rect 58948 16292 58972 16294
rect 59028 16292 59034 16294
rect 58726 16283 59034 16292
rect 58726 15260 59034 15269
rect 58726 15258 58732 15260
rect 58788 15258 58812 15260
rect 58868 15258 58892 15260
rect 58948 15258 58972 15260
rect 59028 15258 59034 15260
rect 58788 15206 58790 15258
rect 58970 15206 58972 15258
rect 58726 15204 58732 15206
rect 58788 15204 58812 15206
rect 58868 15204 58892 15206
rect 58948 15204 58972 15206
rect 59028 15204 59034 15206
rect 58726 15195 59034 15204
rect 58532 14816 58584 14822
rect 58532 14758 58584 14764
rect 58440 14068 58492 14074
rect 58440 14010 58492 14016
rect 58452 13394 58480 14010
rect 58440 13388 58492 13394
rect 58440 13330 58492 13336
rect 58072 12912 58124 12918
rect 58072 12854 58124 12860
rect 58440 12844 58492 12850
rect 58440 12786 58492 12792
rect 58452 12434 58480 12786
rect 57440 9540 57560 9568
rect 57716 12406 57836 12434
rect 58360 12406 58480 12434
rect 57440 6866 57468 9540
rect 57716 7342 57744 12406
rect 57796 8832 57848 8838
rect 57796 8774 57848 8780
rect 57808 7410 57836 8774
rect 57888 8424 57940 8430
rect 57888 8366 57940 8372
rect 57900 8090 57928 8366
rect 58164 8356 58216 8362
rect 58164 8298 58216 8304
rect 57888 8084 57940 8090
rect 57888 8026 57940 8032
rect 57888 7948 57940 7954
rect 57888 7890 57940 7896
rect 57900 7546 57928 7890
rect 58176 7886 58204 8298
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 58176 7546 58204 7822
rect 57888 7540 57940 7546
rect 57888 7482 57940 7488
rect 58164 7540 58216 7546
rect 58164 7482 58216 7488
rect 57796 7404 57848 7410
rect 57796 7346 57848 7352
rect 57704 7336 57756 7342
rect 57704 7278 57756 7284
rect 57428 6860 57480 6866
rect 57428 6802 57480 6808
rect 57612 6724 57664 6730
rect 57612 6666 57664 6672
rect 57704 6724 57756 6730
rect 57704 6666 57756 6672
rect 58256 6724 58308 6730
rect 58256 6666 58308 6672
rect 57244 4208 57296 4214
rect 57244 4150 57296 4156
rect 57336 4208 57388 4214
rect 57336 4150 57388 4156
rect 57428 4140 57480 4146
rect 57428 4082 57480 4088
rect 57152 3732 57204 3738
rect 57152 3674 57204 3680
rect 56876 3392 56928 3398
rect 56876 3334 56928 3340
rect 55128 2644 55180 2650
rect 55128 2586 55180 2592
rect 56600 2644 56652 2650
rect 56600 2586 56652 2592
rect 56784 2644 56836 2650
rect 56784 2586 56836 2592
rect 56784 2508 56836 2514
rect 56784 2450 56836 2456
rect 55600 2378 55720 2394
rect 56152 2378 56364 2394
rect 55600 2372 55732 2378
rect 55600 2366 55680 2372
rect 55600 800 55628 2366
rect 55680 2314 55732 2320
rect 56152 2372 56376 2378
rect 56152 2366 56324 2372
rect 56152 800 56180 2366
rect 56324 2314 56376 2320
rect 56796 1306 56824 2450
rect 56888 2446 56916 3334
rect 57244 2984 57296 2990
rect 57244 2926 57296 2932
rect 56968 2848 57020 2854
rect 56968 2790 57020 2796
rect 56980 2446 57008 2790
rect 56876 2440 56928 2446
rect 56876 2382 56928 2388
rect 56968 2440 57020 2446
rect 56968 2382 57020 2388
rect 56704 1278 56824 1306
rect 56704 800 56732 1278
rect 57256 800 57284 2926
rect 57440 2650 57468 4082
rect 57624 3942 57652 6666
rect 57716 5370 57744 6666
rect 58268 6458 58296 6666
rect 58256 6452 58308 6458
rect 58256 6394 58308 6400
rect 58360 5846 58388 12406
rect 58544 11762 58572 14758
rect 58726 14172 59034 14181
rect 58726 14170 58732 14172
rect 58788 14170 58812 14172
rect 58868 14170 58892 14172
rect 58948 14170 58972 14172
rect 59028 14170 59034 14172
rect 58788 14118 58790 14170
rect 58970 14118 58972 14170
rect 58726 14116 58732 14118
rect 58788 14116 58812 14118
rect 58868 14116 58892 14118
rect 58948 14116 58972 14118
rect 59028 14116 59034 14118
rect 58726 14107 59034 14116
rect 58726 13084 59034 13093
rect 58726 13082 58732 13084
rect 58788 13082 58812 13084
rect 58868 13082 58892 13084
rect 58948 13082 58972 13084
rect 59028 13082 59034 13084
rect 58788 13030 58790 13082
rect 58970 13030 58972 13082
rect 58726 13028 58732 13030
rect 58788 13028 58812 13030
rect 58868 13028 58892 13030
rect 58948 13028 58972 13030
rect 59028 13028 59034 13030
rect 58726 13019 59034 13028
rect 58726 11996 59034 12005
rect 58726 11994 58732 11996
rect 58788 11994 58812 11996
rect 58868 11994 58892 11996
rect 58948 11994 58972 11996
rect 59028 11994 59034 11996
rect 58788 11942 58790 11994
rect 58970 11942 58972 11994
rect 58726 11940 58732 11942
rect 58788 11940 58812 11942
rect 58868 11940 58892 11942
rect 58948 11940 58972 11942
rect 59028 11940 59034 11942
rect 58726 11931 59034 11940
rect 58532 11756 58584 11762
rect 58532 11698 58584 11704
rect 58440 11280 58492 11286
rect 58440 11222 58492 11228
rect 58452 10674 58480 11222
rect 58726 10908 59034 10917
rect 58726 10906 58732 10908
rect 58788 10906 58812 10908
rect 58868 10906 58892 10908
rect 58948 10906 58972 10908
rect 59028 10906 59034 10908
rect 58788 10854 58790 10906
rect 58970 10854 58972 10906
rect 58726 10852 58732 10854
rect 58788 10852 58812 10854
rect 58868 10852 58892 10854
rect 58948 10852 58972 10854
rect 59028 10852 59034 10854
rect 58726 10843 59034 10852
rect 58440 10668 58492 10674
rect 58440 10610 58492 10616
rect 58726 9820 59034 9829
rect 58726 9818 58732 9820
rect 58788 9818 58812 9820
rect 58868 9818 58892 9820
rect 58948 9818 58972 9820
rect 59028 9818 59034 9820
rect 58788 9766 58790 9818
rect 58970 9766 58972 9818
rect 58726 9764 58732 9766
rect 58788 9764 58812 9766
rect 58868 9764 58892 9766
rect 58948 9764 58972 9766
rect 59028 9764 59034 9766
rect 58726 9755 59034 9764
rect 58440 8968 58492 8974
rect 58440 8910 58492 8916
rect 58452 8090 58480 8910
rect 58726 8732 59034 8741
rect 58726 8730 58732 8732
rect 58788 8730 58812 8732
rect 58868 8730 58892 8732
rect 58948 8730 58972 8732
rect 59028 8730 59034 8732
rect 58788 8678 58790 8730
rect 58970 8678 58972 8730
rect 58726 8676 58732 8678
rect 58788 8676 58812 8678
rect 58868 8676 58892 8678
rect 58948 8676 58972 8678
rect 59028 8676 59034 8678
rect 58726 8667 59034 8676
rect 58440 8084 58492 8090
rect 58440 8026 58492 8032
rect 58726 7644 59034 7653
rect 58726 7642 58732 7644
rect 58788 7642 58812 7644
rect 58868 7642 58892 7644
rect 58948 7642 58972 7644
rect 59028 7642 59034 7644
rect 58788 7590 58790 7642
rect 58970 7590 58972 7642
rect 58726 7588 58732 7590
rect 58788 7588 58812 7590
rect 58868 7588 58892 7590
rect 58948 7588 58972 7590
rect 59028 7588 59034 7590
rect 58726 7579 59034 7588
rect 58440 6860 58492 6866
rect 58440 6802 58492 6808
rect 58348 5840 58400 5846
rect 58348 5782 58400 5788
rect 57704 5364 57756 5370
rect 57704 5306 57756 5312
rect 57612 3936 57664 3942
rect 57612 3878 57664 3884
rect 57716 3058 57744 5306
rect 58452 5234 58480 6802
rect 58726 6556 59034 6565
rect 58726 6554 58732 6556
rect 58788 6554 58812 6556
rect 58868 6554 58892 6556
rect 58948 6554 58972 6556
rect 59028 6554 59034 6556
rect 58788 6502 58790 6554
rect 58970 6502 58972 6554
rect 58726 6500 58732 6502
rect 58788 6500 58812 6502
rect 58868 6500 58892 6502
rect 58948 6500 58972 6502
rect 59028 6500 59034 6502
rect 58726 6491 59034 6500
rect 58532 5704 58584 5710
rect 58532 5646 58584 5652
rect 58440 5228 58492 5234
rect 58440 5170 58492 5176
rect 57888 5024 57940 5030
rect 57888 4966 57940 4972
rect 57900 4826 57928 4966
rect 57888 4820 57940 4826
rect 57888 4762 57940 4768
rect 57796 4548 57848 4554
rect 57796 4490 57848 4496
rect 57704 3052 57756 3058
rect 57704 2994 57756 3000
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 57808 800 57836 4490
rect 58256 3732 58308 3738
rect 58256 3674 58308 3680
rect 58268 3482 58296 3674
rect 58176 3466 58296 3482
rect 58164 3460 58296 3466
rect 58216 3454 58296 3460
rect 58164 3402 58216 3408
rect 58544 3194 58572 5646
rect 58726 5468 59034 5477
rect 58726 5466 58732 5468
rect 58788 5466 58812 5468
rect 58868 5466 58892 5468
rect 58948 5466 58972 5468
rect 59028 5466 59034 5468
rect 58788 5414 58790 5466
rect 58970 5414 58972 5466
rect 58726 5412 58732 5414
rect 58788 5412 58812 5414
rect 58868 5412 58892 5414
rect 58948 5412 58972 5414
rect 59028 5412 59034 5414
rect 58726 5403 59034 5412
rect 58624 4548 58676 4554
rect 58624 4490 58676 4496
rect 58532 3188 58584 3194
rect 58532 3130 58584 3136
rect 58348 2984 58400 2990
rect 58348 2926 58400 2932
rect 58360 800 58388 2926
rect 58636 1986 58664 4490
rect 58726 4380 59034 4389
rect 58726 4378 58732 4380
rect 58788 4378 58812 4380
rect 58868 4378 58892 4380
rect 58948 4378 58972 4380
rect 59028 4378 59034 4380
rect 58788 4326 58790 4378
rect 58970 4326 58972 4378
rect 58726 4324 58732 4326
rect 58788 4324 58812 4326
rect 58868 4324 58892 4326
rect 58948 4324 58972 4326
rect 59028 4324 59034 4326
rect 58726 4315 59034 4324
rect 58726 3292 59034 3301
rect 58726 3290 58732 3292
rect 58788 3290 58812 3292
rect 58868 3290 58892 3292
rect 58948 3290 58972 3292
rect 59028 3290 59034 3292
rect 58788 3238 58790 3290
rect 58970 3238 58972 3290
rect 58726 3236 58732 3238
rect 58788 3236 58812 3238
rect 58868 3236 58892 3238
rect 58948 3236 58972 3238
rect 59028 3236 59034 3238
rect 58726 3227 59034 3236
rect 58726 2204 59034 2213
rect 58726 2202 58732 2204
rect 58788 2202 58812 2204
rect 58868 2202 58892 2204
rect 58948 2202 58972 2204
rect 59028 2202 59034 2204
rect 58788 2150 58790 2202
rect 58970 2150 58972 2202
rect 58726 2148 58732 2150
rect 58788 2148 58812 2150
rect 58868 2148 58892 2150
rect 58948 2148 58972 2150
rect 59028 2148 59034 2150
rect 58726 2139 59034 2148
rect 58636 1958 58940 1986
rect 58912 800 58940 1958
rect 54036 734 54248 762
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
<< via2 >>
rect 8178 27770 8234 27772
rect 8258 27770 8314 27772
rect 8338 27770 8394 27772
rect 8418 27770 8474 27772
rect 8178 27718 8224 27770
rect 8224 27718 8234 27770
rect 8258 27718 8288 27770
rect 8288 27718 8300 27770
rect 8300 27718 8314 27770
rect 8338 27718 8352 27770
rect 8352 27718 8364 27770
rect 8364 27718 8394 27770
rect 8418 27718 8428 27770
rect 8428 27718 8474 27770
rect 8178 27716 8234 27718
rect 8258 27716 8314 27718
rect 8338 27716 8394 27718
rect 8418 27716 8474 27718
rect 22622 27770 22678 27772
rect 22702 27770 22758 27772
rect 22782 27770 22838 27772
rect 22862 27770 22918 27772
rect 22622 27718 22668 27770
rect 22668 27718 22678 27770
rect 22702 27718 22732 27770
rect 22732 27718 22744 27770
rect 22744 27718 22758 27770
rect 22782 27718 22796 27770
rect 22796 27718 22808 27770
rect 22808 27718 22838 27770
rect 22862 27718 22872 27770
rect 22872 27718 22918 27770
rect 22622 27716 22678 27718
rect 22702 27716 22758 27718
rect 22782 27716 22838 27718
rect 22862 27716 22918 27718
rect 37066 27770 37122 27772
rect 37146 27770 37202 27772
rect 37226 27770 37282 27772
rect 37306 27770 37362 27772
rect 37066 27718 37112 27770
rect 37112 27718 37122 27770
rect 37146 27718 37176 27770
rect 37176 27718 37188 27770
rect 37188 27718 37202 27770
rect 37226 27718 37240 27770
rect 37240 27718 37252 27770
rect 37252 27718 37282 27770
rect 37306 27718 37316 27770
rect 37316 27718 37362 27770
rect 37066 27716 37122 27718
rect 37146 27716 37202 27718
rect 37226 27716 37282 27718
rect 37306 27716 37362 27718
rect 51510 27770 51566 27772
rect 51590 27770 51646 27772
rect 51670 27770 51726 27772
rect 51750 27770 51806 27772
rect 51510 27718 51556 27770
rect 51556 27718 51566 27770
rect 51590 27718 51620 27770
rect 51620 27718 51632 27770
rect 51632 27718 51646 27770
rect 51670 27718 51684 27770
rect 51684 27718 51696 27770
rect 51696 27718 51726 27770
rect 51750 27718 51760 27770
rect 51760 27718 51806 27770
rect 51510 27716 51566 27718
rect 51590 27716 51646 27718
rect 51670 27716 51726 27718
rect 51750 27716 51806 27718
rect 15400 27226 15456 27228
rect 15480 27226 15536 27228
rect 15560 27226 15616 27228
rect 15640 27226 15696 27228
rect 15400 27174 15446 27226
rect 15446 27174 15456 27226
rect 15480 27174 15510 27226
rect 15510 27174 15522 27226
rect 15522 27174 15536 27226
rect 15560 27174 15574 27226
rect 15574 27174 15586 27226
rect 15586 27174 15616 27226
rect 15640 27174 15650 27226
rect 15650 27174 15696 27226
rect 15400 27172 15456 27174
rect 15480 27172 15536 27174
rect 15560 27172 15616 27174
rect 15640 27172 15696 27174
rect 29844 27226 29900 27228
rect 29924 27226 29980 27228
rect 30004 27226 30060 27228
rect 30084 27226 30140 27228
rect 29844 27174 29890 27226
rect 29890 27174 29900 27226
rect 29924 27174 29954 27226
rect 29954 27174 29966 27226
rect 29966 27174 29980 27226
rect 30004 27174 30018 27226
rect 30018 27174 30030 27226
rect 30030 27174 30060 27226
rect 30084 27174 30094 27226
rect 30094 27174 30140 27226
rect 29844 27172 29900 27174
rect 29924 27172 29980 27174
rect 30004 27172 30060 27174
rect 30084 27172 30140 27174
rect 44288 27226 44344 27228
rect 44368 27226 44424 27228
rect 44448 27226 44504 27228
rect 44528 27226 44584 27228
rect 44288 27174 44334 27226
rect 44334 27174 44344 27226
rect 44368 27174 44398 27226
rect 44398 27174 44410 27226
rect 44410 27174 44424 27226
rect 44448 27174 44462 27226
rect 44462 27174 44474 27226
rect 44474 27174 44504 27226
rect 44528 27174 44538 27226
rect 44538 27174 44584 27226
rect 44288 27172 44344 27174
rect 44368 27172 44424 27174
rect 44448 27172 44504 27174
rect 44528 27172 44584 27174
rect 8178 26682 8234 26684
rect 8258 26682 8314 26684
rect 8338 26682 8394 26684
rect 8418 26682 8474 26684
rect 8178 26630 8224 26682
rect 8224 26630 8234 26682
rect 8258 26630 8288 26682
rect 8288 26630 8300 26682
rect 8300 26630 8314 26682
rect 8338 26630 8352 26682
rect 8352 26630 8364 26682
rect 8364 26630 8394 26682
rect 8418 26630 8428 26682
rect 8428 26630 8474 26682
rect 8178 26628 8234 26630
rect 8258 26628 8314 26630
rect 8338 26628 8394 26630
rect 8418 26628 8474 26630
rect 15400 26138 15456 26140
rect 15480 26138 15536 26140
rect 15560 26138 15616 26140
rect 15640 26138 15696 26140
rect 15400 26086 15446 26138
rect 15446 26086 15456 26138
rect 15480 26086 15510 26138
rect 15510 26086 15522 26138
rect 15522 26086 15536 26138
rect 15560 26086 15574 26138
rect 15574 26086 15586 26138
rect 15586 26086 15616 26138
rect 15640 26086 15650 26138
rect 15650 26086 15696 26138
rect 15400 26084 15456 26086
rect 15480 26084 15536 26086
rect 15560 26084 15616 26086
rect 15640 26084 15696 26086
rect 8178 25594 8234 25596
rect 8258 25594 8314 25596
rect 8338 25594 8394 25596
rect 8418 25594 8474 25596
rect 8178 25542 8224 25594
rect 8224 25542 8234 25594
rect 8258 25542 8288 25594
rect 8288 25542 8300 25594
rect 8300 25542 8314 25594
rect 8338 25542 8352 25594
rect 8352 25542 8364 25594
rect 8364 25542 8394 25594
rect 8418 25542 8428 25594
rect 8428 25542 8474 25594
rect 8178 25540 8234 25542
rect 8258 25540 8314 25542
rect 8338 25540 8394 25542
rect 8418 25540 8474 25542
rect 8178 24506 8234 24508
rect 8258 24506 8314 24508
rect 8338 24506 8394 24508
rect 8418 24506 8474 24508
rect 8178 24454 8224 24506
rect 8224 24454 8234 24506
rect 8258 24454 8288 24506
rect 8288 24454 8300 24506
rect 8300 24454 8314 24506
rect 8338 24454 8352 24506
rect 8352 24454 8364 24506
rect 8364 24454 8394 24506
rect 8418 24454 8428 24506
rect 8428 24454 8474 24506
rect 8178 24452 8234 24454
rect 8258 24452 8314 24454
rect 8338 24452 8394 24454
rect 8418 24452 8474 24454
rect 2502 11192 2558 11248
rect 2778 11092 2780 11112
rect 2780 11092 2832 11112
rect 2832 11092 2834 11112
rect 2778 11056 2834 11092
rect 938 3440 994 3496
rect 1582 4004 1638 4040
rect 1582 3984 1584 4004
rect 1584 3984 1636 4004
rect 1636 3984 1638 4004
rect 2226 2932 2228 2952
rect 2228 2932 2280 2952
rect 2280 2932 2282 2952
rect 2226 2896 2282 2932
rect 4434 11228 4436 11248
rect 4436 11228 4488 11248
rect 4488 11228 4490 11248
rect 4434 11192 4490 11228
rect 4434 11092 4436 11112
rect 4436 11092 4488 11112
rect 4488 11092 4490 11112
rect 4434 11056 4490 11092
rect 4802 3984 4858 4040
rect 8178 23418 8234 23420
rect 8258 23418 8314 23420
rect 8338 23418 8394 23420
rect 8418 23418 8474 23420
rect 8178 23366 8224 23418
rect 8224 23366 8234 23418
rect 8258 23366 8288 23418
rect 8288 23366 8300 23418
rect 8300 23366 8314 23418
rect 8338 23366 8352 23418
rect 8352 23366 8364 23418
rect 8364 23366 8394 23418
rect 8418 23366 8428 23418
rect 8428 23366 8474 23418
rect 8178 23364 8234 23366
rect 8258 23364 8314 23366
rect 8338 23364 8394 23366
rect 8418 23364 8474 23366
rect 8178 22330 8234 22332
rect 8258 22330 8314 22332
rect 8338 22330 8394 22332
rect 8418 22330 8474 22332
rect 8178 22278 8224 22330
rect 8224 22278 8234 22330
rect 8258 22278 8288 22330
rect 8288 22278 8300 22330
rect 8300 22278 8314 22330
rect 8338 22278 8352 22330
rect 8352 22278 8364 22330
rect 8364 22278 8394 22330
rect 8418 22278 8428 22330
rect 8428 22278 8474 22330
rect 8178 22276 8234 22278
rect 8258 22276 8314 22278
rect 8338 22276 8394 22278
rect 8418 22276 8474 22278
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 10046 19352 10102 19408
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 9770 16652 9826 16688
rect 9770 16632 9772 16652
rect 9772 16632 9824 16652
rect 9824 16632 9826 16652
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 9678 9424 9734 9480
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 7194 4140 7250 4176
rect 7194 4120 7196 4140
rect 7196 4120 7248 4140
rect 7248 4120 7250 4140
rect 6366 2932 6368 2952
rect 6368 2932 6420 2952
rect 6420 2932 6422 2952
rect 6366 2896 6422 2932
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 9218 4140 9274 4176
rect 9218 4120 9220 4140
rect 9220 4120 9272 4140
rect 9272 4120 9274 4140
rect 8114 2932 8116 2952
rect 8116 2932 8168 2952
rect 8168 2932 8170 2952
rect 8114 2896 8170 2932
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 9954 6316 10010 6352
rect 9954 6296 9956 6316
rect 9956 6296 10008 6316
rect 10008 6296 10010 6316
rect 10598 6724 10654 6760
rect 10598 6704 10600 6724
rect 10600 6704 10652 6724
rect 10652 6704 10654 6724
rect 10506 3984 10562 4040
rect 11058 11056 11114 11112
rect 11702 6840 11758 6896
rect 11334 6724 11390 6760
rect 11334 6704 11336 6724
rect 11336 6704 11388 6724
rect 11388 6704 11390 6724
rect 15400 25050 15456 25052
rect 15480 25050 15536 25052
rect 15560 25050 15616 25052
rect 15640 25050 15696 25052
rect 15400 24998 15446 25050
rect 15446 24998 15456 25050
rect 15480 24998 15510 25050
rect 15510 24998 15522 25050
rect 15522 24998 15536 25050
rect 15560 24998 15574 25050
rect 15574 24998 15586 25050
rect 15586 24998 15616 25050
rect 15640 24998 15650 25050
rect 15650 24998 15696 25050
rect 15400 24996 15456 24998
rect 15480 24996 15536 24998
rect 15560 24996 15616 24998
rect 15640 24996 15696 24998
rect 15400 23962 15456 23964
rect 15480 23962 15536 23964
rect 15560 23962 15616 23964
rect 15640 23962 15696 23964
rect 15400 23910 15446 23962
rect 15446 23910 15456 23962
rect 15480 23910 15510 23962
rect 15510 23910 15522 23962
rect 15522 23910 15536 23962
rect 15560 23910 15574 23962
rect 15574 23910 15586 23962
rect 15586 23910 15616 23962
rect 15640 23910 15650 23962
rect 15650 23910 15696 23962
rect 15400 23908 15456 23910
rect 15480 23908 15536 23910
rect 15560 23908 15616 23910
rect 15640 23908 15696 23910
rect 15400 22874 15456 22876
rect 15480 22874 15536 22876
rect 15560 22874 15616 22876
rect 15640 22874 15696 22876
rect 15400 22822 15446 22874
rect 15446 22822 15456 22874
rect 15480 22822 15510 22874
rect 15510 22822 15522 22874
rect 15522 22822 15536 22874
rect 15560 22822 15574 22874
rect 15574 22822 15586 22874
rect 15586 22822 15616 22874
rect 15640 22822 15650 22874
rect 15650 22822 15696 22874
rect 15400 22820 15456 22822
rect 15480 22820 15536 22822
rect 15560 22820 15616 22822
rect 15640 22820 15696 22822
rect 15400 21786 15456 21788
rect 15480 21786 15536 21788
rect 15560 21786 15616 21788
rect 15640 21786 15696 21788
rect 15400 21734 15446 21786
rect 15446 21734 15456 21786
rect 15480 21734 15510 21786
rect 15510 21734 15522 21786
rect 15522 21734 15536 21786
rect 15560 21734 15574 21786
rect 15574 21734 15586 21786
rect 15586 21734 15616 21786
rect 15640 21734 15650 21786
rect 15650 21734 15696 21786
rect 15400 21732 15456 21734
rect 15480 21732 15536 21734
rect 15560 21732 15616 21734
rect 15640 21732 15696 21734
rect 15400 20698 15456 20700
rect 15480 20698 15536 20700
rect 15560 20698 15616 20700
rect 15640 20698 15696 20700
rect 15400 20646 15446 20698
rect 15446 20646 15456 20698
rect 15480 20646 15510 20698
rect 15510 20646 15522 20698
rect 15522 20646 15536 20698
rect 15560 20646 15574 20698
rect 15574 20646 15586 20698
rect 15586 20646 15616 20698
rect 15640 20646 15650 20698
rect 15650 20646 15696 20698
rect 15400 20644 15456 20646
rect 15480 20644 15536 20646
rect 15560 20644 15616 20646
rect 15640 20644 15696 20646
rect 12898 6160 12954 6216
rect 15400 19610 15456 19612
rect 15480 19610 15536 19612
rect 15560 19610 15616 19612
rect 15640 19610 15696 19612
rect 15400 19558 15446 19610
rect 15446 19558 15456 19610
rect 15480 19558 15510 19610
rect 15510 19558 15522 19610
rect 15522 19558 15536 19610
rect 15560 19558 15574 19610
rect 15574 19558 15586 19610
rect 15586 19558 15616 19610
rect 15640 19558 15650 19610
rect 15650 19558 15696 19610
rect 15400 19556 15456 19558
rect 15480 19556 15536 19558
rect 15560 19556 15616 19558
rect 15640 19556 15696 19558
rect 15400 18522 15456 18524
rect 15480 18522 15536 18524
rect 15560 18522 15616 18524
rect 15640 18522 15696 18524
rect 15400 18470 15446 18522
rect 15446 18470 15456 18522
rect 15480 18470 15510 18522
rect 15510 18470 15522 18522
rect 15522 18470 15536 18522
rect 15560 18470 15574 18522
rect 15574 18470 15586 18522
rect 15586 18470 15616 18522
rect 15640 18470 15650 18522
rect 15650 18470 15696 18522
rect 15400 18468 15456 18470
rect 15480 18468 15536 18470
rect 15560 18468 15616 18470
rect 15640 18468 15696 18470
rect 15400 17434 15456 17436
rect 15480 17434 15536 17436
rect 15560 17434 15616 17436
rect 15640 17434 15696 17436
rect 15400 17382 15446 17434
rect 15446 17382 15456 17434
rect 15480 17382 15510 17434
rect 15510 17382 15522 17434
rect 15522 17382 15536 17434
rect 15560 17382 15574 17434
rect 15574 17382 15586 17434
rect 15586 17382 15616 17434
rect 15640 17382 15650 17434
rect 15650 17382 15696 17434
rect 15400 17380 15456 17382
rect 15480 17380 15536 17382
rect 15560 17380 15616 17382
rect 15640 17380 15696 17382
rect 15400 16346 15456 16348
rect 15480 16346 15536 16348
rect 15560 16346 15616 16348
rect 15640 16346 15696 16348
rect 15400 16294 15446 16346
rect 15446 16294 15456 16346
rect 15480 16294 15510 16346
rect 15510 16294 15522 16346
rect 15522 16294 15536 16346
rect 15560 16294 15574 16346
rect 15574 16294 15586 16346
rect 15586 16294 15616 16346
rect 15640 16294 15650 16346
rect 15650 16294 15696 16346
rect 15400 16292 15456 16294
rect 15480 16292 15536 16294
rect 15560 16292 15616 16294
rect 15640 16292 15696 16294
rect 15400 15258 15456 15260
rect 15480 15258 15536 15260
rect 15560 15258 15616 15260
rect 15640 15258 15696 15260
rect 15400 15206 15446 15258
rect 15446 15206 15456 15258
rect 15480 15206 15510 15258
rect 15510 15206 15522 15258
rect 15522 15206 15536 15258
rect 15560 15206 15574 15258
rect 15574 15206 15586 15258
rect 15586 15206 15616 15258
rect 15640 15206 15650 15258
rect 15650 15206 15696 15258
rect 15400 15204 15456 15206
rect 15480 15204 15536 15206
rect 15560 15204 15616 15206
rect 15640 15204 15696 15206
rect 15400 14170 15456 14172
rect 15480 14170 15536 14172
rect 15560 14170 15616 14172
rect 15640 14170 15696 14172
rect 15400 14118 15446 14170
rect 15446 14118 15456 14170
rect 15480 14118 15510 14170
rect 15510 14118 15522 14170
rect 15522 14118 15536 14170
rect 15560 14118 15574 14170
rect 15574 14118 15586 14170
rect 15586 14118 15616 14170
rect 15640 14118 15650 14170
rect 15650 14118 15696 14170
rect 15400 14116 15456 14118
rect 15480 14116 15536 14118
rect 15560 14116 15616 14118
rect 15640 14116 15696 14118
rect 15400 13082 15456 13084
rect 15480 13082 15536 13084
rect 15560 13082 15616 13084
rect 15640 13082 15696 13084
rect 15400 13030 15446 13082
rect 15446 13030 15456 13082
rect 15480 13030 15510 13082
rect 15510 13030 15522 13082
rect 15522 13030 15536 13082
rect 15560 13030 15574 13082
rect 15574 13030 15586 13082
rect 15586 13030 15616 13082
rect 15640 13030 15650 13082
rect 15650 13030 15696 13082
rect 15400 13028 15456 13030
rect 15480 13028 15536 13030
rect 15560 13028 15616 13030
rect 15640 13028 15696 13030
rect 15400 11994 15456 11996
rect 15480 11994 15536 11996
rect 15560 11994 15616 11996
rect 15640 11994 15696 11996
rect 15400 11942 15446 11994
rect 15446 11942 15456 11994
rect 15480 11942 15510 11994
rect 15510 11942 15522 11994
rect 15522 11942 15536 11994
rect 15560 11942 15574 11994
rect 15574 11942 15586 11994
rect 15586 11942 15616 11994
rect 15640 11942 15650 11994
rect 15650 11942 15696 11994
rect 15400 11940 15456 11942
rect 15480 11940 15536 11942
rect 15560 11940 15616 11942
rect 15640 11940 15696 11942
rect 15400 10906 15456 10908
rect 15480 10906 15536 10908
rect 15560 10906 15616 10908
rect 15640 10906 15696 10908
rect 15400 10854 15446 10906
rect 15446 10854 15456 10906
rect 15480 10854 15510 10906
rect 15510 10854 15522 10906
rect 15522 10854 15536 10906
rect 15560 10854 15574 10906
rect 15574 10854 15586 10906
rect 15586 10854 15616 10906
rect 15640 10854 15650 10906
rect 15650 10854 15696 10906
rect 15400 10852 15456 10854
rect 15480 10852 15536 10854
rect 15560 10852 15616 10854
rect 15640 10852 15696 10854
rect 22622 26682 22678 26684
rect 22702 26682 22758 26684
rect 22782 26682 22838 26684
rect 22862 26682 22918 26684
rect 22622 26630 22668 26682
rect 22668 26630 22678 26682
rect 22702 26630 22732 26682
rect 22732 26630 22744 26682
rect 22744 26630 22758 26682
rect 22782 26630 22796 26682
rect 22796 26630 22808 26682
rect 22808 26630 22838 26682
rect 22862 26630 22872 26682
rect 22872 26630 22918 26682
rect 22622 26628 22678 26630
rect 22702 26628 22758 26630
rect 22782 26628 22838 26630
rect 22862 26628 22918 26630
rect 15400 9818 15456 9820
rect 15480 9818 15536 9820
rect 15560 9818 15616 9820
rect 15640 9818 15696 9820
rect 15400 9766 15446 9818
rect 15446 9766 15456 9818
rect 15480 9766 15510 9818
rect 15510 9766 15522 9818
rect 15522 9766 15536 9818
rect 15560 9766 15574 9818
rect 15574 9766 15586 9818
rect 15586 9766 15616 9818
rect 15640 9766 15650 9818
rect 15650 9766 15696 9818
rect 15400 9764 15456 9766
rect 15480 9764 15536 9766
rect 15560 9764 15616 9766
rect 15640 9764 15696 9766
rect 15400 8730 15456 8732
rect 15480 8730 15536 8732
rect 15560 8730 15616 8732
rect 15640 8730 15696 8732
rect 15400 8678 15446 8730
rect 15446 8678 15456 8730
rect 15480 8678 15510 8730
rect 15510 8678 15522 8730
rect 15522 8678 15536 8730
rect 15560 8678 15574 8730
rect 15574 8678 15586 8730
rect 15586 8678 15616 8730
rect 15640 8678 15650 8730
rect 15650 8678 15696 8730
rect 15400 8676 15456 8678
rect 15480 8676 15536 8678
rect 15560 8676 15616 8678
rect 15640 8676 15696 8678
rect 15400 7642 15456 7644
rect 15480 7642 15536 7644
rect 15560 7642 15616 7644
rect 15640 7642 15696 7644
rect 15400 7590 15446 7642
rect 15446 7590 15456 7642
rect 15480 7590 15510 7642
rect 15510 7590 15522 7642
rect 15522 7590 15536 7642
rect 15560 7590 15574 7642
rect 15574 7590 15586 7642
rect 15586 7590 15616 7642
rect 15640 7590 15650 7642
rect 15650 7590 15696 7642
rect 15400 7588 15456 7590
rect 15480 7588 15536 7590
rect 15560 7588 15616 7590
rect 15640 7588 15696 7590
rect 15400 6554 15456 6556
rect 15480 6554 15536 6556
rect 15560 6554 15616 6556
rect 15640 6554 15696 6556
rect 15400 6502 15446 6554
rect 15446 6502 15456 6554
rect 15480 6502 15510 6554
rect 15510 6502 15522 6554
rect 15522 6502 15536 6554
rect 15560 6502 15574 6554
rect 15574 6502 15586 6554
rect 15586 6502 15616 6554
rect 15640 6502 15650 6554
rect 15650 6502 15696 6554
rect 15400 6500 15456 6502
rect 15480 6500 15536 6502
rect 15560 6500 15616 6502
rect 15640 6500 15696 6502
rect 15400 5466 15456 5468
rect 15480 5466 15536 5468
rect 15560 5466 15616 5468
rect 15640 5466 15696 5468
rect 15400 5414 15446 5466
rect 15446 5414 15456 5466
rect 15480 5414 15510 5466
rect 15510 5414 15522 5466
rect 15522 5414 15536 5466
rect 15560 5414 15574 5466
rect 15574 5414 15586 5466
rect 15586 5414 15616 5466
rect 15640 5414 15650 5466
rect 15650 5414 15696 5466
rect 15400 5412 15456 5414
rect 15480 5412 15536 5414
rect 15560 5412 15616 5414
rect 15640 5412 15696 5414
rect 15400 4378 15456 4380
rect 15480 4378 15536 4380
rect 15560 4378 15616 4380
rect 15640 4378 15696 4380
rect 15400 4326 15446 4378
rect 15446 4326 15456 4378
rect 15480 4326 15510 4378
rect 15510 4326 15522 4378
rect 15522 4326 15536 4378
rect 15560 4326 15574 4378
rect 15574 4326 15586 4378
rect 15586 4326 15616 4378
rect 15640 4326 15650 4378
rect 15650 4326 15696 4378
rect 15400 4324 15456 4326
rect 15480 4324 15536 4326
rect 15560 4324 15616 4326
rect 15640 4324 15696 4326
rect 15400 3290 15456 3292
rect 15480 3290 15536 3292
rect 15560 3290 15616 3292
rect 15640 3290 15696 3292
rect 15400 3238 15446 3290
rect 15446 3238 15456 3290
rect 15480 3238 15510 3290
rect 15510 3238 15522 3290
rect 15522 3238 15536 3290
rect 15560 3238 15574 3290
rect 15574 3238 15586 3290
rect 15586 3238 15616 3290
rect 15640 3238 15650 3290
rect 15650 3238 15696 3290
rect 15400 3236 15456 3238
rect 15480 3236 15536 3238
rect 15560 3236 15616 3238
rect 15640 3236 15696 3238
rect 22622 25594 22678 25596
rect 22702 25594 22758 25596
rect 22782 25594 22838 25596
rect 22862 25594 22918 25596
rect 22622 25542 22668 25594
rect 22668 25542 22678 25594
rect 22702 25542 22732 25594
rect 22732 25542 22744 25594
rect 22744 25542 22758 25594
rect 22782 25542 22796 25594
rect 22796 25542 22808 25594
rect 22808 25542 22838 25594
rect 22862 25542 22872 25594
rect 22872 25542 22918 25594
rect 22622 25540 22678 25542
rect 22702 25540 22758 25542
rect 22782 25540 22838 25542
rect 22862 25540 22918 25542
rect 22622 24506 22678 24508
rect 22702 24506 22758 24508
rect 22782 24506 22838 24508
rect 22862 24506 22918 24508
rect 22622 24454 22668 24506
rect 22668 24454 22678 24506
rect 22702 24454 22732 24506
rect 22732 24454 22744 24506
rect 22744 24454 22758 24506
rect 22782 24454 22796 24506
rect 22796 24454 22808 24506
rect 22808 24454 22838 24506
rect 22862 24454 22872 24506
rect 22872 24454 22918 24506
rect 22622 24452 22678 24454
rect 22702 24452 22758 24454
rect 22782 24452 22838 24454
rect 22862 24452 22918 24454
rect 22622 23418 22678 23420
rect 22702 23418 22758 23420
rect 22782 23418 22838 23420
rect 22862 23418 22918 23420
rect 22622 23366 22668 23418
rect 22668 23366 22678 23418
rect 22702 23366 22732 23418
rect 22732 23366 22744 23418
rect 22744 23366 22758 23418
rect 22782 23366 22796 23418
rect 22796 23366 22808 23418
rect 22808 23366 22838 23418
rect 22862 23366 22872 23418
rect 22872 23366 22918 23418
rect 22622 23364 22678 23366
rect 22702 23364 22758 23366
rect 22782 23364 22838 23366
rect 22862 23364 22918 23366
rect 16946 7812 17002 7848
rect 16946 7792 16948 7812
rect 16948 7792 17000 7812
rect 17000 7792 17002 7812
rect 15400 2202 15456 2204
rect 15480 2202 15536 2204
rect 15560 2202 15616 2204
rect 15640 2202 15696 2204
rect 15400 2150 15446 2202
rect 15446 2150 15456 2202
rect 15480 2150 15510 2202
rect 15510 2150 15522 2202
rect 15522 2150 15536 2202
rect 15560 2150 15574 2202
rect 15574 2150 15586 2202
rect 15586 2150 15616 2202
rect 15640 2150 15650 2202
rect 15650 2150 15696 2202
rect 15400 2148 15456 2150
rect 15480 2148 15536 2150
rect 15560 2148 15616 2150
rect 15640 2148 15696 2150
rect 16762 3984 16818 4040
rect 17866 4256 17922 4312
rect 18234 3848 18290 3904
rect 18510 3984 18566 4040
rect 18878 4256 18934 4312
rect 19246 3848 19302 3904
rect 22622 22330 22678 22332
rect 22702 22330 22758 22332
rect 22782 22330 22838 22332
rect 22862 22330 22918 22332
rect 22622 22278 22668 22330
rect 22668 22278 22678 22330
rect 22702 22278 22732 22330
rect 22732 22278 22744 22330
rect 22744 22278 22758 22330
rect 22782 22278 22796 22330
rect 22796 22278 22808 22330
rect 22808 22278 22838 22330
rect 22862 22278 22872 22330
rect 22872 22278 22918 22330
rect 22622 22276 22678 22278
rect 22702 22276 22758 22278
rect 22782 22276 22838 22278
rect 22862 22276 22918 22278
rect 22622 21242 22678 21244
rect 22702 21242 22758 21244
rect 22782 21242 22838 21244
rect 22862 21242 22918 21244
rect 22622 21190 22668 21242
rect 22668 21190 22678 21242
rect 22702 21190 22732 21242
rect 22732 21190 22744 21242
rect 22744 21190 22758 21242
rect 22782 21190 22796 21242
rect 22796 21190 22808 21242
rect 22808 21190 22838 21242
rect 22862 21190 22872 21242
rect 22872 21190 22918 21242
rect 22622 21188 22678 21190
rect 22702 21188 22758 21190
rect 22782 21188 22838 21190
rect 22862 21188 22918 21190
rect 22622 20154 22678 20156
rect 22702 20154 22758 20156
rect 22782 20154 22838 20156
rect 22862 20154 22918 20156
rect 22622 20102 22668 20154
rect 22668 20102 22678 20154
rect 22702 20102 22732 20154
rect 22732 20102 22744 20154
rect 22744 20102 22758 20154
rect 22782 20102 22796 20154
rect 22796 20102 22808 20154
rect 22808 20102 22838 20154
rect 22862 20102 22872 20154
rect 22872 20102 22918 20154
rect 22622 20100 22678 20102
rect 22702 20100 22758 20102
rect 22782 20100 22838 20102
rect 22862 20100 22918 20102
rect 22622 19066 22678 19068
rect 22702 19066 22758 19068
rect 22782 19066 22838 19068
rect 22862 19066 22918 19068
rect 22622 19014 22668 19066
rect 22668 19014 22678 19066
rect 22702 19014 22732 19066
rect 22732 19014 22744 19066
rect 22744 19014 22758 19066
rect 22782 19014 22796 19066
rect 22796 19014 22808 19066
rect 22808 19014 22838 19066
rect 22862 19014 22872 19066
rect 22872 19014 22918 19066
rect 22622 19012 22678 19014
rect 22702 19012 22758 19014
rect 22782 19012 22838 19014
rect 22862 19012 22918 19014
rect 22622 17978 22678 17980
rect 22702 17978 22758 17980
rect 22782 17978 22838 17980
rect 22862 17978 22918 17980
rect 22622 17926 22668 17978
rect 22668 17926 22678 17978
rect 22702 17926 22732 17978
rect 22732 17926 22744 17978
rect 22744 17926 22758 17978
rect 22782 17926 22796 17978
rect 22796 17926 22808 17978
rect 22808 17926 22838 17978
rect 22862 17926 22872 17978
rect 22872 17926 22918 17978
rect 22622 17924 22678 17926
rect 22702 17924 22758 17926
rect 22782 17924 22838 17926
rect 22862 17924 22918 17926
rect 22622 16890 22678 16892
rect 22702 16890 22758 16892
rect 22782 16890 22838 16892
rect 22862 16890 22918 16892
rect 22622 16838 22668 16890
rect 22668 16838 22678 16890
rect 22702 16838 22732 16890
rect 22732 16838 22744 16890
rect 22744 16838 22758 16890
rect 22782 16838 22796 16890
rect 22796 16838 22808 16890
rect 22808 16838 22838 16890
rect 22862 16838 22872 16890
rect 22872 16838 22918 16890
rect 22622 16836 22678 16838
rect 22702 16836 22758 16838
rect 22782 16836 22838 16838
rect 22862 16836 22918 16838
rect 22622 15802 22678 15804
rect 22702 15802 22758 15804
rect 22782 15802 22838 15804
rect 22862 15802 22918 15804
rect 22622 15750 22668 15802
rect 22668 15750 22678 15802
rect 22702 15750 22732 15802
rect 22732 15750 22744 15802
rect 22744 15750 22758 15802
rect 22782 15750 22796 15802
rect 22796 15750 22808 15802
rect 22808 15750 22838 15802
rect 22862 15750 22872 15802
rect 22872 15750 22918 15802
rect 22622 15748 22678 15750
rect 22702 15748 22758 15750
rect 22782 15748 22838 15750
rect 22862 15748 22918 15750
rect 22622 14714 22678 14716
rect 22702 14714 22758 14716
rect 22782 14714 22838 14716
rect 22862 14714 22918 14716
rect 22622 14662 22668 14714
rect 22668 14662 22678 14714
rect 22702 14662 22732 14714
rect 22732 14662 22744 14714
rect 22744 14662 22758 14714
rect 22782 14662 22796 14714
rect 22796 14662 22808 14714
rect 22808 14662 22838 14714
rect 22862 14662 22872 14714
rect 22872 14662 22918 14714
rect 22622 14660 22678 14662
rect 22702 14660 22758 14662
rect 22782 14660 22838 14662
rect 22862 14660 22918 14662
rect 22622 13626 22678 13628
rect 22702 13626 22758 13628
rect 22782 13626 22838 13628
rect 22862 13626 22918 13628
rect 22622 13574 22668 13626
rect 22668 13574 22678 13626
rect 22702 13574 22732 13626
rect 22732 13574 22744 13626
rect 22744 13574 22758 13626
rect 22782 13574 22796 13626
rect 22796 13574 22808 13626
rect 22808 13574 22838 13626
rect 22862 13574 22872 13626
rect 22872 13574 22918 13626
rect 22622 13572 22678 13574
rect 22702 13572 22758 13574
rect 22782 13572 22838 13574
rect 22862 13572 22918 13574
rect 22622 12538 22678 12540
rect 22702 12538 22758 12540
rect 22782 12538 22838 12540
rect 22862 12538 22918 12540
rect 22622 12486 22668 12538
rect 22668 12486 22678 12538
rect 22702 12486 22732 12538
rect 22732 12486 22744 12538
rect 22744 12486 22758 12538
rect 22782 12486 22796 12538
rect 22796 12486 22808 12538
rect 22808 12486 22838 12538
rect 22862 12486 22872 12538
rect 22872 12486 22918 12538
rect 22622 12484 22678 12486
rect 22702 12484 22758 12486
rect 22782 12484 22838 12486
rect 22862 12484 22918 12486
rect 23478 12144 23534 12200
rect 22622 11450 22678 11452
rect 22702 11450 22758 11452
rect 22782 11450 22838 11452
rect 22862 11450 22918 11452
rect 22622 11398 22668 11450
rect 22668 11398 22678 11450
rect 22702 11398 22732 11450
rect 22732 11398 22744 11450
rect 22744 11398 22758 11450
rect 22782 11398 22796 11450
rect 22796 11398 22808 11450
rect 22808 11398 22838 11450
rect 22862 11398 22872 11450
rect 22872 11398 22918 11450
rect 22622 11396 22678 11398
rect 22702 11396 22758 11398
rect 22782 11396 22838 11398
rect 22862 11396 22918 11398
rect 22006 10104 22062 10160
rect 22622 10362 22678 10364
rect 22702 10362 22758 10364
rect 22782 10362 22838 10364
rect 22862 10362 22918 10364
rect 22622 10310 22668 10362
rect 22668 10310 22678 10362
rect 22702 10310 22732 10362
rect 22732 10310 22744 10362
rect 22744 10310 22758 10362
rect 22782 10310 22796 10362
rect 22796 10310 22808 10362
rect 22808 10310 22838 10362
rect 22862 10310 22872 10362
rect 22872 10310 22918 10362
rect 22622 10308 22678 10310
rect 22702 10308 22758 10310
rect 22782 10308 22838 10310
rect 22862 10308 22918 10310
rect 22558 10104 22614 10160
rect 22622 9274 22678 9276
rect 22702 9274 22758 9276
rect 22782 9274 22838 9276
rect 22862 9274 22918 9276
rect 22622 9222 22668 9274
rect 22668 9222 22678 9274
rect 22702 9222 22732 9274
rect 22732 9222 22744 9274
rect 22744 9222 22758 9274
rect 22782 9222 22796 9274
rect 22796 9222 22808 9274
rect 22808 9222 22838 9274
rect 22862 9222 22872 9274
rect 22872 9222 22918 9274
rect 22622 9220 22678 9222
rect 22702 9220 22758 9222
rect 22782 9220 22838 9222
rect 22862 9220 22918 9222
rect 22006 7692 22008 7712
rect 22008 7692 22060 7712
rect 22060 7692 22062 7712
rect 22006 7656 22062 7692
rect 22622 8186 22678 8188
rect 22702 8186 22758 8188
rect 22782 8186 22838 8188
rect 22862 8186 22918 8188
rect 22622 8134 22668 8186
rect 22668 8134 22678 8186
rect 22702 8134 22732 8186
rect 22732 8134 22744 8186
rect 22744 8134 22758 8186
rect 22782 8134 22796 8186
rect 22796 8134 22808 8186
rect 22808 8134 22838 8186
rect 22862 8134 22872 8186
rect 22872 8134 22918 8186
rect 22622 8132 22678 8134
rect 22702 8132 22758 8134
rect 22782 8132 22838 8134
rect 22862 8132 22918 8134
rect 22622 7098 22678 7100
rect 22702 7098 22758 7100
rect 22782 7098 22838 7100
rect 22862 7098 22918 7100
rect 22622 7046 22668 7098
rect 22668 7046 22678 7098
rect 22702 7046 22732 7098
rect 22732 7046 22744 7098
rect 22744 7046 22758 7098
rect 22782 7046 22796 7098
rect 22796 7046 22808 7098
rect 22808 7046 22838 7098
rect 22862 7046 22872 7098
rect 22872 7046 22918 7098
rect 22622 7044 22678 7046
rect 22702 7044 22758 7046
rect 22782 7044 22838 7046
rect 22862 7044 22918 7046
rect 22006 5072 22062 5128
rect 21638 3304 21694 3360
rect 21454 3052 21510 3088
rect 21454 3032 21456 3052
rect 21456 3032 21508 3052
rect 21508 3032 21510 3052
rect 22622 6010 22678 6012
rect 22702 6010 22758 6012
rect 22782 6010 22838 6012
rect 22862 6010 22918 6012
rect 22622 5958 22668 6010
rect 22668 5958 22678 6010
rect 22702 5958 22732 6010
rect 22732 5958 22744 6010
rect 22744 5958 22758 6010
rect 22782 5958 22796 6010
rect 22796 5958 22808 6010
rect 22808 5958 22838 6010
rect 22862 5958 22872 6010
rect 22872 5958 22918 6010
rect 22622 5956 22678 5958
rect 22702 5956 22758 5958
rect 22782 5956 22838 5958
rect 22862 5956 22918 5958
rect 22622 4922 22678 4924
rect 22702 4922 22758 4924
rect 22782 4922 22838 4924
rect 22862 4922 22918 4924
rect 22622 4870 22668 4922
rect 22668 4870 22678 4922
rect 22702 4870 22732 4922
rect 22732 4870 22744 4922
rect 22744 4870 22758 4922
rect 22782 4870 22796 4922
rect 22796 4870 22808 4922
rect 22808 4870 22838 4922
rect 22862 4870 22872 4922
rect 22872 4870 22918 4922
rect 22622 4868 22678 4870
rect 22702 4868 22758 4870
rect 22782 4868 22838 4870
rect 22862 4868 22918 4870
rect 22622 3834 22678 3836
rect 22702 3834 22758 3836
rect 22782 3834 22838 3836
rect 22862 3834 22918 3836
rect 22622 3782 22668 3834
rect 22668 3782 22678 3834
rect 22702 3782 22732 3834
rect 22732 3782 22744 3834
rect 22744 3782 22758 3834
rect 22782 3782 22796 3834
rect 22796 3782 22808 3834
rect 22808 3782 22838 3834
rect 22862 3782 22872 3834
rect 22872 3782 22918 3834
rect 22622 3780 22678 3782
rect 22702 3780 22758 3782
rect 22782 3780 22838 3782
rect 22862 3780 22918 3782
rect 22098 3304 22154 3360
rect 22742 3068 22744 3088
rect 22744 3068 22796 3088
rect 22796 3068 22798 3088
rect 22742 3032 22798 3068
rect 22622 2746 22678 2748
rect 22702 2746 22758 2748
rect 22782 2746 22838 2748
rect 22862 2746 22918 2748
rect 22622 2694 22668 2746
rect 22668 2694 22678 2746
rect 22702 2694 22732 2746
rect 22732 2694 22744 2746
rect 22744 2694 22758 2746
rect 22782 2694 22796 2746
rect 22796 2694 22808 2746
rect 22808 2694 22838 2746
rect 22862 2694 22872 2746
rect 22872 2694 22918 2746
rect 22622 2692 22678 2694
rect 22702 2692 22758 2694
rect 22782 2692 22838 2694
rect 22862 2692 22918 2694
rect 29844 26138 29900 26140
rect 29924 26138 29980 26140
rect 30004 26138 30060 26140
rect 30084 26138 30140 26140
rect 29844 26086 29890 26138
rect 29890 26086 29900 26138
rect 29924 26086 29954 26138
rect 29954 26086 29966 26138
rect 29966 26086 29980 26138
rect 30004 26086 30018 26138
rect 30018 26086 30030 26138
rect 30030 26086 30060 26138
rect 30084 26086 30094 26138
rect 30094 26086 30140 26138
rect 29844 26084 29900 26086
rect 29924 26084 29980 26086
rect 30004 26084 30060 26086
rect 30084 26084 30140 26086
rect 29844 25050 29900 25052
rect 29924 25050 29980 25052
rect 30004 25050 30060 25052
rect 30084 25050 30140 25052
rect 29844 24998 29890 25050
rect 29890 24998 29900 25050
rect 29924 24998 29954 25050
rect 29954 24998 29966 25050
rect 29966 24998 29980 25050
rect 30004 24998 30018 25050
rect 30018 24998 30030 25050
rect 30030 24998 30060 25050
rect 30084 24998 30094 25050
rect 30094 24998 30140 25050
rect 29844 24996 29900 24998
rect 29924 24996 29980 24998
rect 30004 24996 30060 24998
rect 30084 24996 30140 24998
rect 37066 26682 37122 26684
rect 37146 26682 37202 26684
rect 37226 26682 37282 26684
rect 37306 26682 37362 26684
rect 37066 26630 37112 26682
rect 37112 26630 37122 26682
rect 37146 26630 37176 26682
rect 37176 26630 37188 26682
rect 37188 26630 37202 26682
rect 37226 26630 37240 26682
rect 37240 26630 37252 26682
rect 37252 26630 37282 26682
rect 37306 26630 37316 26682
rect 37316 26630 37362 26682
rect 37066 26628 37122 26630
rect 37146 26628 37202 26630
rect 37226 26628 37282 26630
rect 37306 26628 37362 26630
rect 29844 23962 29900 23964
rect 29924 23962 29980 23964
rect 30004 23962 30060 23964
rect 30084 23962 30140 23964
rect 29844 23910 29890 23962
rect 29890 23910 29900 23962
rect 29924 23910 29954 23962
rect 29954 23910 29966 23962
rect 29966 23910 29980 23962
rect 30004 23910 30018 23962
rect 30018 23910 30030 23962
rect 30030 23910 30060 23962
rect 30084 23910 30094 23962
rect 30094 23910 30140 23962
rect 29844 23908 29900 23910
rect 29924 23908 29980 23910
rect 30004 23908 30060 23910
rect 30084 23908 30140 23910
rect 29844 22874 29900 22876
rect 29924 22874 29980 22876
rect 30004 22874 30060 22876
rect 30084 22874 30140 22876
rect 29844 22822 29890 22874
rect 29890 22822 29900 22874
rect 29924 22822 29954 22874
rect 29954 22822 29966 22874
rect 29966 22822 29980 22874
rect 30004 22822 30018 22874
rect 30018 22822 30030 22874
rect 30030 22822 30060 22874
rect 30084 22822 30094 22874
rect 30094 22822 30140 22874
rect 29844 22820 29900 22822
rect 29924 22820 29980 22822
rect 30004 22820 30060 22822
rect 30084 22820 30140 22822
rect 29844 21786 29900 21788
rect 29924 21786 29980 21788
rect 30004 21786 30060 21788
rect 30084 21786 30140 21788
rect 29844 21734 29890 21786
rect 29890 21734 29900 21786
rect 29924 21734 29954 21786
rect 29954 21734 29966 21786
rect 29966 21734 29980 21786
rect 30004 21734 30018 21786
rect 30018 21734 30030 21786
rect 30030 21734 30060 21786
rect 30084 21734 30094 21786
rect 30094 21734 30140 21786
rect 29844 21732 29900 21734
rect 29924 21732 29980 21734
rect 30004 21732 30060 21734
rect 30084 21732 30140 21734
rect 37066 25594 37122 25596
rect 37146 25594 37202 25596
rect 37226 25594 37282 25596
rect 37306 25594 37362 25596
rect 37066 25542 37112 25594
rect 37112 25542 37122 25594
rect 37146 25542 37176 25594
rect 37176 25542 37188 25594
rect 37188 25542 37202 25594
rect 37226 25542 37240 25594
rect 37240 25542 37252 25594
rect 37252 25542 37282 25594
rect 37306 25542 37316 25594
rect 37316 25542 37362 25594
rect 37066 25540 37122 25542
rect 37146 25540 37202 25542
rect 37226 25540 37282 25542
rect 37306 25540 37362 25542
rect 37066 24506 37122 24508
rect 37146 24506 37202 24508
rect 37226 24506 37282 24508
rect 37306 24506 37362 24508
rect 37066 24454 37112 24506
rect 37112 24454 37122 24506
rect 37146 24454 37176 24506
rect 37176 24454 37188 24506
rect 37188 24454 37202 24506
rect 37226 24454 37240 24506
rect 37240 24454 37252 24506
rect 37252 24454 37282 24506
rect 37306 24454 37316 24506
rect 37316 24454 37362 24506
rect 37066 24452 37122 24454
rect 37146 24452 37202 24454
rect 37226 24452 37282 24454
rect 37306 24452 37362 24454
rect 26054 7384 26110 7440
rect 26422 7656 26478 7712
rect 26606 2896 26662 2952
rect 27618 12180 27620 12200
rect 27620 12180 27672 12200
rect 27672 12180 27674 12200
rect 27618 12144 27674 12180
rect 29844 20698 29900 20700
rect 29924 20698 29980 20700
rect 30004 20698 30060 20700
rect 30084 20698 30140 20700
rect 29844 20646 29890 20698
rect 29890 20646 29900 20698
rect 29924 20646 29954 20698
rect 29954 20646 29966 20698
rect 29966 20646 29980 20698
rect 30004 20646 30018 20698
rect 30018 20646 30030 20698
rect 30030 20646 30060 20698
rect 30084 20646 30094 20698
rect 30094 20646 30140 20698
rect 29844 20644 29900 20646
rect 29924 20644 29980 20646
rect 30004 20644 30060 20646
rect 30084 20644 30140 20646
rect 29844 19610 29900 19612
rect 29924 19610 29980 19612
rect 30004 19610 30060 19612
rect 30084 19610 30140 19612
rect 29844 19558 29890 19610
rect 29890 19558 29900 19610
rect 29924 19558 29954 19610
rect 29954 19558 29966 19610
rect 29966 19558 29980 19610
rect 30004 19558 30018 19610
rect 30018 19558 30030 19610
rect 30030 19558 30060 19610
rect 30084 19558 30094 19610
rect 30094 19558 30140 19610
rect 29844 19556 29900 19558
rect 29924 19556 29980 19558
rect 30004 19556 30060 19558
rect 30084 19556 30140 19558
rect 29844 18522 29900 18524
rect 29924 18522 29980 18524
rect 30004 18522 30060 18524
rect 30084 18522 30140 18524
rect 29844 18470 29890 18522
rect 29890 18470 29900 18522
rect 29924 18470 29954 18522
rect 29954 18470 29966 18522
rect 29966 18470 29980 18522
rect 30004 18470 30018 18522
rect 30018 18470 30030 18522
rect 30030 18470 30060 18522
rect 30084 18470 30094 18522
rect 30094 18470 30140 18522
rect 29844 18468 29900 18470
rect 29924 18468 29980 18470
rect 30004 18468 30060 18470
rect 30084 18468 30140 18470
rect 29844 17434 29900 17436
rect 29924 17434 29980 17436
rect 30004 17434 30060 17436
rect 30084 17434 30140 17436
rect 29844 17382 29890 17434
rect 29890 17382 29900 17434
rect 29924 17382 29954 17434
rect 29954 17382 29966 17434
rect 29966 17382 29980 17434
rect 30004 17382 30018 17434
rect 30018 17382 30030 17434
rect 30030 17382 30060 17434
rect 30084 17382 30094 17434
rect 30094 17382 30140 17434
rect 29844 17380 29900 17382
rect 29924 17380 29980 17382
rect 30004 17380 30060 17382
rect 30084 17380 30140 17382
rect 27158 4120 27214 4176
rect 26790 3576 26846 3632
rect 29844 16346 29900 16348
rect 29924 16346 29980 16348
rect 30004 16346 30060 16348
rect 30084 16346 30140 16348
rect 29844 16294 29890 16346
rect 29890 16294 29900 16346
rect 29924 16294 29954 16346
rect 29954 16294 29966 16346
rect 29966 16294 29980 16346
rect 30004 16294 30018 16346
rect 30018 16294 30030 16346
rect 30030 16294 30060 16346
rect 30084 16294 30094 16346
rect 30094 16294 30140 16346
rect 29844 16292 29900 16294
rect 29924 16292 29980 16294
rect 30004 16292 30060 16294
rect 30084 16292 30140 16294
rect 29844 15258 29900 15260
rect 29924 15258 29980 15260
rect 30004 15258 30060 15260
rect 30084 15258 30140 15260
rect 29844 15206 29890 15258
rect 29890 15206 29900 15258
rect 29924 15206 29954 15258
rect 29954 15206 29966 15258
rect 29966 15206 29980 15258
rect 30004 15206 30018 15258
rect 30018 15206 30030 15258
rect 30030 15206 30060 15258
rect 30084 15206 30094 15258
rect 30094 15206 30140 15258
rect 29844 15204 29900 15206
rect 29924 15204 29980 15206
rect 30004 15204 30060 15206
rect 30084 15204 30140 15206
rect 29844 14170 29900 14172
rect 29924 14170 29980 14172
rect 30004 14170 30060 14172
rect 30084 14170 30140 14172
rect 29844 14118 29890 14170
rect 29890 14118 29900 14170
rect 29924 14118 29954 14170
rect 29954 14118 29966 14170
rect 29966 14118 29980 14170
rect 30004 14118 30018 14170
rect 30018 14118 30030 14170
rect 30030 14118 30060 14170
rect 30084 14118 30094 14170
rect 30094 14118 30140 14170
rect 29844 14116 29900 14118
rect 29924 14116 29980 14118
rect 30004 14116 30060 14118
rect 30084 14116 30140 14118
rect 28906 5072 28962 5128
rect 29844 13082 29900 13084
rect 29924 13082 29980 13084
rect 30004 13082 30060 13084
rect 30084 13082 30140 13084
rect 29844 13030 29890 13082
rect 29890 13030 29900 13082
rect 29924 13030 29954 13082
rect 29954 13030 29966 13082
rect 29966 13030 29980 13082
rect 30004 13030 30018 13082
rect 30018 13030 30030 13082
rect 30030 13030 30060 13082
rect 30084 13030 30094 13082
rect 30094 13030 30140 13082
rect 29844 13028 29900 13030
rect 29924 13028 29980 13030
rect 30004 13028 30060 13030
rect 30084 13028 30140 13030
rect 29844 11994 29900 11996
rect 29924 11994 29980 11996
rect 30004 11994 30060 11996
rect 30084 11994 30140 11996
rect 29844 11942 29890 11994
rect 29890 11942 29900 11994
rect 29924 11942 29954 11994
rect 29954 11942 29966 11994
rect 29966 11942 29980 11994
rect 30004 11942 30018 11994
rect 30018 11942 30030 11994
rect 30030 11942 30060 11994
rect 30084 11942 30094 11994
rect 30094 11942 30140 11994
rect 29844 11940 29900 11942
rect 29924 11940 29980 11942
rect 30004 11940 30060 11942
rect 30084 11940 30140 11942
rect 29844 10906 29900 10908
rect 29924 10906 29980 10908
rect 30004 10906 30060 10908
rect 30084 10906 30140 10908
rect 29844 10854 29890 10906
rect 29890 10854 29900 10906
rect 29924 10854 29954 10906
rect 29954 10854 29966 10906
rect 29966 10854 29980 10906
rect 30004 10854 30018 10906
rect 30018 10854 30030 10906
rect 30030 10854 30060 10906
rect 30084 10854 30094 10906
rect 30094 10854 30140 10906
rect 29844 10852 29900 10854
rect 29924 10852 29980 10854
rect 30004 10852 30060 10854
rect 30084 10852 30140 10854
rect 29844 9818 29900 9820
rect 29924 9818 29980 9820
rect 30004 9818 30060 9820
rect 30084 9818 30140 9820
rect 29844 9766 29890 9818
rect 29890 9766 29900 9818
rect 29924 9766 29954 9818
rect 29954 9766 29966 9818
rect 29966 9766 29980 9818
rect 30004 9766 30018 9818
rect 30018 9766 30030 9818
rect 30030 9766 30060 9818
rect 30084 9766 30094 9818
rect 30094 9766 30140 9818
rect 29844 9764 29900 9766
rect 29924 9764 29980 9766
rect 30004 9764 30060 9766
rect 30084 9764 30140 9766
rect 29844 8730 29900 8732
rect 29924 8730 29980 8732
rect 30004 8730 30060 8732
rect 30084 8730 30140 8732
rect 29844 8678 29890 8730
rect 29890 8678 29900 8730
rect 29924 8678 29954 8730
rect 29954 8678 29966 8730
rect 29966 8678 29980 8730
rect 30004 8678 30018 8730
rect 30018 8678 30030 8730
rect 30030 8678 30060 8730
rect 30084 8678 30094 8730
rect 30094 8678 30140 8730
rect 29844 8676 29900 8678
rect 29924 8676 29980 8678
rect 30004 8676 30060 8678
rect 30084 8676 30140 8678
rect 29844 7642 29900 7644
rect 29924 7642 29980 7644
rect 30004 7642 30060 7644
rect 30084 7642 30140 7644
rect 29844 7590 29890 7642
rect 29890 7590 29900 7642
rect 29924 7590 29954 7642
rect 29954 7590 29966 7642
rect 29966 7590 29980 7642
rect 30004 7590 30018 7642
rect 30018 7590 30030 7642
rect 30030 7590 30060 7642
rect 30084 7590 30094 7642
rect 30094 7590 30140 7642
rect 29844 7588 29900 7590
rect 29924 7588 29980 7590
rect 30004 7588 30060 7590
rect 30084 7588 30140 7590
rect 29844 6554 29900 6556
rect 29924 6554 29980 6556
rect 30004 6554 30060 6556
rect 30084 6554 30140 6556
rect 29844 6502 29890 6554
rect 29890 6502 29900 6554
rect 29924 6502 29954 6554
rect 29954 6502 29966 6554
rect 29966 6502 29980 6554
rect 30004 6502 30018 6554
rect 30018 6502 30030 6554
rect 30030 6502 30060 6554
rect 30084 6502 30094 6554
rect 30094 6502 30140 6554
rect 29844 6500 29900 6502
rect 29924 6500 29980 6502
rect 30004 6500 30060 6502
rect 30084 6500 30140 6502
rect 29844 5466 29900 5468
rect 29924 5466 29980 5468
rect 30004 5466 30060 5468
rect 30084 5466 30140 5468
rect 29844 5414 29890 5466
rect 29890 5414 29900 5466
rect 29924 5414 29954 5466
rect 29954 5414 29966 5466
rect 29966 5414 29980 5466
rect 30004 5414 30018 5466
rect 30018 5414 30030 5466
rect 30030 5414 30060 5466
rect 30084 5414 30094 5466
rect 30094 5414 30140 5466
rect 29844 5412 29900 5414
rect 29924 5412 29980 5414
rect 30004 5412 30060 5414
rect 30084 5412 30140 5414
rect 29844 4378 29900 4380
rect 29924 4378 29980 4380
rect 30004 4378 30060 4380
rect 30084 4378 30140 4380
rect 29844 4326 29890 4378
rect 29890 4326 29900 4378
rect 29924 4326 29954 4378
rect 29954 4326 29966 4378
rect 29966 4326 29980 4378
rect 30004 4326 30018 4378
rect 30018 4326 30030 4378
rect 30030 4326 30060 4378
rect 30084 4326 30094 4378
rect 30094 4326 30140 4378
rect 29844 4324 29900 4326
rect 29924 4324 29980 4326
rect 30004 4324 30060 4326
rect 30084 4324 30140 4326
rect 30010 4140 30066 4176
rect 30010 4120 30012 4140
rect 30012 4120 30064 4140
rect 30064 4120 30066 4140
rect 30194 3440 30250 3496
rect 29844 3290 29900 3292
rect 29924 3290 29980 3292
rect 30004 3290 30060 3292
rect 30084 3290 30140 3292
rect 29844 3238 29890 3290
rect 29890 3238 29900 3290
rect 29924 3238 29954 3290
rect 29954 3238 29966 3290
rect 29966 3238 29980 3290
rect 30004 3238 30018 3290
rect 30018 3238 30030 3290
rect 30030 3238 30060 3290
rect 30084 3238 30094 3290
rect 30094 3238 30140 3290
rect 29844 3236 29900 3238
rect 29924 3236 29980 3238
rect 30004 3236 30060 3238
rect 30084 3236 30140 3238
rect 34242 16632 34298 16688
rect 32678 7792 32734 7848
rect 33598 7404 33654 7440
rect 33598 7384 33600 7404
rect 33600 7384 33652 7404
rect 33652 7384 33654 7404
rect 34978 9580 35034 9616
rect 34978 9560 34980 9580
rect 34980 9560 35032 9580
rect 35032 9560 35034 9580
rect 33506 3032 33562 3088
rect 29844 2202 29900 2204
rect 29924 2202 29980 2204
rect 30004 2202 30060 2204
rect 30084 2202 30140 2204
rect 29844 2150 29890 2202
rect 29890 2150 29900 2202
rect 29924 2150 29954 2202
rect 29954 2150 29966 2202
rect 29966 2150 29980 2202
rect 30004 2150 30018 2202
rect 30018 2150 30030 2202
rect 30030 2150 30060 2202
rect 30084 2150 30094 2202
rect 30094 2150 30140 2202
rect 29844 2148 29900 2150
rect 29924 2148 29980 2150
rect 30004 2148 30060 2150
rect 30084 2148 30140 2150
rect 37066 23418 37122 23420
rect 37146 23418 37202 23420
rect 37226 23418 37282 23420
rect 37306 23418 37362 23420
rect 37066 23366 37112 23418
rect 37112 23366 37122 23418
rect 37146 23366 37176 23418
rect 37176 23366 37188 23418
rect 37188 23366 37202 23418
rect 37226 23366 37240 23418
rect 37240 23366 37252 23418
rect 37252 23366 37282 23418
rect 37306 23366 37316 23418
rect 37316 23366 37362 23418
rect 37066 23364 37122 23366
rect 37146 23364 37202 23366
rect 37226 23364 37282 23366
rect 37306 23364 37362 23366
rect 37066 22330 37122 22332
rect 37146 22330 37202 22332
rect 37226 22330 37282 22332
rect 37306 22330 37362 22332
rect 37066 22278 37112 22330
rect 37112 22278 37122 22330
rect 37146 22278 37176 22330
rect 37176 22278 37188 22330
rect 37188 22278 37202 22330
rect 37226 22278 37240 22330
rect 37240 22278 37252 22330
rect 37252 22278 37282 22330
rect 37306 22278 37316 22330
rect 37316 22278 37362 22330
rect 37066 22276 37122 22278
rect 37146 22276 37202 22278
rect 37226 22276 37282 22278
rect 37306 22276 37362 22278
rect 37066 21242 37122 21244
rect 37146 21242 37202 21244
rect 37226 21242 37282 21244
rect 37306 21242 37362 21244
rect 37066 21190 37112 21242
rect 37112 21190 37122 21242
rect 37146 21190 37176 21242
rect 37176 21190 37188 21242
rect 37188 21190 37202 21242
rect 37226 21190 37240 21242
rect 37240 21190 37252 21242
rect 37252 21190 37282 21242
rect 37306 21190 37316 21242
rect 37316 21190 37362 21242
rect 37066 21188 37122 21190
rect 37146 21188 37202 21190
rect 37226 21188 37282 21190
rect 37306 21188 37362 21190
rect 37066 20154 37122 20156
rect 37146 20154 37202 20156
rect 37226 20154 37282 20156
rect 37306 20154 37362 20156
rect 37066 20102 37112 20154
rect 37112 20102 37122 20154
rect 37146 20102 37176 20154
rect 37176 20102 37188 20154
rect 37188 20102 37202 20154
rect 37226 20102 37240 20154
rect 37240 20102 37252 20154
rect 37252 20102 37282 20154
rect 37306 20102 37316 20154
rect 37316 20102 37362 20154
rect 37066 20100 37122 20102
rect 37146 20100 37202 20102
rect 37226 20100 37282 20102
rect 37306 20100 37362 20102
rect 37066 19066 37122 19068
rect 37146 19066 37202 19068
rect 37226 19066 37282 19068
rect 37306 19066 37362 19068
rect 37066 19014 37112 19066
rect 37112 19014 37122 19066
rect 37146 19014 37176 19066
rect 37176 19014 37188 19066
rect 37188 19014 37202 19066
rect 37226 19014 37240 19066
rect 37240 19014 37252 19066
rect 37252 19014 37282 19066
rect 37306 19014 37316 19066
rect 37316 19014 37362 19066
rect 37066 19012 37122 19014
rect 37146 19012 37202 19014
rect 37226 19012 37282 19014
rect 37306 19012 37362 19014
rect 37066 17978 37122 17980
rect 37146 17978 37202 17980
rect 37226 17978 37282 17980
rect 37306 17978 37362 17980
rect 37066 17926 37112 17978
rect 37112 17926 37122 17978
rect 37146 17926 37176 17978
rect 37176 17926 37188 17978
rect 37188 17926 37202 17978
rect 37226 17926 37240 17978
rect 37240 17926 37252 17978
rect 37252 17926 37282 17978
rect 37306 17926 37316 17978
rect 37316 17926 37362 17978
rect 37066 17924 37122 17926
rect 37146 17924 37202 17926
rect 37226 17924 37282 17926
rect 37306 17924 37362 17926
rect 37066 16890 37122 16892
rect 37146 16890 37202 16892
rect 37226 16890 37282 16892
rect 37306 16890 37362 16892
rect 37066 16838 37112 16890
rect 37112 16838 37122 16890
rect 37146 16838 37176 16890
rect 37176 16838 37188 16890
rect 37188 16838 37202 16890
rect 37226 16838 37240 16890
rect 37240 16838 37252 16890
rect 37252 16838 37282 16890
rect 37306 16838 37316 16890
rect 37316 16838 37362 16890
rect 37066 16836 37122 16838
rect 37146 16836 37202 16838
rect 37226 16836 37282 16838
rect 37306 16836 37362 16838
rect 37066 15802 37122 15804
rect 37146 15802 37202 15804
rect 37226 15802 37282 15804
rect 37306 15802 37362 15804
rect 37066 15750 37112 15802
rect 37112 15750 37122 15802
rect 37146 15750 37176 15802
rect 37176 15750 37188 15802
rect 37188 15750 37202 15802
rect 37226 15750 37240 15802
rect 37240 15750 37252 15802
rect 37252 15750 37282 15802
rect 37306 15750 37316 15802
rect 37316 15750 37362 15802
rect 37066 15748 37122 15750
rect 37146 15748 37202 15750
rect 37226 15748 37282 15750
rect 37306 15748 37362 15750
rect 37066 14714 37122 14716
rect 37146 14714 37202 14716
rect 37226 14714 37282 14716
rect 37306 14714 37362 14716
rect 37066 14662 37112 14714
rect 37112 14662 37122 14714
rect 37146 14662 37176 14714
rect 37176 14662 37188 14714
rect 37188 14662 37202 14714
rect 37226 14662 37240 14714
rect 37240 14662 37252 14714
rect 37252 14662 37282 14714
rect 37306 14662 37316 14714
rect 37316 14662 37362 14714
rect 37066 14660 37122 14662
rect 37146 14660 37202 14662
rect 37226 14660 37282 14662
rect 37306 14660 37362 14662
rect 34794 3984 34850 4040
rect 37066 13626 37122 13628
rect 37146 13626 37202 13628
rect 37226 13626 37282 13628
rect 37306 13626 37362 13628
rect 37066 13574 37112 13626
rect 37112 13574 37122 13626
rect 37146 13574 37176 13626
rect 37176 13574 37188 13626
rect 37188 13574 37202 13626
rect 37226 13574 37240 13626
rect 37240 13574 37252 13626
rect 37252 13574 37282 13626
rect 37306 13574 37316 13626
rect 37316 13574 37362 13626
rect 37066 13572 37122 13574
rect 37146 13572 37202 13574
rect 37226 13572 37282 13574
rect 37306 13572 37362 13574
rect 37066 12538 37122 12540
rect 37146 12538 37202 12540
rect 37226 12538 37282 12540
rect 37306 12538 37362 12540
rect 37066 12486 37112 12538
rect 37112 12486 37122 12538
rect 37146 12486 37176 12538
rect 37176 12486 37188 12538
rect 37188 12486 37202 12538
rect 37226 12486 37240 12538
rect 37240 12486 37252 12538
rect 37252 12486 37282 12538
rect 37306 12486 37316 12538
rect 37316 12486 37362 12538
rect 37066 12484 37122 12486
rect 37146 12484 37202 12486
rect 37226 12484 37282 12486
rect 37306 12484 37362 12486
rect 37066 11450 37122 11452
rect 37146 11450 37202 11452
rect 37226 11450 37282 11452
rect 37306 11450 37362 11452
rect 37066 11398 37112 11450
rect 37112 11398 37122 11450
rect 37146 11398 37176 11450
rect 37176 11398 37188 11450
rect 37188 11398 37202 11450
rect 37226 11398 37240 11450
rect 37240 11398 37252 11450
rect 37252 11398 37282 11450
rect 37306 11398 37316 11450
rect 37316 11398 37362 11450
rect 37066 11396 37122 11398
rect 37146 11396 37202 11398
rect 37226 11396 37282 11398
rect 37306 11396 37362 11398
rect 37066 10362 37122 10364
rect 37146 10362 37202 10364
rect 37226 10362 37282 10364
rect 37306 10362 37362 10364
rect 37066 10310 37112 10362
rect 37112 10310 37122 10362
rect 37146 10310 37176 10362
rect 37176 10310 37188 10362
rect 37188 10310 37202 10362
rect 37226 10310 37240 10362
rect 37240 10310 37252 10362
rect 37252 10310 37282 10362
rect 37306 10310 37316 10362
rect 37316 10310 37362 10362
rect 37066 10308 37122 10310
rect 37146 10308 37202 10310
rect 37226 10308 37282 10310
rect 37306 10308 37362 10310
rect 36634 9968 36690 10024
rect 37094 9968 37150 10024
rect 38106 11056 38162 11112
rect 37066 9274 37122 9276
rect 37146 9274 37202 9276
rect 37226 9274 37282 9276
rect 37306 9274 37362 9276
rect 37066 9222 37112 9274
rect 37112 9222 37122 9274
rect 37146 9222 37176 9274
rect 37176 9222 37188 9274
rect 37188 9222 37202 9274
rect 37226 9222 37240 9274
rect 37240 9222 37252 9274
rect 37252 9222 37282 9274
rect 37306 9222 37316 9274
rect 37316 9222 37362 9274
rect 37066 9220 37122 9222
rect 37146 9220 37202 9222
rect 37226 9220 37282 9222
rect 37306 9220 37362 9222
rect 37066 8186 37122 8188
rect 37146 8186 37202 8188
rect 37226 8186 37282 8188
rect 37306 8186 37362 8188
rect 37066 8134 37112 8186
rect 37112 8134 37122 8186
rect 37146 8134 37176 8186
rect 37176 8134 37188 8186
rect 37188 8134 37202 8186
rect 37226 8134 37240 8186
rect 37240 8134 37252 8186
rect 37252 8134 37282 8186
rect 37306 8134 37316 8186
rect 37316 8134 37362 8186
rect 37066 8132 37122 8134
rect 37146 8132 37202 8134
rect 37226 8132 37282 8134
rect 37306 8132 37362 8134
rect 37066 7098 37122 7100
rect 37146 7098 37202 7100
rect 37226 7098 37282 7100
rect 37306 7098 37362 7100
rect 37066 7046 37112 7098
rect 37112 7046 37122 7098
rect 37146 7046 37176 7098
rect 37176 7046 37188 7098
rect 37188 7046 37202 7098
rect 37226 7046 37240 7098
rect 37240 7046 37252 7098
rect 37252 7046 37282 7098
rect 37306 7046 37316 7098
rect 37316 7046 37362 7098
rect 37066 7044 37122 7046
rect 37146 7044 37202 7046
rect 37226 7044 37282 7046
rect 37306 7044 37362 7046
rect 37066 6010 37122 6012
rect 37146 6010 37202 6012
rect 37226 6010 37282 6012
rect 37306 6010 37362 6012
rect 37066 5958 37112 6010
rect 37112 5958 37122 6010
rect 37146 5958 37176 6010
rect 37176 5958 37188 6010
rect 37188 5958 37202 6010
rect 37226 5958 37240 6010
rect 37240 5958 37252 6010
rect 37252 5958 37282 6010
rect 37306 5958 37316 6010
rect 37316 5958 37362 6010
rect 37066 5956 37122 5958
rect 37146 5956 37202 5958
rect 37226 5956 37282 5958
rect 37306 5956 37362 5958
rect 37066 4922 37122 4924
rect 37146 4922 37202 4924
rect 37226 4922 37282 4924
rect 37306 4922 37362 4924
rect 37066 4870 37112 4922
rect 37112 4870 37122 4922
rect 37146 4870 37176 4922
rect 37176 4870 37188 4922
rect 37188 4870 37202 4922
rect 37226 4870 37240 4922
rect 37240 4870 37252 4922
rect 37252 4870 37282 4922
rect 37306 4870 37316 4922
rect 37316 4870 37362 4922
rect 37066 4868 37122 4870
rect 37146 4868 37202 4870
rect 37226 4868 37282 4870
rect 37306 4868 37362 4870
rect 37066 3834 37122 3836
rect 37146 3834 37202 3836
rect 37226 3834 37282 3836
rect 37306 3834 37362 3836
rect 37066 3782 37112 3834
rect 37112 3782 37122 3834
rect 37146 3782 37176 3834
rect 37176 3782 37188 3834
rect 37188 3782 37202 3834
rect 37226 3782 37240 3834
rect 37240 3782 37252 3834
rect 37252 3782 37282 3834
rect 37306 3782 37316 3834
rect 37316 3782 37362 3834
rect 37066 3780 37122 3782
rect 37146 3780 37202 3782
rect 37226 3780 37282 3782
rect 37306 3780 37362 3782
rect 39946 13504 40002 13560
rect 44288 26138 44344 26140
rect 44368 26138 44424 26140
rect 44448 26138 44504 26140
rect 44528 26138 44584 26140
rect 44288 26086 44334 26138
rect 44334 26086 44344 26138
rect 44368 26086 44398 26138
rect 44398 26086 44410 26138
rect 44410 26086 44424 26138
rect 44448 26086 44462 26138
rect 44462 26086 44474 26138
rect 44474 26086 44504 26138
rect 44528 26086 44538 26138
rect 44538 26086 44584 26138
rect 44288 26084 44344 26086
rect 44368 26084 44424 26086
rect 44448 26084 44504 26086
rect 44528 26084 44584 26086
rect 44288 25050 44344 25052
rect 44368 25050 44424 25052
rect 44448 25050 44504 25052
rect 44528 25050 44584 25052
rect 44288 24998 44334 25050
rect 44334 24998 44344 25050
rect 44368 24998 44398 25050
rect 44398 24998 44410 25050
rect 44410 24998 44424 25050
rect 44448 24998 44462 25050
rect 44462 24998 44474 25050
rect 44474 24998 44504 25050
rect 44528 24998 44538 25050
rect 44538 24998 44584 25050
rect 44288 24996 44344 24998
rect 44368 24996 44424 24998
rect 44448 24996 44504 24998
rect 44528 24996 44584 24998
rect 44288 23962 44344 23964
rect 44368 23962 44424 23964
rect 44448 23962 44504 23964
rect 44528 23962 44584 23964
rect 44288 23910 44334 23962
rect 44334 23910 44344 23962
rect 44368 23910 44398 23962
rect 44398 23910 44410 23962
rect 44410 23910 44424 23962
rect 44448 23910 44462 23962
rect 44462 23910 44474 23962
rect 44474 23910 44504 23962
rect 44528 23910 44538 23962
rect 44538 23910 44584 23962
rect 44288 23908 44344 23910
rect 44368 23908 44424 23910
rect 44448 23908 44504 23910
rect 44528 23908 44584 23910
rect 44288 22874 44344 22876
rect 44368 22874 44424 22876
rect 44448 22874 44504 22876
rect 44528 22874 44584 22876
rect 44288 22822 44334 22874
rect 44334 22822 44344 22874
rect 44368 22822 44398 22874
rect 44398 22822 44410 22874
rect 44410 22822 44424 22874
rect 44448 22822 44462 22874
rect 44462 22822 44474 22874
rect 44474 22822 44504 22874
rect 44528 22822 44538 22874
rect 44538 22822 44584 22874
rect 44288 22820 44344 22822
rect 44368 22820 44424 22822
rect 44448 22820 44504 22822
rect 44528 22820 44584 22822
rect 44288 21786 44344 21788
rect 44368 21786 44424 21788
rect 44448 21786 44504 21788
rect 44528 21786 44584 21788
rect 44288 21734 44334 21786
rect 44334 21734 44344 21786
rect 44368 21734 44398 21786
rect 44398 21734 44410 21786
rect 44410 21734 44424 21786
rect 44448 21734 44462 21786
rect 44462 21734 44474 21786
rect 44474 21734 44504 21786
rect 44528 21734 44538 21786
rect 44538 21734 44584 21786
rect 44288 21732 44344 21734
rect 44368 21732 44424 21734
rect 44448 21732 44504 21734
rect 44528 21732 44584 21734
rect 37554 3984 37610 4040
rect 37002 3440 37058 3496
rect 37066 2746 37122 2748
rect 37146 2746 37202 2748
rect 37226 2746 37282 2748
rect 37306 2746 37362 2748
rect 37066 2694 37112 2746
rect 37112 2694 37122 2746
rect 37146 2694 37176 2746
rect 37176 2694 37188 2746
rect 37188 2694 37202 2746
rect 37226 2694 37240 2746
rect 37240 2694 37252 2746
rect 37252 2694 37282 2746
rect 37306 2694 37316 2746
rect 37316 2694 37362 2746
rect 37066 2692 37122 2694
rect 37146 2692 37202 2694
rect 37226 2692 37282 2694
rect 37306 2692 37362 2694
rect 37922 2896 37978 2952
rect 39578 3884 39580 3904
rect 39580 3884 39632 3904
rect 39632 3884 39634 3904
rect 39578 3848 39634 3884
rect 44288 20698 44344 20700
rect 44368 20698 44424 20700
rect 44448 20698 44504 20700
rect 44528 20698 44584 20700
rect 44288 20646 44334 20698
rect 44334 20646 44344 20698
rect 44368 20646 44398 20698
rect 44398 20646 44410 20698
rect 44410 20646 44424 20698
rect 44448 20646 44462 20698
rect 44462 20646 44474 20698
rect 44474 20646 44504 20698
rect 44528 20646 44538 20698
rect 44538 20646 44584 20698
rect 44288 20644 44344 20646
rect 44368 20644 44424 20646
rect 44448 20644 44504 20646
rect 44528 20644 44584 20646
rect 45742 25472 45798 25528
rect 49882 25492 49938 25528
rect 51510 26682 51566 26684
rect 51590 26682 51646 26684
rect 51670 26682 51726 26684
rect 51750 26682 51806 26684
rect 51510 26630 51556 26682
rect 51556 26630 51566 26682
rect 51590 26630 51620 26682
rect 51620 26630 51632 26682
rect 51632 26630 51646 26682
rect 51670 26630 51684 26682
rect 51684 26630 51696 26682
rect 51696 26630 51726 26682
rect 51750 26630 51760 26682
rect 51760 26630 51806 26682
rect 51510 26628 51566 26630
rect 51590 26628 51646 26630
rect 51670 26628 51726 26630
rect 51750 26628 51806 26630
rect 58732 27226 58788 27228
rect 58812 27226 58868 27228
rect 58892 27226 58948 27228
rect 58972 27226 59028 27228
rect 58732 27174 58778 27226
rect 58778 27174 58788 27226
rect 58812 27174 58842 27226
rect 58842 27174 58854 27226
rect 58854 27174 58868 27226
rect 58892 27174 58906 27226
rect 58906 27174 58918 27226
rect 58918 27174 58948 27226
rect 58972 27174 58982 27226
rect 58982 27174 59028 27226
rect 58732 27172 58788 27174
rect 58812 27172 58868 27174
rect 58892 27172 58948 27174
rect 58972 27172 59028 27174
rect 49882 25472 49884 25492
rect 49884 25472 49936 25492
rect 49936 25472 49938 25492
rect 44288 19610 44344 19612
rect 44368 19610 44424 19612
rect 44448 19610 44504 19612
rect 44528 19610 44584 19612
rect 44288 19558 44334 19610
rect 44334 19558 44344 19610
rect 44368 19558 44398 19610
rect 44398 19558 44410 19610
rect 44410 19558 44424 19610
rect 44448 19558 44462 19610
rect 44462 19558 44474 19610
rect 44474 19558 44504 19610
rect 44528 19558 44538 19610
rect 44538 19558 44584 19610
rect 44288 19556 44344 19558
rect 44368 19556 44424 19558
rect 44448 19556 44504 19558
rect 44528 19556 44584 19558
rect 44288 18522 44344 18524
rect 44368 18522 44424 18524
rect 44448 18522 44504 18524
rect 44528 18522 44584 18524
rect 44288 18470 44334 18522
rect 44334 18470 44344 18522
rect 44368 18470 44398 18522
rect 44398 18470 44410 18522
rect 44410 18470 44424 18522
rect 44448 18470 44462 18522
rect 44462 18470 44474 18522
rect 44474 18470 44504 18522
rect 44528 18470 44538 18522
rect 44538 18470 44584 18522
rect 44288 18468 44344 18470
rect 44368 18468 44424 18470
rect 44448 18468 44504 18470
rect 44528 18468 44584 18470
rect 44288 17434 44344 17436
rect 44368 17434 44424 17436
rect 44448 17434 44504 17436
rect 44528 17434 44584 17436
rect 44288 17382 44334 17434
rect 44334 17382 44344 17434
rect 44368 17382 44398 17434
rect 44398 17382 44410 17434
rect 44410 17382 44424 17434
rect 44448 17382 44462 17434
rect 44462 17382 44474 17434
rect 44474 17382 44504 17434
rect 44528 17382 44538 17434
rect 44538 17382 44584 17434
rect 44288 17380 44344 17382
rect 44368 17380 44424 17382
rect 44448 17380 44504 17382
rect 44528 17380 44584 17382
rect 44288 16346 44344 16348
rect 44368 16346 44424 16348
rect 44448 16346 44504 16348
rect 44528 16346 44584 16348
rect 44288 16294 44334 16346
rect 44334 16294 44344 16346
rect 44368 16294 44398 16346
rect 44398 16294 44410 16346
rect 44410 16294 44424 16346
rect 44448 16294 44462 16346
rect 44462 16294 44474 16346
rect 44474 16294 44504 16346
rect 44528 16294 44538 16346
rect 44538 16294 44584 16346
rect 44288 16292 44344 16294
rect 44368 16292 44424 16294
rect 44448 16292 44504 16294
rect 44528 16292 44584 16294
rect 44288 15258 44344 15260
rect 44368 15258 44424 15260
rect 44448 15258 44504 15260
rect 44528 15258 44584 15260
rect 44288 15206 44334 15258
rect 44334 15206 44344 15258
rect 44368 15206 44398 15258
rect 44398 15206 44410 15258
rect 44410 15206 44424 15258
rect 44448 15206 44462 15258
rect 44462 15206 44474 15258
rect 44474 15206 44504 15258
rect 44528 15206 44538 15258
rect 44538 15206 44584 15258
rect 44288 15204 44344 15206
rect 44368 15204 44424 15206
rect 44448 15204 44504 15206
rect 44528 15204 44584 15206
rect 44288 14170 44344 14172
rect 44368 14170 44424 14172
rect 44448 14170 44504 14172
rect 44528 14170 44584 14172
rect 44288 14118 44334 14170
rect 44334 14118 44344 14170
rect 44368 14118 44398 14170
rect 44398 14118 44410 14170
rect 44410 14118 44424 14170
rect 44448 14118 44462 14170
rect 44462 14118 44474 14170
rect 44474 14118 44504 14170
rect 44528 14118 44538 14170
rect 44538 14118 44584 14170
rect 44288 14116 44344 14118
rect 44368 14116 44424 14118
rect 44448 14116 44504 14118
rect 44528 14116 44584 14118
rect 44288 13082 44344 13084
rect 44368 13082 44424 13084
rect 44448 13082 44504 13084
rect 44528 13082 44584 13084
rect 44288 13030 44334 13082
rect 44334 13030 44344 13082
rect 44368 13030 44398 13082
rect 44398 13030 44410 13082
rect 44410 13030 44424 13082
rect 44448 13030 44462 13082
rect 44462 13030 44474 13082
rect 44474 13030 44504 13082
rect 44528 13030 44538 13082
rect 44538 13030 44584 13082
rect 44288 13028 44344 13030
rect 44368 13028 44424 13030
rect 44448 13028 44504 13030
rect 44528 13028 44584 13030
rect 49606 22072 49662 22128
rect 44288 11994 44344 11996
rect 44368 11994 44424 11996
rect 44448 11994 44504 11996
rect 44528 11994 44584 11996
rect 44288 11942 44334 11994
rect 44334 11942 44344 11994
rect 44368 11942 44398 11994
rect 44398 11942 44410 11994
rect 44410 11942 44424 11994
rect 44448 11942 44462 11994
rect 44462 11942 44474 11994
rect 44474 11942 44504 11994
rect 44528 11942 44538 11994
rect 44538 11942 44584 11994
rect 44288 11940 44344 11942
rect 44368 11940 44424 11942
rect 44448 11940 44504 11942
rect 44528 11940 44584 11942
rect 44288 10906 44344 10908
rect 44368 10906 44424 10908
rect 44448 10906 44504 10908
rect 44528 10906 44584 10908
rect 44288 10854 44334 10906
rect 44334 10854 44344 10906
rect 44368 10854 44398 10906
rect 44398 10854 44410 10906
rect 44410 10854 44424 10906
rect 44448 10854 44462 10906
rect 44462 10854 44474 10906
rect 44474 10854 44504 10906
rect 44528 10854 44538 10906
rect 44538 10854 44584 10906
rect 44288 10852 44344 10854
rect 44368 10852 44424 10854
rect 44448 10852 44504 10854
rect 44528 10852 44584 10854
rect 44288 9818 44344 9820
rect 44368 9818 44424 9820
rect 44448 9818 44504 9820
rect 44528 9818 44584 9820
rect 44288 9766 44334 9818
rect 44334 9766 44344 9818
rect 44368 9766 44398 9818
rect 44398 9766 44410 9818
rect 44410 9766 44424 9818
rect 44448 9766 44462 9818
rect 44462 9766 44474 9818
rect 44474 9766 44504 9818
rect 44528 9766 44538 9818
rect 44538 9766 44584 9818
rect 44288 9764 44344 9766
rect 44368 9764 44424 9766
rect 44448 9764 44504 9766
rect 44528 9764 44584 9766
rect 44288 8730 44344 8732
rect 44368 8730 44424 8732
rect 44448 8730 44504 8732
rect 44528 8730 44584 8732
rect 44288 8678 44334 8730
rect 44334 8678 44344 8730
rect 44368 8678 44398 8730
rect 44398 8678 44410 8730
rect 44410 8678 44424 8730
rect 44448 8678 44462 8730
rect 44462 8678 44474 8730
rect 44474 8678 44504 8730
rect 44528 8678 44538 8730
rect 44538 8678 44584 8730
rect 44288 8676 44344 8678
rect 44368 8676 44424 8678
rect 44448 8676 44504 8678
rect 44528 8676 44584 8678
rect 46202 13504 46258 13560
rect 45374 7828 45376 7848
rect 45376 7828 45428 7848
rect 45428 7828 45430 7848
rect 45374 7792 45430 7828
rect 44288 7642 44344 7644
rect 44368 7642 44424 7644
rect 44448 7642 44504 7644
rect 44528 7642 44584 7644
rect 44288 7590 44334 7642
rect 44334 7590 44344 7642
rect 44368 7590 44398 7642
rect 44398 7590 44410 7642
rect 44410 7590 44424 7642
rect 44448 7590 44462 7642
rect 44462 7590 44474 7642
rect 44474 7590 44504 7642
rect 44528 7590 44538 7642
rect 44538 7590 44584 7642
rect 44288 7588 44344 7590
rect 44368 7588 44424 7590
rect 44448 7588 44504 7590
rect 44528 7588 44584 7590
rect 41234 2760 41290 2816
rect 46478 12144 46534 12200
rect 46478 11076 46534 11112
rect 46478 11056 46480 11076
rect 46480 11056 46532 11076
rect 46532 11056 46534 11076
rect 46202 7792 46258 7848
rect 44288 6554 44344 6556
rect 44368 6554 44424 6556
rect 44448 6554 44504 6556
rect 44528 6554 44584 6556
rect 44288 6502 44334 6554
rect 44334 6502 44344 6554
rect 44368 6502 44398 6554
rect 44398 6502 44410 6554
rect 44410 6502 44424 6554
rect 44448 6502 44462 6554
rect 44462 6502 44474 6554
rect 44474 6502 44504 6554
rect 44528 6502 44538 6554
rect 44538 6502 44584 6554
rect 44288 6500 44344 6502
rect 44368 6500 44424 6502
rect 44448 6500 44504 6502
rect 44528 6500 44584 6502
rect 46846 7828 46848 7848
rect 46848 7828 46900 7848
rect 46900 7828 46902 7848
rect 46846 7792 46902 7828
rect 44288 5466 44344 5468
rect 44368 5466 44424 5468
rect 44448 5466 44504 5468
rect 44528 5466 44584 5468
rect 44288 5414 44334 5466
rect 44334 5414 44344 5466
rect 44368 5414 44398 5466
rect 44398 5414 44410 5466
rect 44410 5414 44424 5466
rect 44448 5414 44462 5466
rect 44462 5414 44474 5466
rect 44474 5414 44504 5466
rect 44528 5414 44538 5466
rect 44538 5414 44584 5466
rect 44288 5412 44344 5414
rect 44368 5412 44424 5414
rect 44448 5412 44504 5414
rect 44528 5412 44584 5414
rect 43442 3984 43498 4040
rect 42246 2896 42302 2952
rect 43350 3460 43406 3496
rect 43350 3440 43352 3460
rect 43352 3440 43404 3460
rect 43404 3440 43406 3460
rect 44288 4378 44344 4380
rect 44368 4378 44424 4380
rect 44448 4378 44504 4380
rect 44528 4378 44584 4380
rect 44288 4326 44334 4378
rect 44334 4326 44344 4378
rect 44368 4326 44398 4378
rect 44398 4326 44410 4378
rect 44410 4326 44424 4378
rect 44448 4326 44462 4378
rect 44462 4326 44474 4378
rect 44474 4326 44504 4378
rect 44528 4326 44538 4378
rect 44538 4326 44584 4378
rect 44288 4324 44344 4326
rect 44368 4324 44424 4326
rect 44448 4324 44504 4326
rect 44528 4324 44584 4326
rect 44178 3884 44180 3904
rect 44180 3884 44232 3904
rect 44232 3884 44234 3904
rect 44178 3848 44234 3884
rect 43902 3576 43958 3632
rect 44288 3290 44344 3292
rect 44368 3290 44424 3292
rect 44448 3290 44504 3292
rect 44528 3290 44584 3292
rect 44288 3238 44334 3290
rect 44334 3238 44344 3290
rect 44368 3238 44398 3290
rect 44398 3238 44410 3290
rect 44410 3238 44424 3290
rect 44448 3238 44462 3290
rect 44462 3238 44474 3290
rect 44474 3238 44504 3290
rect 44528 3238 44538 3290
rect 44538 3238 44584 3290
rect 44288 3236 44344 3238
rect 44368 3236 44424 3238
rect 44448 3236 44504 3238
rect 44528 3236 44584 3238
rect 44288 2202 44344 2204
rect 44368 2202 44424 2204
rect 44448 2202 44504 2204
rect 44528 2202 44584 2204
rect 44288 2150 44334 2202
rect 44334 2150 44344 2202
rect 44368 2150 44398 2202
rect 44398 2150 44410 2202
rect 44410 2150 44424 2202
rect 44448 2150 44462 2202
rect 44462 2150 44474 2202
rect 44474 2150 44504 2202
rect 44528 2150 44538 2202
rect 44538 2150 44584 2202
rect 44288 2148 44344 2150
rect 44368 2148 44424 2150
rect 44448 2148 44504 2150
rect 44528 2148 44584 2150
rect 44822 2760 44878 2816
rect 46386 3984 46442 4040
rect 47214 3440 47270 3496
rect 49514 12144 49570 12200
rect 48410 11056 48466 11112
rect 51510 25594 51566 25596
rect 51590 25594 51646 25596
rect 51670 25594 51726 25596
rect 51750 25594 51806 25596
rect 51510 25542 51556 25594
rect 51556 25542 51566 25594
rect 51590 25542 51620 25594
rect 51620 25542 51632 25594
rect 51632 25542 51646 25594
rect 51670 25542 51684 25594
rect 51684 25542 51696 25594
rect 51696 25542 51726 25594
rect 51750 25542 51760 25594
rect 51760 25542 51806 25594
rect 51510 25540 51566 25542
rect 51590 25540 51646 25542
rect 51670 25540 51726 25542
rect 51750 25540 51806 25542
rect 58732 26138 58788 26140
rect 58812 26138 58868 26140
rect 58892 26138 58948 26140
rect 58972 26138 59028 26140
rect 58732 26086 58778 26138
rect 58778 26086 58788 26138
rect 58812 26086 58842 26138
rect 58842 26086 58854 26138
rect 58854 26086 58868 26138
rect 58892 26086 58906 26138
rect 58906 26086 58918 26138
rect 58918 26086 58948 26138
rect 58972 26086 58982 26138
rect 58982 26086 59028 26138
rect 58732 26084 58788 26086
rect 58812 26084 58868 26086
rect 58892 26084 58948 26086
rect 58972 26084 59028 26086
rect 51510 24506 51566 24508
rect 51590 24506 51646 24508
rect 51670 24506 51726 24508
rect 51750 24506 51806 24508
rect 51510 24454 51556 24506
rect 51556 24454 51566 24506
rect 51590 24454 51620 24506
rect 51620 24454 51632 24506
rect 51632 24454 51646 24506
rect 51670 24454 51684 24506
rect 51684 24454 51696 24506
rect 51696 24454 51726 24506
rect 51750 24454 51760 24506
rect 51760 24454 51806 24506
rect 51510 24452 51566 24454
rect 51590 24452 51646 24454
rect 51670 24452 51726 24454
rect 51750 24452 51806 24454
rect 51510 23418 51566 23420
rect 51590 23418 51646 23420
rect 51670 23418 51726 23420
rect 51750 23418 51806 23420
rect 51510 23366 51556 23418
rect 51556 23366 51566 23418
rect 51590 23366 51620 23418
rect 51620 23366 51632 23418
rect 51632 23366 51646 23418
rect 51670 23366 51684 23418
rect 51684 23366 51696 23418
rect 51696 23366 51726 23418
rect 51750 23366 51760 23418
rect 51760 23366 51806 23418
rect 51510 23364 51566 23366
rect 51590 23364 51646 23366
rect 51670 23364 51726 23366
rect 51750 23364 51806 23366
rect 51510 22330 51566 22332
rect 51590 22330 51646 22332
rect 51670 22330 51726 22332
rect 51750 22330 51806 22332
rect 51510 22278 51556 22330
rect 51556 22278 51566 22330
rect 51590 22278 51620 22330
rect 51620 22278 51632 22330
rect 51632 22278 51646 22330
rect 51670 22278 51684 22330
rect 51684 22278 51696 22330
rect 51696 22278 51726 22330
rect 51750 22278 51760 22330
rect 51760 22278 51806 22330
rect 51510 22276 51566 22278
rect 51590 22276 51646 22278
rect 51670 22276 51726 22278
rect 51750 22276 51806 22278
rect 51510 21242 51566 21244
rect 51590 21242 51646 21244
rect 51670 21242 51726 21244
rect 51750 21242 51806 21244
rect 51510 21190 51556 21242
rect 51556 21190 51566 21242
rect 51590 21190 51620 21242
rect 51620 21190 51632 21242
rect 51632 21190 51646 21242
rect 51670 21190 51684 21242
rect 51684 21190 51696 21242
rect 51696 21190 51726 21242
rect 51750 21190 51760 21242
rect 51760 21190 51806 21242
rect 51510 21188 51566 21190
rect 51590 21188 51646 21190
rect 51670 21188 51726 21190
rect 51750 21188 51806 21190
rect 51510 20154 51566 20156
rect 51590 20154 51646 20156
rect 51670 20154 51726 20156
rect 51750 20154 51806 20156
rect 51510 20102 51556 20154
rect 51556 20102 51566 20154
rect 51590 20102 51620 20154
rect 51620 20102 51632 20154
rect 51632 20102 51646 20154
rect 51670 20102 51684 20154
rect 51684 20102 51696 20154
rect 51696 20102 51726 20154
rect 51750 20102 51760 20154
rect 51760 20102 51806 20154
rect 51510 20100 51566 20102
rect 51590 20100 51646 20102
rect 51670 20100 51726 20102
rect 51750 20100 51806 20102
rect 51510 19066 51566 19068
rect 51590 19066 51646 19068
rect 51670 19066 51726 19068
rect 51750 19066 51806 19068
rect 51510 19014 51556 19066
rect 51556 19014 51566 19066
rect 51590 19014 51620 19066
rect 51620 19014 51632 19066
rect 51632 19014 51646 19066
rect 51670 19014 51684 19066
rect 51684 19014 51696 19066
rect 51696 19014 51726 19066
rect 51750 19014 51760 19066
rect 51760 19014 51806 19066
rect 51510 19012 51566 19014
rect 51590 19012 51646 19014
rect 51670 19012 51726 19014
rect 51750 19012 51806 19014
rect 51510 17978 51566 17980
rect 51590 17978 51646 17980
rect 51670 17978 51726 17980
rect 51750 17978 51806 17980
rect 51510 17926 51556 17978
rect 51556 17926 51566 17978
rect 51590 17926 51620 17978
rect 51620 17926 51632 17978
rect 51632 17926 51646 17978
rect 51670 17926 51684 17978
rect 51684 17926 51696 17978
rect 51696 17926 51726 17978
rect 51750 17926 51760 17978
rect 51760 17926 51806 17978
rect 51510 17924 51566 17926
rect 51590 17924 51646 17926
rect 51670 17924 51726 17926
rect 51750 17924 51806 17926
rect 51510 16890 51566 16892
rect 51590 16890 51646 16892
rect 51670 16890 51726 16892
rect 51750 16890 51806 16892
rect 51510 16838 51556 16890
rect 51556 16838 51566 16890
rect 51590 16838 51620 16890
rect 51620 16838 51632 16890
rect 51632 16838 51646 16890
rect 51670 16838 51684 16890
rect 51684 16838 51696 16890
rect 51696 16838 51726 16890
rect 51750 16838 51760 16890
rect 51760 16838 51806 16890
rect 51510 16836 51566 16838
rect 51590 16836 51646 16838
rect 51670 16836 51726 16838
rect 51750 16836 51806 16838
rect 51510 15802 51566 15804
rect 51590 15802 51646 15804
rect 51670 15802 51726 15804
rect 51750 15802 51806 15804
rect 51510 15750 51556 15802
rect 51556 15750 51566 15802
rect 51590 15750 51620 15802
rect 51620 15750 51632 15802
rect 51632 15750 51646 15802
rect 51670 15750 51684 15802
rect 51684 15750 51696 15802
rect 51696 15750 51726 15802
rect 51750 15750 51760 15802
rect 51760 15750 51806 15802
rect 51510 15748 51566 15750
rect 51590 15748 51646 15750
rect 51670 15748 51726 15750
rect 51750 15748 51806 15750
rect 51510 14714 51566 14716
rect 51590 14714 51646 14716
rect 51670 14714 51726 14716
rect 51750 14714 51806 14716
rect 51510 14662 51556 14714
rect 51556 14662 51566 14714
rect 51590 14662 51620 14714
rect 51620 14662 51632 14714
rect 51632 14662 51646 14714
rect 51670 14662 51684 14714
rect 51684 14662 51696 14714
rect 51696 14662 51726 14714
rect 51750 14662 51760 14714
rect 51760 14662 51806 14714
rect 51510 14660 51566 14662
rect 51590 14660 51646 14662
rect 51670 14660 51726 14662
rect 51750 14660 51806 14662
rect 51510 13626 51566 13628
rect 51590 13626 51646 13628
rect 51670 13626 51726 13628
rect 51750 13626 51806 13628
rect 51510 13574 51556 13626
rect 51556 13574 51566 13626
rect 51590 13574 51620 13626
rect 51620 13574 51632 13626
rect 51632 13574 51646 13626
rect 51670 13574 51684 13626
rect 51684 13574 51696 13626
rect 51696 13574 51726 13626
rect 51750 13574 51760 13626
rect 51760 13574 51806 13626
rect 51510 13572 51566 13574
rect 51590 13572 51646 13574
rect 51670 13572 51726 13574
rect 51750 13572 51806 13574
rect 51510 12538 51566 12540
rect 51590 12538 51646 12540
rect 51670 12538 51726 12540
rect 51750 12538 51806 12540
rect 51510 12486 51556 12538
rect 51556 12486 51566 12538
rect 51590 12486 51620 12538
rect 51620 12486 51632 12538
rect 51632 12486 51646 12538
rect 51670 12486 51684 12538
rect 51684 12486 51696 12538
rect 51696 12486 51726 12538
rect 51750 12486 51760 12538
rect 51760 12486 51806 12538
rect 51510 12484 51566 12486
rect 51590 12484 51646 12486
rect 51670 12484 51726 12486
rect 51750 12484 51806 12486
rect 51262 12144 51318 12200
rect 51510 11450 51566 11452
rect 51590 11450 51646 11452
rect 51670 11450 51726 11452
rect 51750 11450 51806 11452
rect 51510 11398 51556 11450
rect 51556 11398 51566 11450
rect 51590 11398 51620 11450
rect 51620 11398 51632 11450
rect 51632 11398 51646 11450
rect 51670 11398 51684 11450
rect 51684 11398 51696 11450
rect 51696 11398 51726 11450
rect 51750 11398 51760 11450
rect 51760 11398 51806 11450
rect 51510 11396 51566 11398
rect 51590 11396 51646 11398
rect 51670 11396 51726 11398
rect 51750 11396 51806 11398
rect 51510 10362 51566 10364
rect 51590 10362 51646 10364
rect 51670 10362 51726 10364
rect 51750 10362 51806 10364
rect 51510 10310 51556 10362
rect 51556 10310 51566 10362
rect 51590 10310 51620 10362
rect 51620 10310 51632 10362
rect 51632 10310 51646 10362
rect 51670 10310 51684 10362
rect 51684 10310 51696 10362
rect 51696 10310 51726 10362
rect 51750 10310 51760 10362
rect 51760 10310 51806 10362
rect 51510 10308 51566 10310
rect 51590 10308 51646 10310
rect 51670 10308 51726 10310
rect 51750 10308 51806 10310
rect 51510 9274 51566 9276
rect 51590 9274 51646 9276
rect 51670 9274 51726 9276
rect 51750 9274 51806 9276
rect 51510 9222 51556 9274
rect 51556 9222 51566 9274
rect 51590 9222 51620 9274
rect 51620 9222 51632 9274
rect 51632 9222 51646 9274
rect 51670 9222 51684 9274
rect 51684 9222 51696 9274
rect 51696 9222 51726 9274
rect 51750 9222 51760 9274
rect 51760 9222 51806 9274
rect 51510 9220 51566 9222
rect 51590 9220 51646 9222
rect 51670 9220 51726 9222
rect 51750 9220 51806 9222
rect 51510 8186 51566 8188
rect 51590 8186 51646 8188
rect 51670 8186 51726 8188
rect 51750 8186 51806 8188
rect 51510 8134 51556 8186
rect 51556 8134 51566 8186
rect 51590 8134 51620 8186
rect 51620 8134 51632 8186
rect 51632 8134 51646 8186
rect 51670 8134 51684 8186
rect 51684 8134 51696 8186
rect 51696 8134 51726 8186
rect 51750 8134 51760 8186
rect 51760 8134 51806 8186
rect 51510 8132 51566 8134
rect 51590 8132 51646 8134
rect 51670 8132 51726 8134
rect 51750 8132 51806 8134
rect 50434 3984 50490 4040
rect 51510 7098 51566 7100
rect 51590 7098 51646 7100
rect 51670 7098 51726 7100
rect 51750 7098 51806 7100
rect 51510 7046 51556 7098
rect 51556 7046 51566 7098
rect 51590 7046 51620 7098
rect 51620 7046 51632 7098
rect 51632 7046 51646 7098
rect 51670 7046 51684 7098
rect 51684 7046 51696 7098
rect 51696 7046 51726 7098
rect 51750 7046 51760 7098
rect 51760 7046 51806 7098
rect 51510 7044 51566 7046
rect 51590 7044 51646 7046
rect 51670 7044 51726 7046
rect 51750 7044 51806 7046
rect 51510 6010 51566 6012
rect 51590 6010 51646 6012
rect 51670 6010 51726 6012
rect 51750 6010 51806 6012
rect 51510 5958 51556 6010
rect 51556 5958 51566 6010
rect 51590 5958 51620 6010
rect 51620 5958 51632 6010
rect 51632 5958 51646 6010
rect 51670 5958 51684 6010
rect 51684 5958 51696 6010
rect 51696 5958 51726 6010
rect 51750 5958 51760 6010
rect 51760 5958 51806 6010
rect 51510 5956 51566 5958
rect 51590 5956 51646 5958
rect 51670 5956 51726 5958
rect 51750 5956 51806 5958
rect 51510 4922 51566 4924
rect 51590 4922 51646 4924
rect 51670 4922 51726 4924
rect 51750 4922 51806 4924
rect 51510 4870 51556 4922
rect 51556 4870 51566 4922
rect 51590 4870 51620 4922
rect 51620 4870 51632 4922
rect 51632 4870 51646 4922
rect 51670 4870 51684 4922
rect 51684 4870 51696 4922
rect 51696 4870 51726 4922
rect 51750 4870 51760 4922
rect 51760 4870 51806 4922
rect 51510 4868 51566 4870
rect 51590 4868 51646 4870
rect 51670 4868 51726 4870
rect 51750 4868 51806 4870
rect 51510 3834 51566 3836
rect 51590 3834 51646 3836
rect 51670 3834 51726 3836
rect 51750 3834 51806 3836
rect 51510 3782 51556 3834
rect 51556 3782 51566 3834
rect 51590 3782 51620 3834
rect 51620 3782 51632 3834
rect 51632 3782 51646 3834
rect 51670 3782 51684 3834
rect 51684 3782 51696 3834
rect 51696 3782 51726 3834
rect 51750 3782 51760 3834
rect 51760 3782 51806 3834
rect 51510 3780 51566 3782
rect 51590 3780 51646 3782
rect 51670 3780 51726 3782
rect 51750 3780 51806 3782
rect 58732 25050 58788 25052
rect 58812 25050 58868 25052
rect 58892 25050 58948 25052
rect 58972 25050 59028 25052
rect 58732 24998 58778 25050
rect 58778 24998 58788 25050
rect 58812 24998 58842 25050
rect 58842 24998 58854 25050
rect 58854 24998 58868 25050
rect 58892 24998 58906 25050
rect 58906 24998 58918 25050
rect 58918 24998 58948 25050
rect 58972 24998 58982 25050
rect 58982 24998 59028 25050
rect 58732 24996 58788 24998
rect 58812 24996 58868 24998
rect 58892 24996 58948 24998
rect 58972 24996 59028 24998
rect 52826 22072 52882 22128
rect 58732 23962 58788 23964
rect 58812 23962 58868 23964
rect 58892 23962 58948 23964
rect 58972 23962 59028 23964
rect 58732 23910 58778 23962
rect 58778 23910 58788 23962
rect 58812 23910 58842 23962
rect 58842 23910 58854 23962
rect 58854 23910 58868 23962
rect 58892 23910 58906 23962
rect 58906 23910 58918 23962
rect 58918 23910 58948 23962
rect 58972 23910 58982 23962
rect 58982 23910 59028 23962
rect 58732 23908 58788 23910
rect 58812 23908 58868 23910
rect 58892 23908 58948 23910
rect 58972 23908 59028 23910
rect 58732 22874 58788 22876
rect 58812 22874 58868 22876
rect 58892 22874 58948 22876
rect 58972 22874 59028 22876
rect 58732 22822 58778 22874
rect 58778 22822 58788 22874
rect 58812 22822 58842 22874
rect 58842 22822 58854 22874
rect 58854 22822 58868 22874
rect 58892 22822 58906 22874
rect 58906 22822 58918 22874
rect 58918 22822 58948 22874
rect 58972 22822 58982 22874
rect 58982 22822 59028 22874
rect 58732 22820 58788 22822
rect 58812 22820 58868 22822
rect 58892 22820 58948 22822
rect 58972 22820 59028 22822
rect 54482 6840 54538 6896
rect 51510 2746 51566 2748
rect 51590 2746 51646 2748
rect 51670 2746 51726 2748
rect 51750 2746 51806 2748
rect 51510 2694 51556 2746
rect 51556 2694 51566 2746
rect 51590 2694 51620 2746
rect 51620 2694 51632 2746
rect 51632 2694 51646 2746
rect 51670 2694 51684 2746
rect 51684 2694 51696 2746
rect 51696 2694 51726 2746
rect 51750 2694 51760 2746
rect 51760 2694 51806 2746
rect 51510 2692 51566 2694
rect 51590 2692 51646 2694
rect 51670 2692 51726 2694
rect 51750 2692 51806 2694
rect 54574 3984 54630 4040
rect 58732 21786 58788 21788
rect 58812 21786 58868 21788
rect 58892 21786 58948 21788
rect 58972 21786 59028 21788
rect 58732 21734 58778 21786
rect 58778 21734 58788 21786
rect 58812 21734 58842 21786
rect 58842 21734 58854 21786
rect 58854 21734 58868 21786
rect 58892 21734 58906 21786
rect 58906 21734 58918 21786
rect 58918 21734 58948 21786
rect 58972 21734 58982 21786
rect 58982 21734 59028 21786
rect 58732 21732 58788 21734
rect 58812 21732 58868 21734
rect 58892 21732 58948 21734
rect 58972 21732 59028 21734
rect 55770 6160 55826 6216
rect 58732 20698 58788 20700
rect 58812 20698 58868 20700
rect 58892 20698 58948 20700
rect 58972 20698 59028 20700
rect 58732 20646 58778 20698
rect 58778 20646 58788 20698
rect 58812 20646 58842 20698
rect 58842 20646 58854 20698
rect 58854 20646 58868 20698
rect 58892 20646 58906 20698
rect 58906 20646 58918 20698
rect 58918 20646 58948 20698
rect 58972 20646 58982 20698
rect 58982 20646 59028 20698
rect 58732 20644 58788 20646
rect 58812 20644 58868 20646
rect 58892 20644 58948 20646
rect 58972 20644 59028 20646
rect 56414 6296 56470 6352
rect 54942 3032 54998 3088
rect 58732 19610 58788 19612
rect 58812 19610 58868 19612
rect 58892 19610 58948 19612
rect 58972 19610 59028 19612
rect 58732 19558 58778 19610
rect 58778 19558 58788 19610
rect 58812 19558 58842 19610
rect 58842 19558 58854 19610
rect 58854 19558 58868 19610
rect 58892 19558 58906 19610
rect 58906 19558 58918 19610
rect 58918 19558 58948 19610
rect 58972 19558 58982 19610
rect 58982 19558 59028 19610
rect 58732 19556 58788 19558
rect 58812 19556 58868 19558
rect 58892 19556 58948 19558
rect 58972 19556 59028 19558
rect 58732 18522 58788 18524
rect 58812 18522 58868 18524
rect 58892 18522 58948 18524
rect 58972 18522 59028 18524
rect 58732 18470 58778 18522
rect 58778 18470 58788 18522
rect 58812 18470 58842 18522
rect 58842 18470 58854 18522
rect 58854 18470 58868 18522
rect 58892 18470 58906 18522
rect 58906 18470 58918 18522
rect 58918 18470 58948 18522
rect 58972 18470 58982 18522
rect 58982 18470 59028 18522
rect 58732 18468 58788 18470
rect 58812 18468 58868 18470
rect 58892 18468 58948 18470
rect 58972 18468 59028 18470
rect 58732 17434 58788 17436
rect 58812 17434 58868 17436
rect 58892 17434 58948 17436
rect 58972 17434 59028 17436
rect 58732 17382 58778 17434
rect 58778 17382 58788 17434
rect 58812 17382 58842 17434
rect 58842 17382 58854 17434
rect 58854 17382 58868 17434
rect 58892 17382 58906 17434
rect 58906 17382 58918 17434
rect 58918 17382 58948 17434
rect 58972 17382 58982 17434
rect 58982 17382 59028 17434
rect 58732 17380 58788 17382
rect 58812 17380 58868 17382
rect 58892 17380 58948 17382
rect 58972 17380 59028 17382
rect 58732 16346 58788 16348
rect 58812 16346 58868 16348
rect 58892 16346 58948 16348
rect 58972 16346 59028 16348
rect 58732 16294 58778 16346
rect 58778 16294 58788 16346
rect 58812 16294 58842 16346
rect 58842 16294 58854 16346
rect 58854 16294 58868 16346
rect 58892 16294 58906 16346
rect 58906 16294 58918 16346
rect 58918 16294 58948 16346
rect 58972 16294 58982 16346
rect 58982 16294 59028 16346
rect 58732 16292 58788 16294
rect 58812 16292 58868 16294
rect 58892 16292 58948 16294
rect 58972 16292 59028 16294
rect 58732 15258 58788 15260
rect 58812 15258 58868 15260
rect 58892 15258 58948 15260
rect 58972 15258 59028 15260
rect 58732 15206 58778 15258
rect 58778 15206 58788 15258
rect 58812 15206 58842 15258
rect 58842 15206 58854 15258
rect 58854 15206 58868 15258
rect 58892 15206 58906 15258
rect 58906 15206 58918 15258
rect 58918 15206 58948 15258
rect 58972 15206 58982 15258
rect 58982 15206 59028 15258
rect 58732 15204 58788 15206
rect 58812 15204 58868 15206
rect 58892 15204 58948 15206
rect 58972 15204 59028 15206
rect 58732 14170 58788 14172
rect 58812 14170 58868 14172
rect 58892 14170 58948 14172
rect 58972 14170 59028 14172
rect 58732 14118 58778 14170
rect 58778 14118 58788 14170
rect 58812 14118 58842 14170
rect 58842 14118 58854 14170
rect 58854 14118 58868 14170
rect 58892 14118 58906 14170
rect 58906 14118 58918 14170
rect 58918 14118 58948 14170
rect 58972 14118 58982 14170
rect 58982 14118 59028 14170
rect 58732 14116 58788 14118
rect 58812 14116 58868 14118
rect 58892 14116 58948 14118
rect 58972 14116 59028 14118
rect 58732 13082 58788 13084
rect 58812 13082 58868 13084
rect 58892 13082 58948 13084
rect 58972 13082 59028 13084
rect 58732 13030 58778 13082
rect 58778 13030 58788 13082
rect 58812 13030 58842 13082
rect 58842 13030 58854 13082
rect 58854 13030 58868 13082
rect 58892 13030 58906 13082
rect 58906 13030 58918 13082
rect 58918 13030 58948 13082
rect 58972 13030 58982 13082
rect 58982 13030 59028 13082
rect 58732 13028 58788 13030
rect 58812 13028 58868 13030
rect 58892 13028 58948 13030
rect 58972 13028 59028 13030
rect 58732 11994 58788 11996
rect 58812 11994 58868 11996
rect 58892 11994 58948 11996
rect 58972 11994 59028 11996
rect 58732 11942 58778 11994
rect 58778 11942 58788 11994
rect 58812 11942 58842 11994
rect 58842 11942 58854 11994
rect 58854 11942 58868 11994
rect 58892 11942 58906 11994
rect 58906 11942 58918 11994
rect 58918 11942 58948 11994
rect 58972 11942 58982 11994
rect 58982 11942 59028 11994
rect 58732 11940 58788 11942
rect 58812 11940 58868 11942
rect 58892 11940 58948 11942
rect 58972 11940 59028 11942
rect 58732 10906 58788 10908
rect 58812 10906 58868 10908
rect 58892 10906 58948 10908
rect 58972 10906 59028 10908
rect 58732 10854 58778 10906
rect 58778 10854 58788 10906
rect 58812 10854 58842 10906
rect 58842 10854 58854 10906
rect 58854 10854 58868 10906
rect 58892 10854 58906 10906
rect 58906 10854 58918 10906
rect 58918 10854 58948 10906
rect 58972 10854 58982 10906
rect 58982 10854 59028 10906
rect 58732 10852 58788 10854
rect 58812 10852 58868 10854
rect 58892 10852 58948 10854
rect 58972 10852 59028 10854
rect 58732 9818 58788 9820
rect 58812 9818 58868 9820
rect 58892 9818 58948 9820
rect 58972 9818 59028 9820
rect 58732 9766 58778 9818
rect 58778 9766 58788 9818
rect 58812 9766 58842 9818
rect 58842 9766 58854 9818
rect 58854 9766 58868 9818
rect 58892 9766 58906 9818
rect 58906 9766 58918 9818
rect 58918 9766 58948 9818
rect 58972 9766 58982 9818
rect 58982 9766 59028 9818
rect 58732 9764 58788 9766
rect 58812 9764 58868 9766
rect 58892 9764 58948 9766
rect 58972 9764 59028 9766
rect 58732 8730 58788 8732
rect 58812 8730 58868 8732
rect 58892 8730 58948 8732
rect 58972 8730 59028 8732
rect 58732 8678 58778 8730
rect 58778 8678 58788 8730
rect 58812 8678 58842 8730
rect 58842 8678 58854 8730
rect 58854 8678 58868 8730
rect 58892 8678 58906 8730
rect 58906 8678 58918 8730
rect 58918 8678 58948 8730
rect 58972 8678 58982 8730
rect 58982 8678 59028 8730
rect 58732 8676 58788 8678
rect 58812 8676 58868 8678
rect 58892 8676 58948 8678
rect 58972 8676 59028 8678
rect 58732 7642 58788 7644
rect 58812 7642 58868 7644
rect 58892 7642 58948 7644
rect 58972 7642 59028 7644
rect 58732 7590 58778 7642
rect 58778 7590 58788 7642
rect 58812 7590 58842 7642
rect 58842 7590 58854 7642
rect 58854 7590 58868 7642
rect 58892 7590 58906 7642
rect 58906 7590 58918 7642
rect 58918 7590 58948 7642
rect 58972 7590 58982 7642
rect 58982 7590 59028 7642
rect 58732 7588 58788 7590
rect 58812 7588 58868 7590
rect 58892 7588 58948 7590
rect 58972 7588 59028 7590
rect 58732 6554 58788 6556
rect 58812 6554 58868 6556
rect 58892 6554 58948 6556
rect 58972 6554 59028 6556
rect 58732 6502 58778 6554
rect 58778 6502 58788 6554
rect 58812 6502 58842 6554
rect 58842 6502 58854 6554
rect 58854 6502 58868 6554
rect 58892 6502 58906 6554
rect 58906 6502 58918 6554
rect 58918 6502 58948 6554
rect 58972 6502 58982 6554
rect 58982 6502 59028 6554
rect 58732 6500 58788 6502
rect 58812 6500 58868 6502
rect 58892 6500 58948 6502
rect 58972 6500 59028 6502
rect 58732 5466 58788 5468
rect 58812 5466 58868 5468
rect 58892 5466 58948 5468
rect 58972 5466 59028 5468
rect 58732 5414 58778 5466
rect 58778 5414 58788 5466
rect 58812 5414 58842 5466
rect 58842 5414 58854 5466
rect 58854 5414 58868 5466
rect 58892 5414 58906 5466
rect 58906 5414 58918 5466
rect 58918 5414 58948 5466
rect 58972 5414 58982 5466
rect 58982 5414 59028 5466
rect 58732 5412 58788 5414
rect 58812 5412 58868 5414
rect 58892 5412 58948 5414
rect 58972 5412 59028 5414
rect 58732 4378 58788 4380
rect 58812 4378 58868 4380
rect 58892 4378 58948 4380
rect 58972 4378 59028 4380
rect 58732 4326 58778 4378
rect 58778 4326 58788 4378
rect 58812 4326 58842 4378
rect 58842 4326 58854 4378
rect 58854 4326 58868 4378
rect 58892 4326 58906 4378
rect 58906 4326 58918 4378
rect 58918 4326 58948 4378
rect 58972 4326 58982 4378
rect 58982 4326 59028 4378
rect 58732 4324 58788 4326
rect 58812 4324 58868 4326
rect 58892 4324 58948 4326
rect 58972 4324 59028 4326
rect 58732 3290 58788 3292
rect 58812 3290 58868 3292
rect 58892 3290 58948 3292
rect 58972 3290 59028 3292
rect 58732 3238 58778 3290
rect 58778 3238 58788 3290
rect 58812 3238 58842 3290
rect 58842 3238 58854 3290
rect 58854 3238 58868 3290
rect 58892 3238 58906 3290
rect 58906 3238 58918 3290
rect 58918 3238 58948 3290
rect 58972 3238 58982 3290
rect 58982 3238 59028 3290
rect 58732 3236 58788 3238
rect 58812 3236 58868 3238
rect 58892 3236 58948 3238
rect 58972 3236 59028 3238
rect 58732 2202 58788 2204
rect 58812 2202 58868 2204
rect 58892 2202 58948 2204
rect 58972 2202 59028 2204
rect 58732 2150 58778 2202
rect 58778 2150 58788 2202
rect 58812 2150 58842 2202
rect 58842 2150 58854 2202
rect 58854 2150 58868 2202
rect 58892 2150 58906 2202
rect 58906 2150 58918 2202
rect 58918 2150 58948 2202
rect 58972 2150 58982 2202
rect 58982 2150 59028 2202
rect 58732 2148 58788 2150
rect 58812 2148 58868 2150
rect 58892 2148 58948 2150
rect 58972 2148 59028 2150
<< metal3 >>
rect 8168 27776 8484 27777
rect 8168 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8484 27776
rect 8168 27711 8484 27712
rect 22612 27776 22928 27777
rect 22612 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22928 27776
rect 22612 27711 22928 27712
rect 37056 27776 37372 27777
rect 37056 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37372 27776
rect 37056 27711 37372 27712
rect 51500 27776 51816 27777
rect 51500 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51816 27776
rect 51500 27711 51816 27712
rect 15390 27232 15706 27233
rect 15390 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15706 27232
rect 15390 27167 15706 27168
rect 29834 27232 30150 27233
rect 29834 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30150 27232
rect 29834 27167 30150 27168
rect 44278 27232 44594 27233
rect 44278 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44594 27232
rect 44278 27167 44594 27168
rect 58722 27232 59038 27233
rect 58722 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59038 27232
rect 58722 27167 59038 27168
rect 8168 26688 8484 26689
rect 8168 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8484 26688
rect 8168 26623 8484 26624
rect 22612 26688 22928 26689
rect 22612 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22928 26688
rect 22612 26623 22928 26624
rect 37056 26688 37372 26689
rect 37056 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37372 26688
rect 37056 26623 37372 26624
rect 51500 26688 51816 26689
rect 51500 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51816 26688
rect 51500 26623 51816 26624
rect 15390 26144 15706 26145
rect 15390 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15706 26144
rect 15390 26079 15706 26080
rect 29834 26144 30150 26145
rect 29834 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30150 26144
rect 29834 26079 30150 26080
rect 44278 26144 44594 26145
rect 44278 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44594 26144
rect 44278 26079 44594 26080
rect 58722 26144 59038 26145
rect 58722 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59038 26144
rect 58722 26079 59038 26080
rect 8168 25600 8484 25601
rect 8168 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8484 25600
rect 8168 25535 8484 25536
rect 22612 25600 22928 25601
rect 22612 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22928 25600
rect 22612 25535 22928 25536
rect 37056 25600 37372 25601
rect 37056 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37372 25600
rect 37056 25535 37372 25536
rect 51500 25600 51816 25601
rect 51500 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51816 25600
rect 51500 25535 51816 25536
rect 45737 25530 45803 25533
rect 49877 25530 49943 25533
rect 45737 25528 49943 25530
rect 45737 25472 45742 25528
rect 45798 25472 49882 25528
rect 49938 25472 49943 25528
rect 45737 25470 49943 25472
rect 45737 25467 45803 25470
rect 49877 25467 49943 25470
rect 15390 25056 15706 25057
rect 15390 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15706 25056
rect 15390 24991 15706 24992
rect 29834 25056 30150 25057
rect 29834 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30150 25056
rect 29834 24991 30150 24992
rect 44278 25056 44594 25057
rect 44278 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44594 25056
rect 44278 24991 44594 24992
rect 58722 25056 59038 25057
rect 58722 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59038 25056
rect 58722 24991 59038 24992
rect 8168 24512 8484 24513
rect 8168 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8484 24512
rect 8168 24447 8484 24448
rect 22612 24512 22928 24513
rect 22612 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22928 24512
rect 22612 24447 22928 24448
rect 37056 24512 37372 24513
rect 37056 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37372 24512
rect 37056 24447 37372 24448
rect 51500 24512 51816 24513
rect 51500 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51816 24512
rect 51500 24447 51816 24448
rect 15390 23968 15706 23969
rect 15390 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15706 23968
rect 15390 23903 15706 23904
rect 29834 23968 30150 23969
rect 29834 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30150 23968
rect 29834 23903 30150 23904
rect 44278 23968 44594 23969
rect 44278 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44594 23968
rect 44278 23903 44594 23904
rect 58722 23968 59038 23969
rect 58722 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59038 23968
rect 58722 23903 59038 23904
rect 8168 23424 8484 23425
rect 8168 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8484 23424
rect 8168 23359 8484 23360
rect 22612 23424 22928 23425
rect 22612 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22928 23424
rect 22612 23359 22928 23360
rect 37056 23424 37372 23425
rect 37056 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37372 23424
rect 37056 23359 37372 23360
rect 51500 23424 51816 23425
rect 51500 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51816 23424
rect 51500 23359 51816 23360
rect 15390 22880 15706 22881
rect 15390 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15706 22880
rect 15390 22815 15706 22816
rect 29834 22880 30150 22881
rect 29834 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30150 22880
rect 29834 22815 30150 22816
rect 44278 22880 44594 22881
rect 44278 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44594 22880
rect 44278 22815 44594 22816
rect 58722 22880 59038 22881
rect 58722 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59038 22880
rect 58722 22815 59038 22816
rect 8168 22336 8484 22337
rect 8168 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8484 22336
rect 8168 22271 8484 22272
rect 22612 22336 22928 22337
rect 22612 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22928 22336
rect 22612 22271 22928 22272
rect 37056 22336 37372 22337
rect 37056 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37372 22336
rect 37056 22271 37372 22272
rect 51500 22336 51816 22337
rect 51500 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51816 22336
rect 51500 22271 51816 22272
rect 49601 22130 49667 22133
rect 52821 22130 52887 22133
rect 49601 22128 52887 22130
rect 49601 22072 49606 22128
rect 49662 22072 52826 22128
rect 52882 22072 52887 22128
rect 49601 22070 52887 22072
rect 49601 22067 49667 22070
rect 52821 22067 52887 22070
rect 15390 21792 15706 21793
rect 15390 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15706 21792
rect 15390 21727 15706 21728
rect 29834 21792 30150 21793
rect 29834 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30150 21792
rect 29834 21727 30150 21728
rect 44278 21792 44594 21793
rect 44278 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44594 21792
rect 44278 21727 44594 21728
rect 58722 21792 59038 21793
rect 58722 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59038 21792
rect 58722 21727 59038 21728
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 22612 21248 22928 21249
rect 22612 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22928 21248
rect 22612 21183 22928 21184
rect 37056 21248 37372 21249
rect 37056 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37372 21248
rect 37056 21183 37372 21184
rect 51500 21248 51816 21249
rect 51500 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51816 21248
rect 51500 21183 51816 21184
rect 15390 20704 15706 20705
rect 15390 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15706 20704
rect 15390 20639 15706 20640
rect 29834 20704 30150 20705
rect 29834 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30150 20704
rect 29834 20639 30150 20640
rect 44278 20704 44594 20705
rect 44278 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44594 20704
rect 44278 20639 44594 20640
rect 58722 20704 59038 20705
rect 58722 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59038 20704
rect 58722 20639 59038 20640
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 22612 20160 22928 20161
rect 22612 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22928 20160
rect 22612 20095 22928 20096
rect 37056 20160 37372 20161
rect 37056 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37372 20160
rect 37056 20095 37372 20096
rect 51500 20160 51816 20161
rect 51500 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51816 20160
rect 51500 20095 51816 20096
rect 15390 19616 15706 19617
rect 15390 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15706 19616
rect 15390 19551 15706 19552
rect 29834 19616 30150 19617
rect 29834 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30150 19616
rect 29834 19551 30150 19552
rect 44278 19616 44594 19617
rect 44278 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44594 19616
rect 44278 19551 44594 19552
rect 58722 19616 59038 19617
rect 58722 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59038 19616
rect 58722 19551 59038 19552
rect 10041 19410 10107 19413
rect 10174 19410 10180 19412
rect 10041 19408 10180 19410
rect 10041 19352 10046 19408
rect 10102 19352 10180 19408
rect 10041 19350 10180 19352
rect 10041 19347 10107 19350
rect 10174 19348 10180 19350
rect 10244 19348 10250 19412
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 22612 19072 22928 19073
rect 22612 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22928 19072
rect 22612 19007 22928 19008
rect 37056 19072 37372 19073
rect 37056 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37372 19072
rect 37056 19007 37372 19008
rect 51500 19072 51816 19073
rect 51500 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51816 19072
rect 51500 19007 51816 19008
rect 15390 18528 15706 18529
rect 15390 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15706 18528
rect 15390 18463 15706 18464
rect 29834 18528 30150 18529
rect 29834 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30150 18528
rect 29834 18463 30150 18464
rect 44278 18528 44594 18529
rect 44278 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44594 18528
rect 44278 18463 44594 18464
rect 58722 18528 59038 18529
rect 58722 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59038 18528
rect 58722 18463 59038 18464
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 22612 17984 22928 17985
rect 22612 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22928 17984
rect 22612 17919 22928 17920
rect 37056 17984 37372 17985
rect 37056 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37372 17984
rect 37056 17919 37372 17920
rect 51500 17984 51816 17985
rect 51500 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51816 17984
rect 51500 17919 51816 17920
rect 15390 17440 15706 17441
rect 15390 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15706 17440
rect 15390 17375 15706 17376
rect 29834 17440 30150 17441
rect 29834 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30150 17440
rect 29834 17375 30150 17376
rect 44278 17440 44594 17441
rect 44278 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44594 17440
rect 44278 17375 44594 17376
rect 58722 17440 59038 17441
rect 58722 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59038 17440
rect 58722 17375 59038 17376
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 22612 16896 22928 16897
rect 22612 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22928 16896
rect 22612 16831 22928 16832
rect 37056 16896 37372 16897
rect 37056 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37372 16896
rect 37056 16831 37372 16832
rect 51500 16896 51816 16897
rect 51500 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51816 16896
rect 51500 16831 51816 16832
rect 9765 16692 9831 16693
rect 34237 16692 34303 16693
rect 9765 16688 9812 16692
rect 9876 16690 9882 16692
rect 9765 16632 9770 16688
rect 9765 16628 9812 16632
rect 9876 16630 9922 16690
rect 34237 16688 34284 16692
rect 34348 16690 34354 16692
rect 34237 16632 34242 16688
rect 9876 16628 9882 16630
rect 34237 16628 34284 16632
rect 34348 16630 34394 16690
rect 34348 16628 34354 16630
rect 9765 16627 9831 16628
rect 34237 16627 34303 16628
rect 15390 16352 15706 16353
rect 15390 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15706 16352
rect 15390 16287 15706 16288
rect 29834 16352 30150 16353
rect 29834 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30150 16352
rect 29834 16287 30150 16288
rect 44278 16352 44594 16353
rect 44278 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44594 16352
rect 44278 16287 44594 16288
rect 58722 16352 59038 16353
rect 58722 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59038 16352
rect 58722 16287 59038 16288
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 22612 15808 22928 15809
rect 22612 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22928 15808
rect 22612 15743 22928 15744
rect 37056 15808 37372 15809
rect 37056 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37372 15808
rect 37056 15743 37372 15744
rect 51500 15808 51816 15809
rect 51500 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51816 15808
rect 51500 15743 51816 15744
rect 15390 15264 15706 15265
rect 15390 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15706 15264
rect 15390 15199 15706 15200
rect 29834 15264 30150 15265
rect 29834 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30150 15264
rect 29834 15199 30150 15200
rect 44278 15264 44594 15265
rect 44278 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44594 15264
rect 44278 15199 44594 15200
rect 58722 15264 59038 15265
rect 58722 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59038 15264
rect 58722 15199 59038 15200
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 22612 14720 22928 14721
rect 22612 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22928 14720
rect 22612 14655 22928 14656
rect 37056 14720 37372 14721
rect 37056 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37372 14720
rect 37056 14655 37372 14656
rect 51500 14720 51816 14721
rect 51500 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51816 14720
rect 51500 14655 51816 14656
rect 15390 14176 15706 14177
rect 15390 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15706 14176
rect 15390 14111 15706 14112
rect 29834 14176 30150 14177
rect 29834 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30150 14176
rect 29834 14111 30150 14112
rect 44278 14176 44594 14177
rect 44278 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44594 14176
rect 44278 14111 44594 14112
rect 58722 14176 59038 14177
rect 58722 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59038 14176
rect 58722 14111 59038 14112
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 22612 13632 22928 13633
rect 22612 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22928 13632
rect 22612 13567 22928 13568
rect 37056 13632 37372 13633
rect 37056 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37372 13632
rect 37056 13567 37372 13568
rect 51500 13632 51816 13633
rect 51500 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51816 13632
rect 51500 13567 51816 13568
rect 39941 13562 40007 13565
rect 46197 13562 46263 13565
rect 39941 13560 46263 13562
rect 39941 13504 39946 13560
rect 40002 13504 46202 13560
rect 46258 13504 46263 13560
rect 39941 13502 46263 13504
rect 39941 13499 40007 13502
rect 46197 13499 46263 13502
rect 15390 13088 15706 13089
rect 15390 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15706 13088
rect 15390 13023 15706 13024
rect 29834 13088 30150 13089
rect 29834 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30150 13088
rect 29834 13023 30150 13024
rect 44278 13088 44594 13089
rect 44278 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44594 13088
rect 44278 13023 44594 13024
rect 58722 13088 59038 13089
rect 58722 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59038 13088
rect 58722 13023 59038 13024
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 22612 12544 22928 12545
rect 22612 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22928 12544
rect 22612 12479 22928 12480
rect 37056 12544 37372 12545
rect 37056 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37372 12544
rect 37056 12479 37372 12480
rect 51500 12544 51816 12545
rect 51500 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51816 12544
rect 51500 12479 51816 12480
rect 23473 12202 23539 12205
rect 27613 12202 27679 12205
rect 23473 12200 27679 12202
rect 23473 12144 23478 12200
rect 23534 12144 27618 12200
rect 27674 12144 27679 12200
rect 23473 12142 27679 12144
rect 23473 12139 23539 12142
rect 27613 12139 27679 12142
rect 46473 12202 46539 12205
rect 49509 12202 49575 12205
rect 51257 12202 51323 12205
rect 46473 12200 51323 12202
rect 46473 12144 46478 12200
rect 46534 12144 49514 12200
rect 49570 12144 51262 12200
rect 51318 12144 51323 12200
rect 46473 12142 51323 12144
rect 46473 12139 46539 12142
rect 49509 12139 49575 12142
rect 51257 12139 51323 12142
rect 15390 12000 15706 12001
rect 15390 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15706 12000
rect 15390 11935 15706 11936
rect 29834 12000 30150 12001
rect 29834 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30150 12000
rect 29834 11935 30150 11936
rect 44278 12000 44594 12001
rect 44278 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44594 12000
rect 44278 11935 44594 11936
rect 58722 12000 59038 12001
rect 58722 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59038 12000
rect 58722 11935 59038 11936
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 22612 11456 22928 11457
rect 22612 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22928 11456
rect 22612 11391 22928 11392
rect 37056 11456 37372 11457
rect 37056 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37372 11456
rect 37056 11391 37372 11392
rect 51500 11456 51816 11457
rect 51500 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51816 11456
rect 51500 11391 51816 11392
rect 2497 11250 2563 11253
rect 4429 11250 4495 11253
rect 2497 11248 4495 11250
rect 2497 11192 2502 11248
rect 2558 11192 4434 11248
rect 4490 11192 4495 11248
rect 2497 11190 4495 11192
rect 2497 11187 2563 11190
rect 4429 11187 4495 11190
rect 2773 11114 2839 11117
rect 4429 11114 4495 11117
rect 2773 11112 4495 11114
rect 2773 11056 2778 11112
rect 2834 11056 4434 11112
rect 4490 11056 4495 11112
rect 2773 11054 4495 11056
rect 2773 11051 2839 11054
rect 4429 11051 4495 11054
rect 10542 11052 10548 11116
rect 10612 11114 10618 11116
rect 11053 11114 11119 11117
rect 10612 11112 11119 11114
rect 10612 11056 11058 11112
rect 11114 11056 11119 11112
rect 10612 11054 11119 11056
rect 10612 11052 10618 11054
rect 11053 11051 11119 11054
rect 37590 11052 37596 11116
rect 37660 11114 37666 11116
rect 38101 11114 38167 11117
rect 37660 11112 38167 11114
rect 37660 11056 38106 11112
rect 38162 11056 38167 11112
rect 37660 11054 38167 11056
rect 37660 11052 37666 11054
rect 38101 11051 38167 11054
rect 46473 11114 46539 11117
rect 48405 11114 48471 11117
rect 46473 11112 48471 11114
rect 46473 11056 46478 11112
rect 46534 11056 48410 11112
rect 48466 11056 48471 11112
rect 46473 11054 48471 11056
rect 46473 11051 46539 11054
rect 48405 11051 48471 11054
rect 15390 10912 15706 10913
rect 15390 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15706 10912
rect 15390 10847 15706 10848
rect 29834 10912 30150 10913
rect 29834 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30150 10912
rect 29834 10847 30150 10848
rect 44278 10912 44594 10913
rect 44278 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44594 10912
rect 44278 10847 44594 10848
rect 58722 10912 59038 10913
rect 58722 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59038 10912
rect 58722 10847 59038 10848
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 22612 10368 22928 10369
rect 22612 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22928 10368
rect 22612 10303 22928 10304
rect 37056 10368 37372 10369
rect 37056 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37372 10368
rect 37056 10303 37372 10304
rect 51500 10368 51816 10369
rect 51500 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51816 10368
rect 51500 10303 51816 10304
rect 22001 10162 22067 10165
rect 22553 10162 22619 10165
rect 22001 10160 22619 10162
rect 22001 10104 22006 10160
rect 22062 10104 22558 10160
rect 22614 10104 22619 10160
rect 22001 10102 22619 10104
rect 22001 10099 22067 10102
rect 22553 10099 22619 10102
rect 36629 10026 36695 10029
rect 37089 10026 37155 10029
rect 36629 10024 37155 10026
rect 36629 9968 36634 10024
rect 36690 9968 37094 10024
rect 37150 9968 37155 10024
rect 36629 9966 37155 9968
rect 36629 9963 36695 9966
rect 37089 9963 37155 9966
rect 15390 9824 15706 9825
rect 15390 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15706 9824
rect 15390 9759 15706 9760
rect 29834 9824 30150 9825
rect 29834 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30150 9824
rect 29834 9759 30150 9760
rect 44278 9824 44594 9825
rect 44278 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44594 9824
rect 44278 9759 44594 9760
rect 58722 9824 59038 9825
rect 58722 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59038 9824
rect 58722 9759 59038 9760
rect 34278 9556 34284 9620
rect 34348 9618 34354 9620
rect 34973 9618 35039 9621
rect 34348 9616 35039 9618
rect 34348 9560 34978 9616
rect 35034 9560 35039 9616
rect 34348 9558 35039 9560
rect 34348 9556 34354 9558
rect 34973 9555 35039 9558
rect 9673 9482 9739 9485
rect 9806 9482 9812 9484
rect 9673 9480 9812 9482
rect 9673 9424 9678 9480
rect 9734 9424 9812 9480
rect 9673 9422 9812 9424
rect 9673 9419 9739 9422
rect 9806 9420 9812 9422
rect 9876 9420 9882 9484
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 22612 9280 22928 9281
rect 22612 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22928 9280
rect 22612 9215 22928 9216
rect 37056 9280 37372 9281
rect 37056 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37372 9280
rect 37056 9215 37372 9216
rect 51500 9280 51816 9281
rect 51500 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51816 9280
rect 51500 9215 51816 9216
rect 15390 8736 15706 8737
rect 15390 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15706 8736
rect 15390 8671 15706 8672
rect 29834 8736 30150 8737
rect 29834 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30150 8736
rect 29834 8671 30150 8672
rect 44278 8736 44594 8737
rect 44278 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44594 8736
rect 44278 8671 44594 8672
rect 58722 8736 59038 8737
rect 58722 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59038 8736
rect 58722 8671 59038 8672
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 22612 8192 22928 8193
rect 22612 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22928 8192
rect 22612 8127 22928 8128
rect 37056 8192 37372 8193
rect 37056 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37372 8192
rect 37056 8127 37372 8128
rect 51500 8192 51816 8193
rect 51500 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51816 8192
rect 51500 8127 51816 8128
rect 16941 7850 17007 7853
rect 32673 7850 32739 7853
rect 16941 7848 32739 7850
rect 16941 7792 16946 7848
rect 17002 7792 32678 7848
rect 32734 7792 32739 7848
rect 16941 7790 32739 7792
rect 16941 7787 17007 7790
rect 32673 7787 32739 7790
rect 45369 7850 45435 7853
rect 46197 7850 46263 7853
rect 46841 7850 46907 7853
rect 45369 7848 46907 7850
rect 45369 7792 45374 7848
rect 45430 7792 46202 7848
rect 46258 7792 46846 7848
rect 46902 7792 46907 7848
rect 45369 7790 46907 7792
rect 45369 7787 45435 7790
rect 46197 7787 46263 7790
rect 46841 7787 46907 7790
rect 22001 7714 22067 7717
rect 26417 7714 26483 7717
rect 22001 7712 26483 7714
rect 22001 7656 22006 7712
rect 22062 7656 26422 7712
rect 26478 7656 26483 7712
rect 22001 7654 26483 7656
rect 22001 7651 22067 7654
rect 26417 7651 26483 7654
rect 15390 7648 15706 7649
rect 15390 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15706 7648
rect 15390 7583 15706 7584
rect 29834 7648 30150 7649
rect 29834 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30150 7648
rect 29834 7583 30150 7584
rect 44278 7648 44594 7649
rect 44278 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44594 7648
rect 44278 7583 44594 7584
rect 58722 7648 59038 7649
rect 58722 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59038 7648
rect 58722 7583 59038 7584
rect 26049 7442 26115 7445
rect 33593 7442 33659 7445
rect 26049 7440 33659 7442
rect 26049 7384 26054 7440
rect 26110 7384 33598 7440
rect 33654 7384 33659 7440
rect 26049 7382 33659 7384
rect 26049 7379 26115 7382
rect 33593 7379 33659 7382
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 22612 7104 22928 7105
rect 22612 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22928 7104
rect 22612 7039 22928 7040
rect 37056 7104 37372 7105
rect 37056 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37372 7104
rect 37056 7039 37372 7040
rect 51500 7104 51816 7105
rect 51500 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51816 7104
rect 51500 7039 51816 7040
rect 11697 6898 11763 6901
rect 54477 6898 54543 6901
rect 11697 6896 54543 6898
rect 11697 6840 11702 6896
rect 11758 6840 54482 6896
rect 54538 6840 54543 6896
rect 11697 6838 54543 6840
rect 11697 6835 11763 6838
rect 54477 6835 54543 6838
rect 10593 6762 10659 6765
rect 11329 6762 11395 6765
rect 10593 6760 11395 6762
rect 10593 6704 10598 6760
rect 10654 6704 11334 6760
rect 11390 6704 11395 6760
rect 10593 6702 11395 6704
rect 10593 6699 10659 6702
rect 11329 6699 11395 6702
rect 15390 6560 15706 6561
rect 15390 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15706 6560
rect 15390 6495 15706 6496
rect 29834 6560 30150 6561
rect 29834 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30150 6560
rect 29834 6495 30150 6496
rect 44278 6560 44594 6561
rect 44278 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44594 6560
rect 44278 6495 44594 6496
rect 58722 6560 59038 6561
rect 58722 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59038 6560
rect 58722 6495 59038 6496
rect 9949 6354 10015 6357
rect 56409 6354 56475 6357
rect 9949 6352 56475 6354
rect 9949 6296 9954 6352
rect 10010 6296 56414 6352
rect 56470 6296 56475 6352
rect 9949 6294 56475 6296
rect 9949 6291 10015 6294
rect 56409 6291 56475 6294
rect 12893 6218 12959 6221
rect 55765 6218 55831 6221
rect 12893 6216 55831 6218
rect 12893 6160 12898 6216
rect 12954 6160 55770 6216
rect 55826 6160 55831 6216
rect 12893 6158 55831 6160
rect 12893 6155 12959 6158
rect 55765 6155 55831 6158
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 22612 6016 22928 6017
rect 22612 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22928 6016
rect 22612 5951 22928 5952
rect 37056 6016 37372 6017
rect 37056 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37372 6016
rect 37056 5951 37372 5952
rect 51500 6016 51816 6017
rect 51500 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51816 6016
rect 51500 5951 51816 5952
rect 15390 5472 15706 5473
rect 15390 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15706 5472
rect 15390 5407 15706 5408
rect 29834 5472 30150 5473
rect 29834 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30150 5472
rect 29834 5407 30150 5408
rect 44278 5472 44594 5473
rect 44278 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44594 5472
rect 44278 5407 44594 5408
rect 58722 5472 59038 5473
rect 58722 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59038 5472
rect 58722 5407 59038 5408
rect 22001 5130 22067 5133
rect 28901 5130 28967 5133
rect 22001 5128 28967 5130
rect 22001 5072 22006 5128
rect 22062 5072 28906 5128
rect 28962 5072 28967 5128
rect 22001 5070 28967 5072
rect 22001 5067 22067 5070
rect 28901 5067 28967 5070
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 22612 4928 22928 4929
rect 22612 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22928 4928
rect 22612 4863 22928 4864
rect 37056 4928 37372 4929
rect 37056 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37372 4928
rect 37056 4863 37372 4864
rect 51500 4928 51816 4929
rect 51500 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51816 4928
rect 51500 4863 51816 4864
rect 15390 4384 15706 4385
rect 15390 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15706 4384
rect 15390 4319 15706 4320
rect 29834 4384 30150 4385
rect 29834 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30150 4384
rect 29834 4319 30150 4320
rect 44278 4384 44594 4385
rect 44278 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44594 4384
rect 44278 4319 44594 4320
rect 58722 4384 59038 4385
rect 58722 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59038 4384
rect 58722 4319 59038 4320
rect 17861 4314 17927 4317
rect 18873 4314 18939 4317
rect 17861 4312 18939 4314
rect 17861 4256 17866 4312
rect 17922 4256 18878 4312
rect 18934 4256 18939 4312
rect 17861 4254 18939 4256
rect 17861 4251 17927 4254
rect 18873 4251 18939 4254
rect 7189 4178 7255 4181
rect 9213 4178 9279 4181
rect 7189 4176 9279 4178
rect 7189 4120 7194 4176
rect 7250 4120 9218 4176
rect 9274 4120 9279 4176
rect 7189 4118 9279 4120
rect 7189 4115 7255 4118
rect 9213 4115 9279 4118
rect 27153 4178 27219 4181
rect 30005 4178 30071 4181
rect 27153 4176 30071 4178
rect 27153 4120 27158 4176
rect 27214 4120 30010 4176
rect 30066 4120 30071 4176
rect 27153 4118 30071 4120
rect 27153 4115 27219 4118
rect 30005 4115 30071 4118
rect 1577 4042 1643 4045
rect 4797 4042 4863 4045
rect 1577 4040 4863 4042
rect 1577 3984 1582 4040
rect 1638 3984 4802 4040
rect 4858 3984 4863 4040
rect 1577 3982 4863 3984
rect 1577 3979 1643 3982
rect 4797 3979 4863 3982
rect 10501 4044 10567 4045
rect 10501 4040 10548 4044
rect 10612 4042 10618 4044
rect 16757 4042 16823 4045
rect 18505 4042 18571 4045
rect 34789 4042 34855 4045
rect 37549 4042 37615 4045
rect 10501 3984 10506 4040
rect 10501 3980 10548 3984
rect 10612 3982 10658 4042
rect 16757 4040 37615 4042
rect 16757 3984 16762 4040
rect 16818 3984 18510 4040
rect 18566 3984 34794 4040
rect 34850 3984 37554 4040
rect 37610 3984 37615 4040
rect 16757 3982 37615 3984
rect 10612 3980 10618 3982
rect 10501 3979 10567 3980
rect 16757 3979 16823 3982
rect 18505 3979 18571 3982
rect 34789 3979 34855 3982
rect 37549 3979 37615 3982
rect 43437 4042 43503 4045
rect 46381 4042 46447 4045
rect 43437 4040 46447 4042
rect 43437 3984 43442 4040
rect 43498 3984 46386 4040
rect 46442 3984 46447 4040
rect 43437 3982 46447 3984
rect 43437 3979 43503 3982
rect 46381 3979 46447 3982
rect 50429 4042 50495 4045
rect 54569 4042 54635 4045
rect 50429 4040 54635 4042
rect 50429 3984 50434 4040
rect 50490 3984 54574 4040
rect 54630 3984 54635 4040
rect 50429 3982 54635 3984
rect 50429 3979 50495 3982
rect 54569 3979 54635 3982
rect 18229 3906 18295 3909
rect 19241 3906 19307 3909
rect 18229 3904 19307 3906
rect 18229 3848 18234 3904
rect 18290 3848 19246 3904
rect 19302 3848 19307 3904
rect 18229 3846 19307 3848
rect 18229 3843 18295 3846
rect 19241 3843 19307 3846
rect 39573 3906 39639 3909
rect 44173 3906 44239 3909
rect 39573 3904 44239 3906
rect 39573 3848 39578 3904
rect 39634 3848 44178 3904
rect 44234 3848 44239 3904
rect 39573 3846 44239 3848
rect 39573 3843 39639 3846
rect 44173 3843 44239 3846
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 22612 3840 22928 3841
rect 22612 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22928 3840
rect 22612 3775 22928 3776
rect 37056 3840 37372 3841
rect 37056 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37372 3840
rect 37056 3775 37372 3776
rect 51500 3840 51816 3841
rect 51500 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51816 3840
rect 51500 3775 51816 3776
rect 26785 3634 26851 3637
rect 43897 3634 43963 3637
rect 26785 3632 43963 3634
rect 26785 3576 26790 3632
rect 26846 3576 43902 3632
rect 43958 3576 43963 3632
rect 26785 3574 43963 3576
rect 26785 3571 26851 3574
rect 43897 3571 43963 3574
rect 933 3498 999 3501
rect 30189 3498 30255 3501
rect 933 3496 30255 3498
rect 933 3440 938 3496
rect 994 3440 30194 3496
rect 30250 3440 30255 3496
rect 933 3438 30255 3440
rect 933 3435 999 3438
rect 30189 3435 30255 3438
rect 36997 3498 37063 3501
rect 37590 3498 37596 3500
rect 36997 3496 37596 3498
rect 36997 3440 37002 3496
rect 37058 3440 37596 3496
rect 36997 3438 37596 3440
rect 36997 3435 37063 3438
rect 37590 3436 37596 3438
rect 37660 3436 37666 3500
rect 43345 3498 43411 3501
rect 47209 3498 47275 3501
rect 43345 3496 47275 3498
rect 43345 3440 43350 3496
rect 43406 3440 47214 3496
rect 47270 3440 47275 3496
rect 43345 3438 47275 3440
rect 43345 3435 43411 3438
rect 47209 3435 47275 3438
rect 21633 3362 21699 3365
rect 22093 3362 22159 3365
rect 21633 3360 22159 3362
rect 21633 3304 21638 3360
rect 21694 3304 22098 3360
rect 22154 3304 22159 3360
rect 21633 3302 22159 3304
rect 21633 3299 21699 3302
rect 22093 3299 22159 3302
rect 15390 3296 15706 3297
rect 15390 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15706 3296
rect 15390 3231 15706 3232
rect 29834 3296 30150 3297
rect 29834 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30150 3296
rect 29834 3231 30150 3232
rect 44278 3296 44594 3297
rect 44278 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44594 3296
rect 44278 3231 44594 3232
rect 58722 3296 59038 3297
rect 58722 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59038 3296
rect 58722 3231 59038 3232
rect 21449 3090 21515 3093
rect 22737 3090 22803 3093
rect 21449 3088 22803 3090
rect 21449 3032 21454 3088
rect 21510 3032 22742 3088
rect 22798 3032 22803 3088
rect 21449 3030 22803 3032
rect 21449 3027 21515 3030
rect 22737 3027 22803 3030
rect 33501 3090 33567 3093
rect 54937 3090 55003 3093
rect 33501 3088 55003 3090
rect 33501 3032 33506 3088
rect 33562 3032 54942 3088
rect 54998 3032 55003 3088
rect 33501 3030 55003 3032
rect 33501 3027 33567 3030
rect 54937 3027 55003 3030
rect 2221 2954 2287 2957
rect 6361 2954 6427 2957
rect 2221 2952 6427 2954
rect 2221 2896 2226 2952
rect 2282 2896 6366 2952
rect 6422 2896 6427 2952
rect 2221 2894 6427 2896
rect 2221 2891 2287 2894
rect 6361 2891 6427 2894
rect 8109 2954 8175 2957
rect 26601 2954 26667 2957
rect 8109 2952 26667 2954
rect 8109 2896 8114 2952
rect 8170 2896 26606 2952
rect 26662 2896 26667 2952
rect 8109 2894 26667 2896
rect 8109 2891 8175 2894
rect 26601 2891 26667 2894
rect 37917 2954 37983 2957
rect 42241 2954 42307 2957
rect 37917 2952 42307 2954
rect 37917 2896 37922 2952
rect 37978 2896 42246 2952
rect 42302 2896 42307 2952
rect 37917 2894 42307 2896
rect 37917 2891 37983 2894
rect 42241 2891 42307 2894
rect 41229 2818 41295 2821
rect 44817 2818 44883 2821
rect 41229 2816 44883 2818
rect 41229 2760 41234 2816
rect 41290 2760 44822 2816
rect 44878 2760 44883 2816
rect 41229 2758 44883 2760
rect 41229 2755 41295 2758
rect 44817 2755 44883 2758
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 22612 2752 22928 2753
rect 22612 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22928 2752
rect 22612 2687 22928 2688
rect 37056 2752 37372 2753
rect 37056 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37372 2752
rect 37056 2687 37372 2688
rect 51500 2752 51816 2753
rect 51500 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51816 2752
rect 51500 2687 51816 2688
rect 15390 2208 15706 2209
rect 15390 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15706 2208
rect 15390 2143 15706 2144
rect 29834 2208 30150 2209
rect 29834 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30150 2208
rect 29834 2143 30150 2144
rect 44278 2208 44594 2209
rect 44278 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44594 2208
rect 44278 2143 44594 2144
rect 58722 2208 59038 2209
rect 58722 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59038 2208
rect 58722 2143 59038 2144
<< via3 >>
rect 8174 27772 8238 27776
rect 8174 27716 8178 27772
rect 8178 27716 8234 27772
rect 8234 27716 8238 27772
rect 8174 27712 8238 27716
rect 8254 27772 8318 27776
rect 8254 27716 8258 27772
rect 8258 27716 8314 27772
rect 8314 27716 8318 27772
rect 8254 27712 8318 27716
rect 8334 27772 8398 27776
rect 8334 27716 8338 27772
rect 8338 27716 8394 27772
rect 8394 27716 8398 27772
rect 8334 27712 8398 27716
rect 8414 27772 8478 27776
rect 8414 27716 8418 27772
rect 8418 27716 8474 27772
rect 8474 27716 8478 27772
rect 8414 27712 8478 27716
rect 22618 27772 22682 27776
rect 22618 27716 22622 27772
rect 22622 27716 22678 27772
rect 22678 27716 22682 27772
rect 22618 27712 22682 27716
rect 22698 27772 22762 27776
rect 22698 27716 22702 27772
rect 22702 27716 22758 27772
rect 22758 27716 22762 27772
rect 22698 27712 22762 27716
rect 22778 27772 22842 27776
rect 22778 27716 22782 27772
rect 22782 27716 22838 27772
rect 22838 27716 22842 27772
rect 22778 27712 22842 27716
rect 22858 27772 22922 27776
rect 22858 27716 22862 27772
rect 22862 27716 22918 27772
rect 22918 27716 22922 27772
rect 22858 27712 22922 27716
rect 37062 27772 37126 27776
rect 37062 27716 37066 27772
rect 37066 27716 37122 27772
rect 37122 27716 37126 27772
rect 37062 27712 37126 27716
rect 37142 27772 37206 27776
rect 37142 27716 37146 27772
rect 37146 27716 37202 27772
rect 37202 27716 37206 27772
rect 37142 27712 37206 27716
rect 37222 27772 37286 27776
rect 37222 27716 37226 27772
rect 37226 27716 37282 27772
rect 37282 27716 37286 27772
rect 37222 27712 37286 27716
rect 37302 27772 37366 27776
rect 37302 27716 37306 27772
rect 37306 27716 37362 27772
rect 37362 27716 37366 27772
rect 37302 27712 37366 27716
rect 51506 27772 51570 27776
rect 51506 27716 51510 27772
rect 51510 27716 51566 27772
rect 51566 27716 51570 27772
rect 51506 27712 51570 27716
rect 51586 27772 51650 27776
rect 51586 27716 51590 27772
rect 51590 27716 51646 27772
rect 51646 27716 51650 27772
rect 51586 27712 51650 27716
rect 51666 27772 51730 27776
rect 51666 27716 51670 27772
rect 51670 27716 51726 27772
rect 51726 27716 51730 27772
rect 51666 27712 51730 27716
rect 51746 27772 51810 27776
rect 51746 27716 51750 27772
rect 51750 27716 51806 27772
rect 51806 27716 51810 27772
rect 51746 27712 51810 27716
rect 15396 27228 15460 27232
rect 15396 27172 15400 27228
rect 15400 27172 15456 27228
rect 15456 27172 15460 27228
rect 15396 27168 15460 27172
rect 15476 27228 15540 27232
rect 15476 27172 15480 27228
rect 15480 27172 15536 27228
rect 15536 27172 15540 27228
rect 15476 27168 15540 27172
rect 15556 27228 15620 27232
rect 15556 27172 15560 27228
rect 15560 27172 15616 27228
rect 15616 27172 15620 27228
rect 15556 27168 15620 27172
rect 15636 27228 15700 27232
rect 15636 27172 15640 27228
rect 15640 27172 15696 27228
rect 15696 27172 15700 27228
rect 15636 27168 15700 27172
rect 29840 27228 29904 27232
rect 29840 27172 29844 27228
rect 29844 27172 29900 27228
rect 29900 27172 29904 27228
rect 29840 27168 29904 27172
rect 29920 27228 29984 27232
rect 29920 27172 29924 27228
rect 29924 27172 29980 27228
rect 29980 27172 29984 27228
rect 29920 27168 29984 27172
rect 30000 27228 30064 27232
rect 30000 27172 30004 27228
rect 30004 27172 30060 27228
rect 30060 27172 30064 27228
rect 30000 27168 30064 27172
rect 30080 27228 30144 27232
rect 30080 27172 30084 27228
rect 30084 27172 30140 27228
rect 30140 27172 30144 27228
rect 30080 27168 30144 27172
rect 44284 27228 44348 27232
rect 44284 27172 44288 27228
rect 44288 27172 44344 27228
rect 44344 27172 44348 27228
rect 44284 27168 44348 27172
rect 44364 27228 44428 27232
rect 44364 27172 44368 27228
rect 44368 27172 44424 27228
rect 44424 27172 44428 27228
rect 44364 27168 44428 27172
rect 44444 27228 44508 27232
rect 44444 27172 44448 27228
rect 44448 27172 44504 27228
rect 44504 27172 44508 27228
rect 44444 27168 44508 27172
rect 44524 27228 44588 27232
rect 44524 27172 44528 27228
rect 44528 27172 44584 27228
rect 44584 27172 44588 27228
rect 44524 27168 44588 27172
rect 58728 27228 58792 27232
rect 58728 27172 58732 27228
rect 58732 27172 58788 27228
rect 58788 27172 58792 27228
rect 58728 27168 58792 27172
rect 58808 27228 58872 27232
rect 58808 27172 58812 27228
rect 58812 27172 58868 27228
rect 58868 27172 58872 27228
rect 58808 27168 58872 27172
rect 58888 27228 58952 27232
rect 58888 27172 58892 27228
rect 58892 27172 58948 27228
rect 58948 27172 58952 27228
rect 58888 27168 58952 27172
rect 58968 27228 59032 27232
rect 58968 27172 58972 27228
rect 58972 27172 59028 27228
rect 59028 27172 59032 27228
rect 58968 27168 59032 27172
rect 8174 26684 8238 26688
rect 8174 26628 8178 26684
rect 8178 26628 8234 26684
rect 8234 26628 8238 26684
rect 8174 26624 8238 26628
rect 8254 26684 8318 26688
rect 8254 26628 8258 26684
rect 8258 26628 8314 26684
rect 8314 26628 8318 26684
rect 8254 26624 8318 26628
rect 8334 26684 8398 26688
rect 8334 26628 8338 26684
rect 8338 26628 8394 26684
rect 8394 26628 8398 26684
rect 8334 26624 8398 26628
rect 8414 26684 8478 26688
rect 8414 26628 8418 26684
rect 8418 26628 8474 26684
rect 8474 26628 8478 26684
rect 8414 26624 8478 26628
rect 22618 26684 22682 26688
rect 22618 26628 22622 26684
rect 22622 26628 22678 26684
rect 22678 26628 22682 26684
rect 22618 26624 22682 26628
rect 22698 26684 22762 26688
rect 22698 26628 22702 26684
rect 22702 26628 22758 26684
rect 22758 26628 22762 26684
rect 22698 26624 22762 26628
rect 22778 26684 22842 26688
rect 22778 26628 22782 26684
rect 22782 26628 22838 26684
rect 22838 26628 22842 26684
rect 22778 26624 22842 26628
rect 22858 26684 22922 26688
rect 22858 26628 22862 26684
rect 22862 26628 22918 26684
rect 22918 26628 22922 26684
rect 22858 26624 22922 26628
rect 37062 26684 37126 26688
rect 37062 26628 37066 26684
rect 37066 26628 37122 26684
rect 37122 26628 37126 26684
rect 37062 26624 37126 26628
rect 37142 26684 37206 26688
rect 37142 26628 37146 26684
rect 37146 26628 37202 26684
rect 37202 26628 37206 26684
rect 37142 26624 37206 26628
rect 37222 26684 37286 26688
rect 37222 26628 37226 26684
rect 37226 26628 37282 26684
rect 37282 26628 37286 26684
rect 37222 26624 37286 26628
rect 37302 26684 37366 26688
rect 37302 26628 37306 26684
rect 37306 26628 37362 26684
rect 37362 26628 37366 26684
rect 37302 26624 37366 26628
rect 51506 26684 51570 26688
rect 51506 26628 51510 26684
rect 51510 26628 51566 26684
rect 51566 26628 51570 26684
rect 51506 26624 51570 26628
rect 51586 26684 51650 26688
rect 51586 26628 51590 26684
rect 51590 26628 51646 26684
rect 51646 26628 51650 26684
rect 51586 26624 51650 26628
rect 51666 26684 51730 26688
rect 51666 26628 51670 26684
rect 51670 26628 51726 26684
rect 51726 26628 51730 26684
rect 51666 26624 51730 26628
rect 51746 26684 51810 26688
rect 51746 26628 51750 26684
rect 51750 26628 51806 26684
rect 51806 26628 51810 26684
rect 51746 26624 51810 26628
rect 15396 26140 15460 26144
rect 15396 26084 15400 26140
rect 15400 26084 15456 26140
rect 15456 26084 15460 26140
rect 15396 26080 15460 26084
rect 15476 26140 15540 26144
rect 15476 26084 15480 26140
rect 15480 26084 15536 26140
rect 15536 26084 15540 26140
rect 15476 26080 15540 26084
rect 15556 26140 15620 26144
rect 15556 26084 15560 26140
rect 15560 26084 15616 26140
rect 15616 26084 15620 26140
rect 15556 26080 15620 26084
rect 15636 26140 15700 26144
rect 15636 26084 15640 26140
rect 15640 26084 15696 26140
rect 15696 26084 15700 26140
rect 15636 26080 15700 26084
rect 29840 26140 29904 26144
rect 29840 26084 29844 26140
rect 29844 26084 29900 26140
rect 29900 26084 29904 26140
rect 29840 26080 29904 26084
rect 29920 26140 29984 26144
rect 29920 26084 29924 26140
rect 29924 26084 29980 26140
rect 29980 26084 29984 26140
rect 29920 26080 29984 26084
rect 30000 26140 30064 26144
rect 30000 26084 30004 26140
rect 30004 26084 30060 26140
rect 30060 26084 30064 26140
rect 30000 26080 30064 26084
rect 30080 26140 30144 26144
rect 30080 26084 30084 26140
rect 30084 26084 30140 26140
rect 30140 26084 30144 26140
rect 30080 26080 30144 26084
rect 44284 26140 44348 26144
rect 44284 26084 44288 26140
rect 44288 26084 44344 26140
rect 44344 26084 44348 26140
rect 44284 26080 44348 26084
rect 44364 26140 44428 26144
rect 44364 26084 44368 26140
rect 44368 26084 44424 26140
rect 44424 26084 44428 26140
rect 44364 26080 44428 26084
rect 44444 26140 44508 26144
rect 44444 26084 44448 26140
rect 44448 26084 44504 26140
rect 44504 26084 44508 26140
rect 44444 26080 44508 26084
rect 44524 26140 44588 26144
rect 44524 26084 44528 26140
rect 44528 26084 44584 26140
rect 44584 26084 44588 26140
rect 44524 26080 44588 26084
rect 58728 26140 58792 26144
rect 58728 26084 58732 26140
rect 58732 26084 58788 26140
rect 58788 26084 58792 26140
rect 58728 26080 58792 26084
rect 58808 26140 58872 26144
rect 58808 26084 58812 26140
rect 58812 26084 58868 26140
rect 58868 26084 58872 26140
rect 58808 26080 58872 26084
rect 58888 26140 58952 26144
rect 58888 26084 58892 26140
rect 58892 26084 58948 26140
rect 58948 26084 58952 26140
rect 58888 26080 58952 26084
rect 58968 26140 59032 26144
rect 58968 26084 58972 26140
rect 58972 26084 59028 26140
rect 59028 26084 59032 26140
rect 58968 26080 59032 26084
rect 8174 25596 8238 25600
rect 8174 25540 8178 25596
rect 8178 25540 8234 25596
rect 8234 25540 8238 25596
rect 8174 25536 8238 25540
rect 8254 25596 8318 25600
rect 8254 25540 8258 25596
rect 8258 25540 8314 25596
rect 8314 25540 8318 25596
rect 8254 25536 8318 25540
rect 8334 25596 8398 25600
rect 8334 25540 8338 25596
rect 8338 25540 8394 25596
rect 8394 25540 8398 25596
rect 8334 25536 8398 25540
rect 8414 25596 8478 25600
rect 8414 25540 8418 25596
rect 8418 25540 8474 25596
rect 8474 25540 8478 25596
rect 8414 25536 8478 25540
rect 22618 25596 22682 25600
rect 22618 25540 22622 25596
rect 22622 25540 22678 25596
rect 22678 25540 22682 25596
rect 22618 25536 22682 25540
rect 22698 25596 22762 25600
rect 22698 25540 22702 25596
rect 22702 25540 22758 25596
rect 22758 25540 22762 25596
rect 22698 25536 22762 25540
rect 22778 25596 22842 25600
rect 22778 25540 22782 25596
rect 22782 25540 22838 25596
rect 22838 25540 22842 25596
rect 22778 25536 22842 25540
rect 22858 25596 22922 25600
rect 22858 25540 22862 25596
rect 22862 25540 22918 25596
rect 22918 25540 22922 25596
rect 22858 25536 22922 25540
rect 37062 25596 37126 25600
rect 37062 25540 37066 25596
rect 37066 25540 37122 25596
rect 37122 25540 37126 25596
rect 37062 25536 37126 25540
rect 37142 25596 37206 25600
rect 37142 25540 37146 25596
rect 37146 25540 37202 25596
rect 37202 25540 37206 25596
rect 37142 25536 37206 25540
rect 37222 25596 37286 25600
rect 37222 25540 37226 25596
rect 37226 25540 37282 25596
rect 37282 25540 37286 25596
rect 37222 25536 37286 25540
rect 37302 25596 37366 25600
rect 37302 25540 37306 25596
rect 37306 25540 37362 25596
rect 37362 25540 37366 25596
rect 37302 25536 37366 25540
rect 51506 25596 51570 25600
rect 51506 25540 51510 25596
rect 51510 25540 51566 25596
rect 51566 25540 51570 25596
rect 51506 25536 51570 25540
rect 51586 25596 51650 25600
rect 51586 25540 51590 25596
rect 51590 25540 51646 25596
rect 51646 25540 51650 25596
rect 51586 25536 51650 25540
rect 51666 25596 51730 25600
rect 51666 25540 51670 25596
rect 51670 25540 51726 25596
rect 51726 25540 51730 25596
rect 51666 25536 51730 25540
rect 51746 25596 51810 25600
rect 51746 25540 51750 25596
rect 51750 25540 51806 25596
rect 51806 25540 51810 25596
rect 51746 25536 51810 25540
rect 15396 25052 15460 25056
rect 15396 24996 15400 25052
rect 15400 24996 15456 25052
rect 15456 24996 15460 25052
rect 15396 24992 15460 24996
rect 15476 25052 15540 25056
rect 15476 24996 15480 25052
rect 15480 24996 15536 25052
rect 15536 24996 15540 25052
rect 15476 24992 15540 24996
rect 15556 25052 15620 25056
rect 15556 24996 15560 25052
rect 15560 24996 15616 25052
rect 15616 24996 15620 25052
rect 15556 24992 15620 24996
rect 15636 25052 15700 25056
rect 15636 24996 15640 25052
rect 15640 24996 15696 25052
rect 15696 24996 15700 25052
rect 15636 24992 15700 24996
rect 29840 25052 29904 25056
rect 29840 24996 29844 25052
rect 29844 24996 29900 25052
rect 29900 24996 29904 25052
rect 29840 24992 29904 24996
rect 29920 25052 29984 25056
rect 29920 24996 29924 25052
rect 29924 24996 29980 25052
rect 29980 24996 29984 25052
rect 29920 24992 29984 24996
rect 30000 25052 30064 25056
rect 30000 24996 30004 25052
rect 30004 24996 30060 25052
rect 30060 24996 30064 25052
rect 30000 24992 30064 24996
rect 30080 25052 30144 25056
rect 30080 24996 30084 25052
rect 30084 24996 30140 25052
rect 30140 24996 30144 25052
rect 30080 24992 30144 24996
rect 44284 25052 44348 25056
rect 44284 24996 44288 25052
rect 44288 24996 44344 25052
rect 44344 24996 44348 25052
rect 44284 24992 44348 24996
rect 44364 25052 44428 25056
rect 44364 24996 44368 25052
rect 44368 24996 44424 25052
rect 44424 24996 44428 25052
rect 44364 24992 44428 24996
rect 44444 25052 44508 25056
rect 44444 24996 44448 25052
rect 44448 24996 44504 25052
rect 44504 24996 44508 25052
rect 44444 24992 44508 24996
rect 44524 25052 44588 25056
rect 44524 24996 44528 25052
rect 44528 24996 44584 25052
rect 44584 24996 44588 25052
rect 44524 24992 44588 24996
rect 58728 25052 58792 25056
rect 58728 24996 58732 25052
rect 58732 24996 58788 25052
rect 58788 24996 58792 25052
rect 58728 24992 58792 24996
rect 58808 25052 58872 25056
rect 58808 24996 58812 25052
rect 58812 24996 58868 25052
rect 58868 24996 58872 25052
rect 58808 24992 58872 24996
rect 58888 25052 58952 25056
rect 58888 24996 58892 25052
rect 58892 24996 58948 25052
rect 58948 24996 58952 25052
rect 58888 24992 58952 24996
rect 58968 25052 59032 25056
rect 58968 24996 58972 25052
rect 58972 24996 59028 25052
rect 59028 24996 59032 25052
rect 58968 24992 59032 24996
rect 8174 24508 8238 24512
rect 8174 24452 8178 24508
rect 8178 24452 8234 24508
rect 8234 24452 8238 24508
rect 8174 24448 8238 24452
rect 8254 24508 8318 24512
rect 8254 24452 8258 24508
rect 8258 24452 8314 24508
rect 8314 24452 8318 24508
rect 8254 24448 8318 24452
rect 8334 24508 8398 24512
rect 8334 24452 8338 24508
rect 8338 24452 8394 24508
rect 8394 24452 8398 24508
rect 8334 24448 8398 24452
rect 8414 24508 8478 24512
rect 8414 24452 8418 24508
rect 8418 24452 8474 24508
rect 8474 24452 8478 24508
rect 8414 24448 8478 24452
rect 22618 24508 22682 24512
rect 22618 24452 22622 24508
rect 22622 24452 22678 24508
rect 22678 24452 22682 24508
rect 22618 24448 22682 24452
rect 22698 24508 22762 24512
rect 22698 24452 22702 24508
rect 22702 24452 22758 24508
rect 22758 24452 22762 24508
rect 22698 24448 22762 24452
rect 22778 24508 22842 24512
rect 22778 24452 22782 24508
rect 22782 24452 22838 24508
rect 22838 24452 22842 24508
rect 22778 24448 22842 24452
rect 22858 24508 22922 24512
rect 22858 24452 22862 24508
rect 22862 24452 22918 24508
rect 22918 24452 22922 24508
rect 22858 24448 22922 24452
rect 37062 24508 37126 24512
rect 37062 24452 37066 24508
rect 37066 24452 37122 24508
rect 37122 24452 37126 24508
rect 37062 24448 37126 24452
rect 37142 24508 37206 24512
rect 37142 24452 37146 24508
rect 37146 24452 37202 24508
rect 37202 24452 37206 24508
rect 37142 24448 37206 24452
rect 37222 24508 37286 24512
rect 37222 24452 37226 24508
rect 37226 24452 37282 24508
rect 37282 24452 37286 24508
rect 37222 24448 37286 24452
rect 37302 24508 37366 24512
rect 37302 24452 37306 24508
rect 37306 24452 37362 24508
rect 37362 24452 37366 24508
rect 37302 24448 37366 24452
rect 51506 24508 51570 24512
rect 51506 24452 51510 24508
rect 51510 24452 51566 24508
rect 51566 24452 51570 24508
rect 51506 24448 51570 24452
rect 51586 24508 51650 24512
rect 51586 24452 51590 24508
rect 51590 24452 51646 24508
rect 51646 24452 51650 24508
rect 51586 24448 51650 24452
rect 51666 24508 51730 24512
rect 51666 24452 51670 24508
rect 51670 24452 51726 24508
rect 51726 24452 51730 24508
rect 51666 24448 51730 24452
rect 51746 24508 51810 24512
rect 51746 24452 51750 24508
rect 51750 24452 51806 24508
rect 51806 24452 51810 24508
rect 51746 24448 51810 24452
rect 15396 23964 15460 23968
rect 15396 23908 15400 23964
rect 15400 23908 15456 23964
rect 15456 23908 15460 23964
rect 15396 23904 15460 23908
rect 15476 23964 15540 23968
rect 15476 23908 15480 23964
rect 15480 23908 15536 23964
rect 15536 23908 15540 23964
rect 15476 23904 15540 23908
rect 15556 23964 15620 23968
rect 15556 23908 15560 23964
rect 15560 23908 15616 23964
rect 15616 23908 15620 23964
rect 15556 23904 15620 23908
rect 15636 23964 15700 23968
rect 15636 23908 15640 23964
rect 15640 23908 15696 23964
rect 15696 23908 15700 23964
rect 15636 23904 15700 23908
rect 29840 23964 29904 23968
rect 29840 23908 29844 23964
rect 29844 23908 29900 23964
rect 29900 23908 29904 23964
rect 29840 23904 29904 23908
rect 29920 23964 29984 23968
rect 29920 23908 29924 23964
rect 29924 23908 29980 23964
rect 29980 23908 29984 23964
rect 29920 23904 29984 23908
rect 30000 23964 30064 23968
rect 30000 23908 30004 23964
rect 30004 23908 30060 23964
rect 30060 23908 30064 23964
rect 30000 23904 30064 23908
rect 30080 23964 30144 23968
rect 30080 23908 30084 23964
rect 30084 23908 30140 23964
rect 30140 23908 30144 23964
rect 30080 23904 30144 23908
rect 44284 23964 44348 23968
rect 44284 23908 44288 23964
rect 44288 23908 44344 23964
rect 44344 23908 44348 23964
rect 44284 23904 44348 23908
rect 44364 23964 44428 23968
rect 44364 23908 44368 23964
rect 44368 23908 44424 23964
rect 44424 23908 44428 23964
rect 44364 23904 44428 23908
rect 44444 23964 44508 23968
rect 44444 23908 44448 23964
rect 44448 23908 44504 23964
rect 44504 23908 44508 23964
rect 44444 23904 44508 23908
rect 44524 23964 44588 23968
rect 44524 23908 44528 23964
rect 44528 23908 44584 23964
rect 44584 23908 44588 23964
rect 44524 23904 44588 23908
rect 58728 23964 58792 23968
rect 58728 23908 58732 23964
rect 58732 23908 58788 23964
rect 58788 23908 58792 23964
rect 58728 23904 58792 23908
rect 58808 23964 58872 23968
rect 58808 23908 58812 23964
rect 58812 23908 58868 23964
rect 58868 23908 58872 23964
rect 58808 23904 58872 23908
rect 58888 23964 58952 23968
rect 58888 23908 58892 23964
rect 58892 23908 58948 23964
rect 58948 23908 58952 23964
rect 58888 23904 58952 23908
rect 58968 23964 59032 23968
rect 58968 23908 58972 23964
rect 58972 23908 59028 23964
rect 59028 23908 59032 23964
rect 58968 23904 59032 23908
rect 8174 23420 8238 23424
rect 8174 23364 8178 23420
rect 8178 23364 8234 23420
rect 8234 23364 8238 23420
rect 8174 23360 8238 23364
rect 8254 23420 8318 23424
rect 8254 23364 8258 23420
rect 8258 23364 8314 23420
rect 8314 23364 8318 23420
rect 8254 23360 8318 23364
rect 8334 23420 8398 23424
rect 8334 23364 8338 23420
rect 8338 23364 8394 23420
rect 8394 23364 8398 23420
rect 8334 23360 8398 23364
rect 8414 23420 8478 23424
rect 8414 23364 8418 23420
rect 8418 23364 8474 23420
rect 8474 23364 8478 23420
rect 8414 23360 8478 23364
rect 22618 23420 22682 23424
rect 22618 23364 22622 23420
rect 22622 23364 22678 23420
rect 22678 23364 22682 23420
rect 22618 23360 22682 23364
rect 22698 23420 22762 23424
rect 22698 23364 22702 23420
rect 22702 23364 22758 23420
rect 22758 23364 22762 23420
rect 22698 23360 22762 23364
rect 22778 23420 22842 23424
rect 22778 23364 22782 23420
rect 22782 23364 22838 23420
rect 22838 23364 22842 23420
rect 22778 23360 22842 23364
rect 22858 23420 22922 23424
rect 22858 23364 22862 23420
rect 22862 23364 22918 23420
rect 22918 23364 22922 23420
rect 22858 23360 22922 23364
rect 37062 23420 37126 23424
rect 37062 23364 37066 23420
rect 37066 23364 37122 23420
rect 37122 23364 37126 23420
rect 37062 23360 37126 23364
rect 37142 23420 37206 23424
rect 37142 23364 37146 23420
rect 37146 23364 37202 23420
rect 37202 23364 37206 23420
rect 37142 23360 37206 23364
rect 37222 23420 37286 23424
rect 37222 23364 37226 23420
rect 37226 23364 37282 23420
rect 37282 23364 37286 23420
rect 37222 23360 37286 23364
rect 37302 23420 37366 23424
rect 37302 23364 37306 23420
rect 37306 23364 37362 23420
rect 37362 23364 37366 23420
rect 37302 23360 37366 23364
rect 51506 23420 51570 23424
rect 51506 23364 51510 23420
rect 51510 23364 51566 23420
rect 51566 23364 51570 23420
rect 51506 23360 51570 23364
rect 51586 23420 51650 23424
rect 51586 23364 51590 23420
rect 51590 23364 51646 23420
rect 51646 23364 51650 23420
rect 51586 23360 51650 23364
rect 51666 23420 51730 23424
rect 51666 23364 51670 23420
rect 51670 23364 51726 23420
rect 51726 23364 51730 23420
rect 51666 23360 51730 23364
rect 51746 23420 51810 23424
rect 51746 23364 51750 23420
rect 51750 23364 51806 23420
rect 51806 23364 51810 23420
rect 51746 23360 51810 23364
rect 15396 22876 15460 22880
rect 15396 22820 15400 22876
rect 15400 22820 15456 22876
rect 15456 22820 15460 22876
rect 15396 22816 15460 22820
rect 15476 22876 15540 22880
rect 15476 22820 15480 22876
rect 15480 22820 15536 22876
rect 15536 22820 15540 22876
rect 15476 22816 15540 22820
rect 15556 22876 15620 22880
rect 15556 22820 15560 22876
rect 15560 22820 15616 22876
rect 15616 22820 15620 22876
rect 15556 22816 15620 22820
rect 15636 22876 15700 22880
rect 15636 22820 15640 22876
rect 15640 22820 15696 22876
rect 15696 22820 15700 22876
rect 15636 22816 15700 22820
rect 29840 22876 29904 22880
rect 29840 22820 29844 22876
rect 29844 22820 29900 22876
rect 29900 22820 29904 22876
rect 29840 22816 29904 22820
rect 29920 22876 29984 22880
rect 29920 22820 29924 22876
rect 29924 22820 29980 22876
rect 29980 22820 29984 22876
rect 29920 22816 29984 22820
rect 30000 22876 30064 22880
rect 30000 22820 30004 22876
rect 30004 22820 30060 22876
rect 30060 22820 30064 22876
rect 30000 22816 30064 22820
rect 30080 22876 30144 22880
rect 30080 22820 30084 22876
rect 30084 22820 30140 22876
rect 30140 22820 30144 22876
rect 30080 22816 30144 22820
rect 44284 22876 44348 22880
rect 44284 22820 44288 22876
rect 44288 22820 44344 22876
rect 44344 22820 44348 22876
rect 44284 22816 44348 22820
rect 44364 22876 44428 22880
rect 44364 22820 44368 22876
rect 44368 22820 44424 22876
rect 44424 22820 44428 22876
rect 44364 22816 44428 22820
rect 44444 22876 44508 22880
rect 44444 22820 44448 22876
rect 44448 22820 44504 22876
rect 44504 22820 44508 22876
rect 44444 22816 44508 22820
rect 44524 22876 44588 22880
rect 44524 22820 44528 22876
rect 44528 22820 44584 22876
rect 44584 22820 44588 22876
rect 44524 22816 44588 22820
rect 58728 22876 58792 22880
rect 58728 22820 58732 22876
rect 58732 22820 58788 22876
rect 58788 22820 58792 22876
rect 58728 22816 58792 22820
rect 58808 22876 58872 22880
rect 58808 22820 58812 22876
rect 58812 22820 58868 22876
rect 58868 22820 58872 22876
rect 58808 22816 58872 22820
rect 58888 22876 58952 22880
rect 58888 22820 58892 22876
rect 58892 22820 58948 22876
rect 58948 22820 58952 22876
rect 58888 22816 58952 22820
rect 58968 22876 59032 22880
rect 58968 22820 58972 22876
rect 58972 22820 59028 22876
rect 59028 22820 59032 22876
rect 58968 22816 59032 22820
rect 8174 22332 8238 22336
rect 8174 22276 8178 22332
rect 8178 22276 8234 22332
rect 8234 22276 8238 22332
rect 8174 22272 8238 22276
rect 8254 22332 8318 22336
rect 8254 22276 8258 22332
rect 8258 22276 8314 22332
rect 8314 22276 8318 22332
rect 8254 22272 8318 22276
rect 8334 22332 8398 22336
rect 8334 22276 8338 22332
rect 8338 22276 8394 22332
rect 8394 22276 8398 22332
rect 8334 22272 8398 22276
rect 8414 22332 8478 22336
rect 8414 22276 8418 22332
rect 8418 22276 8474 22332
rect 8474 22276 8478 22332
rect 8414 22272 8478 22276
rect 22618 22332 22682 22336
rect 22618 22276 22622 22332
rect 22622 22276 22678 22332
rect 22678 22276 22682 22332
rect 22618 22272 22682 22276
rect 22698 22332 22762 22336
rect 22698 22276 22702 22332
rect 22702 22276 22758 22332
rect 22758 22276 22762 22332
rect 22698 22272 22762 22276
rect 22778 22332 22842 22336
rect 22778 22276 22782 22332
rect 22782 22276 22838 22332
rect 22838 22276 22842 22332
rect 22778 22272 22842 22276
rect 22858 22332 22922 22336
rect 22858 22276 22862 22332
rect 22862 22276 22918 22332
rect 22918 22276 22922 22332
rect 22858 22272 22922 22276
rect 37062 22332 37126 22336
rect 37062 22276 37066 22332
rect 37066 22276 37122 22332
rect 37122 22276 37126 22332
rect 37062 22272 37126 22276
rect 37142 22332 37206 22336
rect 37142 22276 37146 22332
rect 37146 22276 37202 22332
rect 37202 22276 37206 22332
rect 37142 22272 37206 22276
rect 37222 22332 37286 22336
rect 37222 22276 37226 22332
rect 37226 22276 37282 22332
rect 37282 22276 37286 22332
rect 37222 22272 37286 22276
rect 37302 22332 37366 22336
rect 37302 22276 37306 22332
rect 37306 22276 37362 22332
rect 37362 22276 37366 22332
rect 37302 22272 37366 22276
rect 51506 22332 51570 22336
rect 51506 22276 51510 22332
rect 51510 22276 51566 22332
rect 51566 22276 51570 22332
rect 51506 22272 51570 22276
rect 51586 22332 51650 22336
rect 51586 22276 51590 22332
rect 51590 22276 51646 22332
rect 51646 22276 51650 22332
rect 51586 22272 51650 22276
rect 51666 22332 51730 22336
rect 51666 22276 51670 22332
rect 51670 22276 51726 22332
rect 51726 22276 51730 22332
rect 51666 22272 51730 22276
rect 51746 22332 51810 22336
rect 51746 22276 51750 22332
rect 51750 22276 51806 22332
rect 51806 22276 51810 22332
rect 51746 22272 51810 22276
rect 15396 21788 15460 21792
rect 15396 21732 15400 21788
rect 15400 21732 15456 21788
rect 15456 21732 15460 21788
rect 15396 21728 15460 21732
rect 15476 21788 15540 21792
rect 15476 21732 15480 21788
rect 15480 21732 15536 21788
rect 15536 21732 15540 21788
rect 15476 21728 15540 21732
rect 15556 21788 15620 21792
rect 15556 21732 15560 21788
rect 15560 21732 15616 21788
rect 15616 21732 15620 21788
rect 15556 21728 15620 21732
rect 15636 21788 15700 21792
rect 15636 21732 15640 21788
rect 15640 21732 15696 21788
rect 15696 21732 15700 21788
rect 15636 21728 15700 21732
rect 29840 21788 29904 21792
rect 29840 21732 29844 21788
rect 29844 21732 29900 21788
rect 29900 21732 29904 21788
rect 29840 21728 29904 21732
rect 29920 21788 29984 21792
rect 29920 21732 29924 21788
rect 29924 21732 29980 21788
rect 29980 21732 29984 21788
rect 29920 21728 29984 21732
rect 30000 21788 30064 21792
rect 30000 21732 30004 21788
rect 30004 21732 30060 21788
rect 30060 21732 30064 21788
rect 30000 21728 30064 21732
rect 30080 21788 30144 21792
rect 30080 21732 30084 21788
rect 30084 21732 30140 21788
rect 30140 21732 30144 21788
rect 30080 21728 30144 21732
rect 44284 21788 44348 21792
rect 44284 21732 44288 21788
rect 44288 21732 44344 21788
rect 44344 21732 44348 21788
rect 44284 21728 44348 21732
rect 44364 21788 44428 21792
rect 44364 21732 44368 21788
rect 44368 21732 44424 21788
rect 44424 21732 44428 21788
rect 44364 21728 44428 21732
rect 44444 21788 44508 21792
rect 44444 21732 44448 21788
rect 44448 21732 44504 21788
rect 44504 21732 44508 21788
rect 44444 21728 44508 21732
rect 44524 21788 44588 21792
rect 44524 21732 44528 21788
rect 44528 21732 44584 21788
rect 44584 21732 44588 21788
rect 44524 21728 44588 21732
rect 58728 21788 58792 21792
rect 58728 21732 58732 21788
rect 58732 21732 58788 21788
rect 58788 21732 58792 21788
rect 58728 21728 58792 21732
rect 58808 21788 58872 21792
rect 58808 21732 58812 21788
rect 58812 21732 58868 21788
rect 58868 21732 58872 21788
rect 58808 21728 58872 21732
rect 58888 21788 58952 21792
rect 58888 21732 58892 21788
rect 58892 21732 58948 21788
rect 58948 21732 58952 21788
rect 58888 21728 58952 21732
rect 58968 21788 59032 21792
rect 58968 21732 58972 21788
rect 58972 21732 59028 21788
rect 59028 21732 59032 21788
rect 58968 21728 59032 21732
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 22618 21244 22682 21248
rect 22618 21188 22622 21244
rect 22622 21188 22678 21244
rect 22678 21188 22682 21244
rect 22618 21184 22682 21188
rect 22698 21244 22762 21248
rect 22698 21188 22702 21244
rect 22702 21188 22758 21244
rect 22758 21188 22762 21244
rect 22698 21184 22762 21188
rect 22778 21244 22842 21248
rect 22778 21188 22782 21244
rect 22782 21188 22838 21244
rect 22838 21188 22842 21244
rect 22778 21184 22842 21188
rect 22858 21244 22922 21248
rect 22858 21188 22862 21244
rect 22862 21188 22918 21244
rect 22918 21188 22922 21244
rect 22858 21184 22922 21188
rect 37062 21244 37126 21248
rect 37062 21188 37066 21244
rect 37066 21188 37122 21244
rect 37122 21188 37126 21244
rect 37062 21184 37126 21188
rect 37142 21244 37206 21248
rect 37142 21188 37146 21244
rect 37146 21188 37202 21244
rect 37202 21188 37206 21244
rect 37142 21184 37206 21188
rect 37222 21244 37286 21248
rect 37222 21188 37226 21244
rect 37226 21188 37282 21244
rect 37282 21188 37286 21244
rect 37222 21184 37286 21188
rect 37302 21244 37366 21248
rect 37302 21188 37306 21244
rect 37306 21188 37362 21244
rect 37362 21188 37366 21244
rect 37302 21184 37366 21188
rect 51506 21244 51570 21248
rect 51506 21188 51510 21244
rect 51510 21188 51566 21244
rect 51566 21188 51570 21244
rect 51506 21184 51570 21188
rect 51586 21244 51650 21248
rect 51586 21188 51590 21244
rect 51590 21188 51646 21244
rect 51646 21188 51650 21244
rect 51586 21184 51650 21188
rect 51666 21244 51730 21248
rect 51666 21188 51670 21244
rect 51670 21188 51726 21244
rect 51726 21188 51730 21244
rect 51666 21184 51730 21188
rect 51746 21244 51810 21248
rect 51746 21188 51750 21244
rect 51750 21188 51806 21244
rect 51806 21188 51810 21244
rect 51746 21184 51810 21188
rect 15396 20700 15460 20704
rect 15396 20644 15400 20700
rect 15400 20644 15456 20700
rect 15456 20644 15460 20700
rect 15396 20640 15460 20644
rect 15476 20700 15540 20704
rect 15476 20644 15480 20700
rect 15480 20644 15536 20700
rect 15536 20644 15540 20700
rect 15476 20640 15540 20644
rect 15556 20700 15620 20704
rect 15556 20644 15560 20700
rect 15560 20644 15616 20700
rect 15616 20644 15620 20700
rect 15556 20640 15620 20644
rect 15636 20700 15700 20704
rect 15636 20644 15640 20700
rect 15640 20644 15696 20700
rect 15696 20644 15700 20700
rect 15636 20640 15700 20644
rect 29840 20700 29904 20704
rect 29840 20644 29844 20700
rect 29844 20644 29900 20700
rect 29900 20644 29904 20700
rect 29840 20640 29904 20644
rect 29920 20700 29984 20704
rect 29920 20644 29924 20700
rect 29924 20644 29980 20700
rect 29980 20644 29984 20700
rect 29920 20640 29984 20644
rect 30000 20700 30064 20704
rect 30000 20644 30004 20700
rect 30004 20644 30060 20700
rect 30060 20644 30064 20700
rect 30000 20640 30064 20644
rect 30080 20700 30144 20704
rect 30080 20644 30084 20700
rect 30084 20644 30140 20700
rect 30140 20644 30144 20700
rect 30080 20640 30144 20644
rect 44284 20700 44348 20704
rect 44284 20644 44288 20700
rect 44288 20644 44344 20700
rect 44344 20644 44348 20700
rect 44284 20640 44348 20644
rect 44364 20700 44428 20704
rect 44364 20644 44368 20700
rect 44368 20644 44424 20700
rect 44424 20644 44428 20700
rect 44364 20640 44428 20644
rect 44444 20700 44508 20704
rect 44444 20644 44448 20700
rect 44448 20644 44504 20700
rect 44504 20644 44508 20700
rect 44444 20640 44508 20644
rect 44524 20700 44588 20704
rect 44524 20644 44528 20700
rect 44528 20644 44584 20700
rect 44584 20644 44588 20700
rect 44524 20640 44588 20644
rect 58728 20700 58792 20704
rect 58728 20644 58732 20700
rect 58732 20644 58788 20700
rect 58788 20644 58792 20700
rect 58728 20640 58792 20644
rect 58808 20700 58872 20704
rect 58808 20644 58812 20700
rect 58812 20644 58868 20700
rect 58868 20644 58872 20700
rect 58808 20640 58872 20644
rect 58888 20700 58952 20704
rect 58888 20644 58892 20700
rect 58892 20644 58948 20700
rect 58948 20644 58952 20700
rect 58888 20640 58952 20644
rect 58968 20700 59032 20704
rect 58968 20644 58972 20700
rect 58972 20644 59028 20700
rect 59028 20644 59032 20700
rect 58968 20640 59032 20644
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 22618 20156 22682 20160
rect 22618 20100 22622 20156
rect 22622 20100 22678 20156
rect 22678 20100 22682 20156
rect 22618 20096 22682 20100
rect 22698 20156 22762 20160
rect 22698 20100 22702 20156
rect 22702 20100 22758 20156
rect 22758 20100 22762 20156
rect 22698 20096 22762 20100
rect 22778 20156 22842 20160
rect 22778 20100 22782 20156
rect 22782 20100 22838 20156
rect 22838 20100 22842 20156
rect 22778 20096 22842 20100
rect 22858 20156 22922 20160
rect 22858 20100 22862 20156
rect 22862 20100 22918 20156
rect 22918 20100 22922 20156
rect 22858 20096 22922 20100
rect 37062 20156 37126 20160
rect 37062 20100 37066 20156
rect 37066 20100 37122 20156
rect 37122 20100 37126 20156
rect 37062 20096 37126 20100
rect 37142 20156 37206 20160
rect 37142 20100 37146 20156
rect 37146 20100 37202 20156
rect 37202 20100 37206 20156
rect 37142 20096 37206 20100
rect 37222 20156 37286 20160
rect 37222 20100 37226 20156
rect 37226 20100 37282 20156
rect 37282 20100 37286 20156
rect 37222 20096 37286 20100
rect 37302 20156 37366 20160
rect 37302 20100 37306 20156
rect 37306 20100 37362 20156
rect 37362 20100 37366 20156
rect 37302 20096 37366 20100
rect 51506 20156 51570 20160
rect 51506 20100 51510 20156
rect 51510 20100 51566 20156
rect 51566 20100 51570 20156
rect 51506 20096 51570 20100
rect 51586 20156 51650 20160
rect 51586 20100 51590 20156
rect 51590 20100 51646 20156
rect 51646 20100 51650 20156
rect 51586 20096 51650 20100
rect 51666 20156 51730 20160
rect 51666 20100 51670 20156
rect 51670 20100 51726 20156
rect 51726 20100 51730 20156
rect 51666 20096 51730 20100
rect 51746 20156 51810 20160
rect 51746 20100 51750 20156
rect 51750 20100 51806 20156
rect 51806 20100 51810 20156
rect 51746 20096 51810 20100
rect 15396 19612 15460 19616
rect 15396 19556 15400 19612
rect 15400 19556 15456 19612
rect 15456 19556 15460 19612
rect 15396 19552 15460 19556
rect 15476 19612 15540 19616
rect 15476 19556 15480 19612
rect 15480 19556 15536 19612
rect 15536 19556 15540 19612
rect 15476 19552 15540 19556
rect 15556 19612 15620 19616
rect 15556 19556 15560 19612
rect 15560 19556 15616 19612
rect 15616 19556 15620 19612
rect 15556 19552 15620 19556
rect 15636 19612 15700 19616
rect 15636 19556 15640 19612
rect 15640 19556 15696 19612
rect 15696 19556 15700 19612
rect 15636 19552 15700 19556
rect 29840 19612 29904 19616
rect 29840 19556 29844 19612
rect 29844 19556 29900 19612
rect 29900 19556 29904 19612
rect 29840 19552 29904 19556
rect 29920 19612 29984 19616
rect 29920 19556 29924 19612
rect 29924 19556 29980 19612
rect 29980 19556 29984 19612
rect 29920 19552 29984 19556
rect 30000 19612 30064 19616
rect 30000 19556 30004 19612
rect 30004 19556 30060 19612
rect 30060 19556 30064 19612
rect 30000 19552 30064 19556
rect 30080 19612 30144 19616
rect 30080 19556 30084 19612
rect 30084 19556 30140 19612
rect 30140 19556 30144 19612
rect 30080 19552 30144 19556
rect 44284 19612 44348 19616
rect 44284 19556 44288 19612
rect 44288 19556 44344 19612
rect 44344 19556 44348 19612
rect 44284 19552 44348 19556
rect 44364 19612 44428 19616
rect 44364 19556 44368 19612
rect 44368 19556 44424 19612
rect 44424 19556 44428 19612
rect 44364 19552 44428 19556
rect 44444 19612 44508 19616
rect 44444 19556 44448 19612
rect 44448 19556 44504 19612
rect 44504 19556 44508 19612
rect 44444 19552 44508 19556
rect 44524 19612 44588 19616
rect 44524 19556 44528 19612
rect 44528 19556 44584 19612
rect 44584 19556 44588 19612
rect 44524 19552 44588 19556
rect 58728 19612 58792 19616
rect 58728 19556 58732 19612
rect 58732 19556 58788 19612
rect 58788 19556 58792 19612
rect 58728 19552 58792 19556
rect 58808 19612 58872 19616
rect 58808 19556 58812 19612
rect 58812 19556 58868 19612
rect 58868 19556 58872 19612
rect 58808 19552 58872 19556
rect 58888 19612 58952 19616
rect 58888 19556 58892 19612
rect 58892 19556 58948 19612
rect 58948 19556 58952 19612
rect 58888 19552 58952 19556
rect 58968 19612 59032 19616
rect 58968 19556 58972 19612
rect 58972 19556 59028 19612
rect 59028 19556 59032 19612
rect 58968 19552 59032 19556
rect 10180 19348 10244 19412
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 22618 19068 22682 19072
rect 22618 19012 22622 19068
rect 22622 19012 22678 19068
rect 22678 19012 22682 19068
rect 22618 19008 22682 19012
rect 22698 19068 22762 19072
rect 22698 19012 22702 19068
rect 22702 19012 22758 19068
rect 22758 19012 22762 19068
rect 22698 19008 22762 19012
rect 22778 19068 22842 19072
rect 22778 19012 22782 19068
rect 22782 19012 22838 19068
rect 22838 19012 22842 19068
rect 22778 19008 22842 19012
rect 22858 19068 22922 19072
rect 22858 19012 22862 19068
rect 22862 19012 22918 19068
rect 22918 19012 22922 19068
rect 22858 19008 22922 19012
rect 37062 19068 37126 19072
rect 37062 19012 37066 19068
rect 37066 19012 37122 19068
rect 37122 19012 37126 19068
rect 37062 19008 37126 19012
rect 37142 19068 37206 19072
rect 37142 19012 37146 19068
rect 37146 19012 37202 19068
rect 37202 19012 37206 19068
rect 37142 19008 37206 19012
rect 37222 19068 37286 19072
rect 37222 19012 37226 19068
rect 37226 19012 37282 19068
rect 37282 19012 37286 19068
rect 37222 19008 37286 19012
rect 37302 19068 37366 19072
rect 37302 19012 37306 19068
rect 37306 19012 37362 19068
rect 37362 19012 37366 19068
rect 37302 19008 37366 19012
rect 51506 19068 51570 19072
rect 51506 19012 51510 19068
rect 51510 19012 51566 19068
rect 51566 19012 51570 19068
rect 51506 19008 51570 19012
rect 51586 19068 51650 19072
rect 51586 19012 51590 19068
rect 51590 19012 51646 19068
rect 51646 19012 51650 19068
rect 51586 19008 51650 19012
rect 51666 19068 51730 19072
rect 51666 19012 51670 19068
rect 51670 19012 51726 19068
rect 51726 19012 51730 19068
rect 51666 19008 51730 19012
rect 51746 19068 51810 19072
rect 51746 19012 51750 19068
rect 51750 19012 51806 19068
rect 51806 19012 51810 19068
rect 51746 19008 51810 19012
rect 15396 18524 15460 18528
rect 15396 18468 15400 18524
rect 15400 18468 15456 18524
rect 15456 18468 15460 18524
rect 15396 18464 15460 18468
rect 15476 18524 15540 18528
rect 15476 18468 15480 18524
rect 15480 18468 15536 18524
rect 15536 18468 15540 18524
rect 15476 18464 15540 18468
rect 15556 18524 15620 18528
rect 15556 18468 15560 18524
rect 15560 18468 15616 18524
rect 15616 18468 15620 18524
rect 15556 18464 15620 18468
rect 15636 18524 15700 18528
rect 15636 18468 15640 18524
rect 15640 18468 15696 18524
rect 15696 18468 15700 18524
rect 15636 18464 15700 18468
rect 29840 18524 29904 18528
rect 29840 18468 29844 18524
rect 29844 18468 29900 18524
rect 29900 18468 29904 18524
rect 29840 18464 29904 18468
rect 29920 18524 29984 18528
rect 29920 18468 29924 18524
rect 29924 18468 29980 18524
rect 29980 18468 29984 18524
rect 29920 18464 29984 18468
rect 30000 18524 30064 18528
rect 30000 18468 30004 18524
rect 30004 18468 30060 18524
rect 30060 18468 30064 18524
rect 30000 18464 30064 18468
rect 30080 18524 30144 18528
rect 30080 18468 30084 18524
rect 30084 18468 30140 18524
rect 30140 18468 30144 18524
rect 30080 18464 30144 18468
rect 44284 18524 44348 18528
rect 44284 18468 44288 18524
rect 44288 18468 44344 18524
rect 44344 18468 44348 18524
rect 44284 18464 44348 18468
rect 44364 18524 44428 18528
rect 44364 18468 44368 18524
rect 44368 18468 44424 18524
rect 44424 18468 44428 18524
rect 44364 18464 44428 18468
rect 44444 18524 44508 18528
rect 44444 18468 44448 18524
rect 44448 18468 44504 18524
rect 44504 18468 44508 18524
rect 44444 18464 44508 18468
rect 44524 18524 44588 18528
rect 44524 18468 44528 18524
rect 44528 18468 44584 18524
rect 44584 18468 44588 18524
rect 44524 18464 44588 18468
rect 58728 18524 58792 18528
rect 58728 18468 58732 18524
rect 58732 18468 58788 18524
rect 58788 18468 58792 18524
rect 58728 18464 58792 18468
rect 58808 18524 58872 18528
rect 58808 18468 58812 18524
rect 58812 18468 58868 18524
rect 58868 18468 58872 18524
rect 58808 18464 58872 18468
rect 58888 18524 58952 18528
rect 58888 18468 58892 18524
rect 58892 18468 58948 18524
rect 58948 18468 58952 18524
rect 58888 18464 58952 18468
rect 58968 18524 59032 18528
rect 58968 18468 58972 18524
rect 58972 18468 59028 18524
rect 59028 18468 59032 18524
rect 58968 18464 59032 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 22618 17980 22682 17984
rect 22618 17924 22622 17980
rect 22622 17924 22678 17980
rect 22678 17924 22682 17980
rect 22618 17920 22682 17924
rect 22698 17980 22762 17984
rect 22698 17924 22702 17980
rect 22702 17924 22758 17980
rect 22758 17924 22762 17980
rect 22698 17920 22762 17924
rect 22778 17980 22842 17984
rect 22778 17924 22782 17980
rect 22782 17924 22838 17980
rect 22838 17924 22842 17980
rect 22778 17920 22842 17924
rect 22858 17980 22922 17984
rect 22858 17924 22862 17980
rect 22862 17924 22918 17980
rect 22918 17924 22922 17980
rect 22858 17920 22922 17924
rect 37062 17980 37126 17984
rect 37062 17924 37066 17980
rect 37066 17924 37122 17980
rect 37122 17924 37126 17980
rect 37062 17920 37126 17924
rect 37142 17980 37206 17984
rect 37142 17924 37146 17980
rect 37146 17924 37202 17980
rect 37202 17924 37206 17980
rect 37142 17920 37206 17924
rect 37222 17980 37286 17984
rect 37222 17924 37226 17980
rect 37226 17924 37282 17980
rect 37282 17924 37286 17980
rect 37222 17920 37286 17924
rect 37302 17980 37366 17984
rect 37302 17924 37306 17980
rect 37306 17924 37362 17980
rect 37362 17924 37366 17980
rect 37302 17920 37366 17924
rect 51506 17980 51570 17984
rect 51506 17924 51510 17980
rect 51510 17924 51566 17980
rect 51566 17924 51570 17980
rect 51506 17920 51570 17924
rect 51586 17980 51650 17984
rect 51586 17924 51590 17980
rect 51590 17924 51646 17980
rect 51646 17924 51650 17980
rect 51586 17920 51650 17924
rect 51666 17980 51730 17984
rect 51666 17924 51670 17980
rect 51670 17924 51726 17980
rect 51726 17924 51730 17980
rect 51666 17920 51730 17924
rect 51746 17980 51810 17984
rect 51746 17924 51750 17980
rect 51750 17924 51806 17980
rect 51806 17924 51810 17980
rect 51746 17920 51810 17924
rect 15396 17436 15460 17440
rect 15396 17380 15400 17436
rect 15400 17380 15456 17436
rect 15456 17380 15460 17436
rect 15396 17376 15460 17380
rect 15476 17436 15540 17440
rect 15476 17380 15480 17436
rect 15480 17380 15536 17436
rect 15536 17380 15540 17436
rect 15476 17376 15540 17380
rect 15556 17436 15620 17440
rect 15556 17380 15560 17436
rect 15560 17380 15616 17436
rect 15616 17380 15620 17436
rect 15556 17376 15620 17380
rect 15636 17436 15700 17440
rect 15636 17380 15640 17436
rect 15640 17380 15696 17436
rect 15696 17380 15700 17436
rect 15636 17376 15700 17380
rect 29840 17436 29904 17440
rect 29840 17380 29844 17436
rect 29844 17380 29900 17436
rect 29900 17380 29904 17436
rect 29840 17376 29904 17380
rect 29920 17436 29984 17440
rect 29920 17380 29924 17436
rect 29924 17380 29980 17436
rect 29980 17380 29984 17436
rect 29920 17376 29984 17380
rect 30000 17436 30064 17440
rect 30000 17380 30004 17436
rect 30004 17380 30060 17436
rect 30060 17380 30064 17436
rect 30000 17376 30064 17380
rect 30080 17436 30144 17440
rect 30080 17380 30084 17436
rect 30084 17380 30140 17436
rect 30140 17380 30144 17436
rect 30080 17376 30144 17380
rect 44284 17436 44348 17440
rect 44284 17380 44288 17436
rect 44288 17380 44344 17436
rect 44344 17380 44348 17436
rect 44284 17376 44348 17380
rect 44364 17436 44428 17440
rect 44364 17380 44368 17436
rect 44368 17380 44424 17436
rect 44424 17380 44428 17436
rect 44364 17376 44428 17380
rect 44444 17436 44508 17440
rect 44444 17380 44448 17436
rect 44448 17380 44504 17436
rect 44504 17380 44508 17436
rect 44444 17376 44508 17380
rect 44524 17436 44588 17440
rect 44524 17380 44528 17436
rect 44528 17380 44584 17436
rect 44584 17380 44588 17436
rect 44524 17376 44588 17380
rect 58728 17436 58792 17440
rect 58728 17380 58732 17436
rect 58732 17380 58788 17436
rect 58788 17380 58792 17436
rect 58728 17376 58792 17380
rect 58808 17436 58872 17440
rect 58808 17380 58812 17436
rect 58812 17380 58868 17436
rect 58868 17380 58872 17436
rect 58808 17376 58872 17380
rect 58888 17436 58952 17440
rect 58888 17380 58892 17436
rect 58892 17380 58948 17436
rect 58948 17380 58952 17436
rect 58888 17376 58952 17380
rect 58968 17436 59032 17440
rect 58968 17380 58972 17436
rect 58972 17380 59028 17436
rect 59028 17380 59032 17436
rect 58968 17376 59032 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 22618 16892 22682 16896
rect 22618 16836 22622 16892
rect 22622 16836 22678 16892
rect 22678 16836 22682 16892
rect 22618 16832 22682 16836
rect 22698 16892 22762 16896
rect 22698 16836 22702 16892
rect 22702 16836 22758 16892
rect 22758 16836 22762 16892
rect 22698 16832 22762 16836
rect 22778 16892 22842 16896
rect 22778 16836 22782 16892
rect 22782 16836 22838 16892
rect 22838 16836 22842 16892
rect 22778 16832 22842 16836
rect 22858 16892 22922 16896
rect 22858 16836 22862 16892
rect 22862 16836 22918 16892
rect 22918 16836 22922 16892
rect 22858 16832 22922 16836
rect 37062 16892 37126 16896
rect 37062 16836 37066 16892
rect 37066 16836 37122 16892
rect 37122 16836 37126 16892
rect 37062 16832 37126 16836
rect 37142 16892 37206 16896
rect 37142 16836 37146 16892
rect 37146 16836 37202 16892
rect 37202 16836 37206 16892
rect 37142 16832 37206 16836
rect 37222 16892 37286 16896
rect 37222 16836 37226 16892
rect 37226 16836 37282 16892
rect 37282 16836 37286 16892
rect 37222 16832 37286 16836
rect 37302 16892 37366 16896
rect 37302 16836 37306 16892
rect 37306 16836 37362 16892
rect 37362 16836 37366 16892
rect 37302 16832 37366 16836
rect 51506 16892 51570 16896
rect 51506 16836 51510 16892
rect 51510 16836 51566 16892
rect 51566 16836 51570 16892
rect 51506 16832 51570 16836
rect 51586 16892 51650 16896
rect 51586 16836 51590 16892
rect 51590 16836 51646 16892
rect 51646 16836 51650 16892
rect 51586 16832 51650 16836
rect 51666 16892 51730 16896
rect 51666 16836 51670 16892
rect 51670 16836 51726 16892
rect 51726 16836 51730 16892
rect 51666 16832 51730 16836
rect 51746 16892 51810 16896
rect 51746 16836 51750 16892
rect 51750 16836 51806 16892
rect 51806 16836 51810 16892
rect 51746 16832 51810 16836
rect 9812 16688 9876 16692
rect 9812 16632 9826 16688
rect 9826 16632 9876 16688
rect 9812 16628 9876 16632
rect 34284 16688 34348 16692
rect 34284 16632 34298 16688
rect 34298 16632 34348 16688
rect 34284 16628 34348 16632
rect 15396 16348 15460 16352
rect 15396 16292 15400 16348
rect 15400 16292 15456 16348
rect 15456 16292 15460 16348
rect 15396 16288 15460 16292
rect 15476 16348 15540 16352
rect 15476 16292 15480 16348
rect 15480 16292 15536 16348
rect 15536 16292 15540 16348
rect 15476 16288 15540 16292
rect 15556 16348 15620 16352
rect 15556 16292 15560 16348
rect 15560 16292 15616 16348
rect 15616 16292 15620 16348
rect 15556 16288 15620 16292
rect 15636 16348 15700 16352
rect 15636 16292 15640 16348
rect 15640 16292 15696 16348
rect 15696 16292 15700 16348
rect 15636 16288 15700 16292
rect 29840 16348 29904 16352
rect 29840 16292 29844 16348
rect 29844 16292 29900 16348
rect 29900 16292 29904 16348
rect 29840 16288 29904 16292
rect 29920 16348 29984 16352
rect 29920 16292 29924 16348
rect 29924 16292 29980 16348
rect 29980 16292 29984 16348
rect 29920 16288 29984 16292
rect 30000 16348 30064 16352
rect 30000 16292 30004 16348
rect 30004 16292 30060 16348
rect 30060 16292 30064 16348
rect 30000 16288 30064 16292
rect 30080 16348 30144 16352
rect 30080 16292 30084 16348
rect 30084 16292 30140 16348
rect 30140 16292 30144 16348
rect 30080 16288 30144 16292
rect 44284 16348 44348 16352
rect 44284 16292 44288 16348
rect 44288 16292 44344 16348
rect 44344 16292 44348 16348
rect 44284 16288 44348 16292
rect 44364 16348 44428 16352
rect 44364 16292 44368 16348
rect 44368 16292 44424 16348
rect 44424 16292 44428 16348
rect 44364 16288 44428 16292
rect 44444 16348 44508 16352
rect 44444 16292 44448 16348
rect 44448 16292 44504 16348
rect 44504 16292 44508 16348
rect 44444 16288 44508 16292
rect 44524 16348 44588 16352
rect 44524 16292 44528 16348
rect 44528 16292 44584 16348
rect 44584 16292 44588 16348
rect 44524 16288 44588 16292
rect 58728 16348 58792 16352
rect 58728 16292 58732 16348
rect 58732 16292 58788 16348
rect 58788 16292 58792 16348
rect 58728 16288 58792 16292
rect 58808 16348 58872 16352
rect 58808 16292 58812 16348
rect 58812 16292 58868 16348
rect 58868 16292 58872 16348
rect 58808 16288 58872 16292
rect 58888 16348 58952 16352
rect 58888 16292 58892 16348
rect 58892 16292 58948 16348
rect 58948 16292 58952 16348
rect 58888 16288 58952 16292
rect 58968 16348 59032 16352
rect 58968 16292 58972 16348
rect 58972 16292 59028 16348
rect 59028 16292 59032 16348
rect 58968 16288 59032 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 22618 15804 22682 15808
rect 22618 15748 22622 15804
rect 22622 15748 22678 15804
rect 22678 15748 22682 15804
rect 22618 15744 22682 15748
rect 22698 15804 22762 15808
rect 22698 15748 22702 15804
rect 22702 15748 22758 15804
rect 22758 15748 22762 15804
rect 22698 15744 22762 15748
rect 22778 15804 22842 15808
rect 22778 15748 22782 15804
rect 22782 15748 22838 15804
rect 22838 15748 22842 15804
rect 22778 15744 22842 15748
rect 22858 15804 22922 15808
rect 22858 15748 22862 15804
rect 22862 15748 22918 15804
rect 22918 15748 22922 15804
rect 22858 15744 22922 15748
rect 37062 15804 37126 15808
rect 37062 15748 37066 15804
rect 37066 15748 37122 15804
rect 37122 15748 37126 15804
rect 37062 15744 37126 15748
rect 37142 15804 37206 15808
rect 37142 15748 37146 15804
rect 37146 15748 37202 15804
rect 37202 15748 37206 15804
rect 37142 15744 37206 15748
rect 37222 15804 37286 15808
rect 37222 15748 37226 15804
rect 37226 15748 37282 15804
rect 37282 15748 37286 15804
rect 37222 15744 37286 15748
rect 37302 15804 37366 15808
rect 37302 15748 37306 15804
rect 37306 15748 37362 15804
rect 37362 15748 37366 15804
rect 37302 15744 37366 15748
rect 51506 15804 51570 15808
rect 51506 15748 51510 15804
rect 51510 15748 51566 15804
rect 51566 15748 51570 15804
rect 51506 15744 51570 15748
rect 51586 15804 51650 15808
rect 51586 15748 51590 15804
rect 51590 15748 51646 15804
rect 51646 15748 51650 15804
rect 51586 15744 51650 15748
rect 51666 15804 51730 15808
rect 51666 15748 51670 15804
rect 51670 15748 51726 15804
rect 51726 15748 51730 15804
rect 51666 15744 51730 15748
rect 51746 15804 51810 15808
rect 51746 15748 51750 15804
rect 51750 15748 51806 15804
rect 51806 15748 51810 15804
rect 51746 15744 51810 15748
rect 15396 15260 15460 15264
rect 15396 15204 15400 15260
rect 15400 15204 15456 15260
rect 15456 15204 15460 15260
rect 15396 15200 15460 15204
rect 15476 15260 15540 15264
rect 15476 15204 15480 15260
rect 15480 15204 15536 15260
rect 15536 15204 15540 15260
rect 15476 15200 15540 15204
rect 15556 15260 15620 15264
rect 15556 15204 15560 15260
rect 15560 15204 15616 15260
rect 15616 15204 15620 15260
rect 15556 15200 15620 15204
rect 15636 15260 15700 15264
rect 15636 15204 15640 15260
rect 15640 15204 15696 15260
rect 15696 15204 15700 15260
rect 15636 15200 15700 15204
rect 29840 15260 29904 15264
rect 29840 15204 29844 15260
rect 29844 15204 29900 15260
rect 29900 15204 29904 15260
rect 29840 15200 29904 15204
rect 29920 15260 29984 15264
rect 29920 15204 29924 15260
rect 29924 15204 29980 15260
rect 29980 15204 29984 15260
rect 29920 15200 29984 15204
rect 30000 15260 30064 15264
rect 30000 15204 30004 15260
rect 30004 15204 30060 15260
rect 30060 15204 30064 15260
rect 30000 15200 30064 15204
rect 30080 15260 30144 15264
rect 30080 15204 30084 15260
rect 30084 15204 30140 15260
rect 30140 15204 30144 15260
rect 30080 15200 30144 15204
rect 44284 15260 44348 15264
rect 44284 15204 44288 15260
rect 44288 15204 44344 15260
rect 44344 15204 44348 15260
rect 44284 15200 44348 15204
rect 44364 15260 44428 15264
rect 44364 15204 44368 15260
rect 44368 15204 44424 15260
rect 44424 15204 44428 15260
rect 44364 15200 44428 15204
rect 44444 15260 44508 15264
rect 44444 15204 44448 15260
rect 44448 15204 44504 15260
rect 44504 15204 44508 15260
rect 44444 15200 44508 15204
rect 44524 15260 44588 15264
rect 44524 15204 44528 15260
rect 44528 15204 44584 15260
rect 44584 15204 44588 15260
rect 44524 15200 44588 15204
rect 58728 15260 58792 15264
rect 58728 15204 58732 15260
rect 58732 15204 58788 15260
rect 58788 15204 58792 15260
rect 58728 15200 58792 15204
rect 58808 15260 58872 15264
rect 58808 15204 58812 15260
rect 58812 15204 58868 15260
rect 58868 15204 58872 15260
rect 58808 15200 58872 15204
rect 58888 15260 58952 15264
rect 58888 15204 58892 15260
rect 58892 15204 58948 15260
rect 58948 15204 58952 15260
rect 58888 15200 58952 15204
rect 58968 15260 59032 15264
rect 58968 15204 58972 15260
rect 58972 15204 59028 15260
rect 59028 15204 59032 15260
rect 58968 15200 59032 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 22618 14716 22682 14720
rect 22618 14660 22622 14716
rect 22622 14660 22678 14716
rect 22678 14660 22682 14716
rect 22618 14656 22682 14660
rect 22698 14716 22762 14720
rect 22698 14660 22702 14716
rect 22702 14660 22758 14716
rect 22758 14660 22762 14716
rect 22698 14656 22762 14660
rect 22778 14716 22842 14720
rect 22778 14660 22782 14716
rect 22782 14660 22838 14716
rect 22838 14660 22842 14716
rect 22778 14656 22842 14660
rect 22858 14716 22922 14720
rect 22858 14660 22862 14716
rect 22862 14660 22918 14716
rect 22918 14660 22922 14716
rect 22858 14656 22922 14660
rect 37062 14716 37126 14720
rect 37062 14660 37066 14716
rect 37066 14660 37122 14716
rect 37122 14660 37126 14716
rect 37062 14656 37126 14660
rect 37142 14716 37206 14720
rect 37142 14660 37146 14716
rect 37146 14660 37202 14716
rect 37202 14660 37206 14716
rect 37142 14656 37206 14660
rect 37222 14716 37286 14720
rect 37222 14660 37226 14716
rect 37226 14660 37282 14716
rect 37282 14660 37286 14716
rect 37222 14656 37286 14660
rect 37302 14716 37366 14720
rect 37302 14660 37306 14716
rect 37306 14660 37362 14716
rect 37362 14660 37366 14716
rect 37302 14656 37366 14660
rect 51506 14716 51570 14720
rect 51506 14660 51510 14716
rect 51510 14660 51566 14716
rect 51566 14660 51570 14716
rect 51506 14656 51570 14660
rect 51586 14716 51650 14720
rect 51586 14660 51590 14716
rect 51590 14660 51646 14716
rect 51646 14660 51650 14716
rect 51586 14656 51650 14660
rect 51666 14716 51730 14720
rect 51666 14660 51670 14716
rect 51670 14660 51726 14716
rect 51726 14660 51730 14716
rect 51666 14656 51730 14660
rect 51746 14716 51810 14720
rect 51746 14660 51750 14716
rect 51750 14660 51806 14716
rect 51806 14660 51810 14716
rect 51746 14656 51810 14660
rect 15396 14172 15460 14176
rect 15396 14116 15400 14172
rect 15400 14116 15456 14172
rect 15456 14116 15460 14172
rect 15396 14112 15460 14116
rect 15476 14172 15540 14176
rect 15476 14116 15480 14172
rect 15480 14116 15536 14172
rect 15536 14116 15540 14172
rect 15476 14112 15540 14116
rect 15556 14172 15620 14176
rect 15556 14116 15560 14172
rect 15560 14116 15616 14172
rect 15616 14116 15620 14172
rect 15556 14112 15620 14116
rect 15636 14172 15700 14176
rect 15636 14116 15640 14172
rect 15640 14116 15696 14172
rect 15696 14116 15700 14172
rect 15636 14112 15700 14116
rect 29840 14172 29904 14176
rect 29840 14116 29844 14172
rect 29844 14116 29900 14172
rect 29900 14116 29904 14172
rect 29840 14112 29904 14116
rect 29920 14172 29984 14176
rect 29920 14116 29924 14172
rect 29924 14116 29980 14172
rect 29980 14116 29984 14172
rect 29920 14112 29984 14116
rect 30000 14172 30064 14176
rect 30000 14116 30004 14172
rect 30004 14116 30060 14172
rect 30060 14116 30064 14172
rect 30000 14112 30064 14116
rect 30080 14172 30144 14176
rect 30080 14116 30084 14172
rect 30084 14116 30140 14172
rect 30140 14116 30144 14172
rect 30080 14112 30144 14116
rect 44284 14172 44348 14176
rect 44284 14116 44288 14172
rect 44288 14116 44344 14172
rect 44344 14116 44348 14172
rect 44284 14112 44348 14116
rect 44364 14172 44428 14176
rect 44364 14116 44368 14172
rect 44368 14116 44424 14172
rect 44424 14116 44428 14172
rect 44364 14112 44428 14116
rect 44444 14172 44508 14176
rect 44444 14116 44448 14172
rect 44448 14116 44504 14172
rect 44504 14116 44508 14172
rect 44444 14112 44508 14116
rect 44524 14172 44588 14176
rect 44524 14116 44528 14172
rect 44528 14116 44584 14172
rect 44584 14116 44588 14172
rect 44524 14112 44588 14116
rect 58728 14172 58792 14176
rect 58728 14116 58732 14172
rect 58732 14116 58788 14172
rect 58788 14116 58792 14172
rect 58728 14112 58792 14116
rect 58808 14172 58872 14176
rect 58808 14116 58812 14172
rect 58812 14116 58868 14172
rect 58868 14116 58872 14172
rect 58808 14112 58872 14116
rect 58888 14172 58952 14176
rect 58888 14116 58892 14172
rect 58892 14116 58948 14172
rect 58948 14116 58952 14172
rect 58888 14112 58952 14116
rect 58968 14172 59032 14176
rect 58968 14116 58972 14172
rect 58972 14116 59028 14172
rect 59028 14116 59032 14172
rect 58968 14112 59032 14116
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 22618 13628 22682 13632
rect 22618 13572 22622 13628
rect 22622 13572 22678 13628
rect 22678 13572 22682 13628
rect 22618 13568 22682 13572
rect 22698 13628 22762 13632
rect 22698 13572 22702 13628
rect 22702 13572 22758 13628
rect 22758 13572 22762 13628
rect 22698 13568 22762 13572
rect 22778 13628 22842 13632
rect 22778 13572 22782 13628
rect 22782 13572 22838 13628
rect 22838 13572 22842 13628
rect 22778 13568 22842 13572
rect 22858 13628 22922 13632
rect 22858 13572 22862 13628
rect 22862 13572 22918 13628
rect 22918 13572 22922 13628
rect 22858 13568 22922 13572
rect 37062 13628 37126 13632
rect 37062 13572 37066 13628
rect 37066 13572 37122 13628
rect 37122 13572 37126 13628
rect 37062 13568 37126 13572
rect 37142 13628 37206 13632
rect 37142 13572 37146 13628
rect 37146 13572 37202 13628
rect 37202 13572 37206 13628
rect 37142 13568 37206 13572
rect 37222 13628 37286 13632
rect 37222 13572 37226 13628
rect 37226 13572 37282 13628
rect 37282 13572 37286 13628
rect 37222 13568 37286 13572
rect 37302 13628 37366 13632
rect 37302 13572 37306 13628
rect 37306 13572 37362 13628
rect 37362 13572 37366 13628
rect 37302 13568 37366 13572
rect 51506 13628 51570 13632
rect 51506 13572 51510 13628
rect 51510 13572 51566 13628
rect 51566 13572 51570 13628
rect 51506 13568 51570 13572
rect 51586 13628 51650 13632
rect 51586 13572 51590 13628
rect 51590 13572 51646 13628
rect 51646 13572 51650 13628
rect 51586 13568 51650 13572
rect 51666 13628 51730 13632
rect 51666 13572 51670 13628
rect 51670 13572 51726 13628
rect 51726 13572 51730 13628
rect 51666 13568 51730 13572
rect 51746 13628 51810 13632
rect 51746 13572 51750 13628
rect 51750 13572 51806 13628
rect 51806 13572 51810 13628
rect 51746 13568 51810 13572
rect 15396 13084 15460 13088
rect 15396 13028 15400 13084
rect 15400 13028 15456 13084
rect 15456 13028 15460 13084
rect 15396 13024 15460 13028
rect 15476 13084 15540 13088
rect 15476 13028 15480 13084
rect 15480 13028 15536 13084
rect 15536 13028 15540 13084
rect 15476 13024 15540 13028
rect 15556 13084 15620 13088
rect 15556 13028 15560 13084
rect 15560 13028 15616 13084
rect 15616 13028 15620 13084
rect 15556 13024 15620 13028
rect 15636 13084 15700 13088
rect 15636 13028 15640 13084
rect 15640 13028 15696 13084
rect 15696 13028 15700 13084
rect 15636 13024 15700 13028
rect 29840 13084 29904 13088
rect 29840 13028 29844 13084
rect 29844 13028 29900 13084
rect 29900 13028 29904 13084
rect 29840 13024 29904 13028
rect 29920 13084 29984 13088
rect 29920 13028 29924 13084
rect 29924 13028 29980 13084
rect 29980 13028 29984 13084
rect 29920 13024 29984 13028
rect 30000 13084 30064 13088
rect 30000 13028 30004 13084
rect 30004 13028 30060 13084
rect 30060 13028 30064 13084
rect 30000 13024 30064 13028
rect 30080 13084 30144 13088
rect 30080 13028 30084 13084
rect 30084 13028 30140 13084
rect 30140 13028 30144 13084
rect 30080 13024 30144 13028
rect 44284 13084 44348 13088
rect 44284 13028 44288 13084
rect 44288 13028 44344 13084
rect 44344 13028 44348 13084
rect 44284 13024 44348 13028
rect 44364 13084 44428 13088
rect 44364 13028 44368 13084
rect 44368 13028 44424 13084
rect 44424 13028 44428 13084
rect 44364 13024 44428 13028
rect 44444 13084 44508 13088
rect 44444 13028 44448 13084
rect 44448 13028 44504 13084
rect 44504 13028 44508 13084
rect 44444 13024 44508 13028
rect 44524 13084 44588 13088
rect 44524 13028 44528 13084
rect 44528 13028 44584 13084
rect 44584 13028 44588 13084
rect 44524 13024 44588 13028
rect 58728 13084 58792 13088
rect 58728 13028 58732 13084
rect 58732 13028 58788 13084
rect 58788 13028 58792 13084
rect 58728 13024 58792 13028
rect 58808 13084 58872 13088
rect 58808 13028 58812 13084
rect 58812 13028 58868 13084
rect 58868 13028 58872 13084
rect 58808 13024 58872 13028
rect 58888 13084 58952 13088
rect 58888 13028 58892 13084
rect 58892 13028 58948 13084
rect 58948 13028 58952 13084
rect 58888 13024 58952 13028
rect 58968 13084 59032 13088
rect 58968 13028 58972 13084
rect 58972 13028 59028 13084
rect 59028 13028 59032 13084
rect 58968 13024 59032 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 22618 12540 22682 12544
rect 22618 12484 22622 12540
rect 22622 12484 22678 12540
rect 22678 12484 22682 12540
rect 22618 12480 22682 12484
rect 22698 12540 22762 12544
rect 22698 12484 22702 12540
rect 22702 12484 22758 12540
rect 22758 12484 22762 12540
rect 22698 12480 22762 12484
rect 22778 12540 22842 12544
rect 22778 12484 22782 12540
rect 22782 12484 22838 12540
rect 22838 12484 22842 12540
rect 22778 12480 22842 12484
rect 22858 12540 22922 12544
rect 22858 12484 22862 12540
rect 22862 12484 22918 12540
rect 22918 12484 22922 12540
rect 22858 12480 22922 12484
rect 37062 12540 37126 12544
rect 37062 12484 37066 12540
rect 37066 12484 37122 12540
rect 37122 12484 37126 12540
rect 37062 12480 37126 12484
rect 37142 12540 37206 12544
rect 37142 12484 37146 12540
rect 37146 12484 37202 12540
rect 37202 12484 37206 12540
rect 37142 12480 37206 12484
rect 37222 12540 37286 12544
rect 37222 12484 37226 12540
rect 37226 12484 37282 12540
rect 37282 12484 37286 12540
rect 37222 12480 37286 12484
rect 37302 12540 37366 12544
rect 37302 12484 37306 12540
rect 37306 12484 37362 12540
rect 37362 12484 37366 12540
rect 37302 12480 37366 12484
rect 51506 12540 51570 12544
rect 51506 12484 51510 12540
rect 51510 12484 51566 12540
rect 51566 12484 51570 12540
rect 51506 12480 51570 12484
rect 51586 12540 51650 12544
rect 51586 12484 51590 12540
rect 51590 12484 51646 12540
rect 51646 12484 51650 12540
rect 51586 12480 51650 12484
rect 51666 12540 51730 12544
rect 51666 12484 51670 12540
rect 51670 12484 51726 12540
rect 51726 12484 51730 12540
rect 51666 12480 51730 12484
rect 51746 12540 51810 12544
rect 51746 12484 51750 12540
rect 51750 12484 51806 12540
rect 51806 12484 51810 12540
rect 51746 12480 51810 12484
rect 15396 11996 15460 12000
rect 15396 11940 15400 11996
rect 15400 11940 15456 11996
rect 15456 11940 15460 11996
rect 15396 11936 15460 11940
rect 15476 11996 15540 12000
rect 15476 11940 15480 11996
rect 15480 11940 15536 11996
rect 15536 11940 15540 11996
rect 15476 11936 15540 11940
rect 15556 11996 15620 12000
rect 15556 11940 15560 11996
rect 15560 11940 15616 11996
rect 15616 11940 15620 11996
rect 15556 11936 15620 11940
rect 15636 11996 15700 12000
rect 15636 11940 15640 11996
rect 15640 11940 15696 11996
rect 15696 11940 15700 11996
rect 15636 11936 15700 11940
rect 29840 11996 29904 12000
rect 29840 11940 29844 11996
rect 29844 11940 29900 11996
rect 29900 11940 29904 11996
rect 29840 11936 29904 11940
rect 29920 11996 29984 12000
rect 29920 11940 29924 11996
rect 29924 11940 29980 11996
rect 29980 11940 29984 11996
rect 29920 11936 29984 11940
rect 30000 11996 30064 12000
rect 30000 11940 30004 11996
rect 30004 11940 30060 11996
rect 30060 11940 30064 11996
rect 30000 11936 30064 11940
rect 30080 11996 30144 12000
rect 30080 11940 30084 11996
rect 30084 11940 30140 11996
rect 30140 11940 30144 11996
rect 30080 11936 30144 11940
rect 44284 11996 44348 12000
rect 44284 11940 44288 11996
rect 44288 11940 44344 11996
rect 44344 11940 44348 11996
rect 44284 11936 44348 11940
rect 44364 11996 44428 12000
rect 44364 11940 44368 11996
rect 44368 11940 44424 11996
rect 44424 11940 44428 11996
rect 44364 11936 44428 11940
rect 44444 11996 44508 12000
rect 44444 11940 44448 11996
rect 44448 11940 44504 11996
rect 44504 11940 44508 11996
rect 44444 11936 44508 11940
rect 44524 11996 44588 12000
rect 44524 11940 44528 11996
rect 44528 11940 44584 11996
rect 44584 11940 44588 11996
rect 44524 11936 44588 11940
rect 58728 11996 58792 12000
rect 58728 11940 58732 11996
rect 58732 11940 58788 11996
rect 58788 11940 58792 11996
rect 58728 11936 58792 11940
rect 58808 11996 58872 12000
rect 58808 11940 58812 11996
rect 58812 11940 58868 11996
rect 58868 11940 58872 11996
rect 58808 11936 58872 11940
rect 58888 11996 58952 12000
rect 58888 11940 58892 11996
rect 58892 11940 58948 11996
rect 58948 11940 58952 11996
rect 58888 11936 58952 11940
rect 58968 11996 59032 12000
rect 58968 11940 58972 11996
rect 58972 11940 59028 11996
rect 59028 11940 59032 11996
rect 58968 11936 59032 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 22618 11452 22682 11456
rect 22618 11396 22622 11452
rect 22622 11396 22678 11452
rect 22678 11396 22682 11452
rect 22618 11392 22682 11396
rect 22698 11452 22762 11456
rect 22698 11396 22702 11452
rect 22702 11396 22758 11452
rect 22758 11396 22762 11452
rect 22698 11392 22762 11396
rect 22778 11452 22842 11456
rect 22778 11396 22782 11452
rect 22782 11396 22838 11452
rect 22838 11396 22842 11452
rect 22778 11392 22842 11396
rect 22858 11452 22922 11456
rect 22858 11396 22862 11452
rect 22862 11396 22918 11452
rect 22918 11396 22922 11452
rect 22858 11392 22922 11396
rect 37062 11452 37126 11456
rect 37062 11396 37066 11452
rect 37066 11396 37122 11452
rect 37122 11396 37126 11452
rect 37062 11392 37126 11396
rect 37142 11452 37206 11456
rect 37142 11396 37146 11452
rect 37146 11396 37202 11452
rect 37202 11396 37206 11452
rect 37142 11392 37206 11396
rect 37222 11452 37286 11456
rect 37222 11396 37226 11452
rect 37226 11396 37282 11452
rect 37282 11396 37286 11452
rect 37222 11392 37286 11396
rect 37302 11452 37366 11456
rect 37302 11396 37306 11452
rect 37306 11396 37362 11452
rect 37362 11396 37366 11452
rect 37302 11392 37366 11396
rect 51506 11452 51570 11456
rect 51506 11396 51510 11452
rect 51510 11396 51566 11452
rect 51566 11396 51570 11452
rect 51506 11392 51570 11396
rect 51586 11452 51650 11456
rect 51586 11396 51590 11452
rect 51590 11396 51646 11452
rect 51646 11396 51650 11452
rect 51586 11392 51650 11396
rect 51666 11452 51730 11456
rect 51666 11396 51670 11452
rect 51670 11396 51726 11452
rect 51726 11396 51730 11452
rect 51666 11392 51730 11396
rect 51746 11452 51810 11456
rect 51746 11396 51750 11452
rect 51750 11396 51806 11452
rect 51806 11396 51810 11452
rect 51746 11392 51810 11396
rect 10548 11052 10612 11116
rect 37596 11052 37660 11116
rect 15396 10908 15460 10912
rect 15396 10852 15400 10908
rect 15400 10852 15456 10908
rect 15456 10852 15460 10908
rect 15396 10848 15460 10852
rect 15476 10908 15540 10912
rect 15476 10852 15480 10908
rect 15480 10852 15536 10908
rect 15536 10852 15540 10908
rect 15476 10848 15540 10852
rect 15556 10908 15620 10912
rect 15556 10852 15560 10908
rect 15560 10852 15616 10908
rect 15616 10852 15620 10908
rect 15556 10848 15620 10852
rect 15636 10908 15700 10912
rect 15636 10852 15640 10908
rect 15640 10852 15696 10908
rect 15696 10852 15700 10908
rect 15636 10848 15700 10852
rect 29840 10908 29904 10912
rect 29840 10852 29844 10908
rect 29844 10852 29900 10908
rect 29900 10852 29904 10908
rect 29840 10848 29904 10852
rect 29920 10908 29984 10912
rect 29920 10852 29924 10908
rect 29924 10852 29980 10908
rect 29980 10852 29984 10908
rect 29920 10848 29984 10852
rect 30000 10908 30064 10912
rect 30000 10852 30004 10908
rect 30004 10852 30060 10908
rect 30060 10852 30064 10908
rect 30000 10848 30064 10852
rect 30080 10908 30144 10912
rect 30080 10852 30084 10908
rect 30084 10852 30140 10908
rect 30140 10852 30144 10908
rect 30080 10848 30144 10852
rect 44284 10908 44348 10912
rect 44284 10852 44288 10908
rect 44288 10852 44344 10908
rect 44344 10852 44348 10908
rect 44284 10848 44348 10852
rect 44364 10908 44428 10912
rect 44364 10852 44368 10908
rect 44368 10852 44424 10908
rect 44424 10852 44428 10908
rect 44364 10848 44428 10852
rect 44444 10908 44508 10912
rect 44444 10852 44448 10908
rect 44448 10852 44504 10908
rect 44504 10852 44508 10908
rect 44444 10848 44508 10852
rect 44524 10908 44588 10912
rect 44524 10852 44528 10908
rect 44528 10852 44584 10908
rect 44584 10852 44588 10908
rect 44524 10848 44588 10852
rect 58728 10908 58792 10912
rect 58728 10852 58732 10908
rect 58732 10852 58788 10908
rect 58788 10852 58792 10908
rect 58728 10848 58792 10852
rect 58808 10908 58872 10912
rect 58808 10852 58812 10908
rect 58812 10852 58868 10908
rect 58868 10852 58872 10908
rect 58808 10848 58872 10852
rect 58888 10908 58952 10912
rect 58888 10852 58892 10908
rect 58892 10852 58948 10908
rect 58948 10852 58952 10908
rect 58888 10848 58952 10852
rect 58968 10908 59032 10912
rect 58968 10852 58972 10908
rect 58972 10852 59028 10908
rect 59028 10852 59032 10908
rect 58968 10848 59032 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 22618 10364 22682 10368
rect 22618 10308 22622 10364
rect 22622 10308 22678 10364
rect 22678 10308 22682 10364
rect 22618 10304 22682 10308
rect 22698 10364 22762 10368
rect 22698 10308 22702 10364
rect 22702 10308 22758 10364
rect 22758 10308 22762 10364
rect 22698 10304 22762 10308
rect 22778 10364 22842 10368
rect 22778 10308 22782 10364
rect 22782 10308 22838 10364
rect 22838 10308 22842 10364
rect 22778 10304 22842 10308
rect 22858 10364 22922 10368
rect 22858 10308 22862 10364
rect 22862 10308 22918 10364
rect 22918 10308 22922 10364
rect 22858 10304 22922 10308
rect 37062 10364 37126 10368
rect 37062 10308 37066 10364
rect 37066 10308 37122 10364
rect 37122 10308 37126 10364
rect 37062 10304 37126 10308
rect 37142 10364 37206 10368
rect 37142 10308 37146 10364
rect 37146 10308 37202 10364
rect 37202 10308 37206 10364
rect 37142 10304 37206 10308
rect 37222 10364 37286 10368
rect 37222 10308 37226 10364
rect 37226 10308 37282 10364
rect 37282 10308 37286 10364
rect 37222 10304 37286 10308
rect 37302 10364 37366 10368
rect 37302 10308 37306 10364
rect 37306 10308 37362 10364
rect 37362 10308 37366 10364
rect 37302 10304 37366 10308
rect 51506 10364 51570 10368
rect 51506 10308 51510 10364
rect 51510 10308 51566 10364
rect 51566 10308 51570 10364
rect 51506 10304 51570 10308
rect 51586 10364 51650 10368
rect 51586 10308 51590 10364
rect 51590 10308 51646 10364
rect 51646 10308 51650 10364
rect 51586 10304 51650 10308
rect 51666 10364 51730 10368
rect 51666 10308 51670 10364
rect 51670 10308 51726 10364
rect 51726 10308 51730 10364
rect 51666 10304 51730 10308
rect 51746 10364 51810 10368
rect 51746 10308 51750 10364
rect 51750 10308 51806 10364
rect 51806 10308 51810 10364
rect 51746 10304 51810 10308
rect 15396 9820 15460 9824
rect 15396 9764 15400 9820
rect 15400 9764 15456 9820
rect 15456 9764 15460 9820
rect 15396 9760 15460 9764
rect 15476 9820 15540 9824
rect 15476 9764 15480 9820
rect 15480 9764 15536 9820
rect 15536 9764 15540 9820
rect 15476 9760 15540 9764
rect 15556 9820 15620 9824
rect 15556 9764 15560 9820
rect 15560 9764 15616 9820
rect 15616 9764 15620 9820
rect 15556 9760 15620 9764
rect 15636 9820 15700 9824
rect 15636 9764 15640 9820
rect 15640 9764 15696 9820
rect 15696 9764 15700 9820
rect 15636 9760 15700 9764
rect 29840 9820 29904 9824
rect 29840 9764 29844 9820
rect 29844 9764 29900 9820
rect 29900 9764 29904 9820
rect 29840 9760 29904 9764
rect 29920 9820 29984 9824
rect 29920 9764 29924 9820
rect 29924 9764 29980 9820
rect 29980 9764 29984 9820
rect 29920 9760 29984 9764
rect 30000 9820 30064 9824
rect 30000 9764 30004 9820
rect 30004 9764 30060 9820
rect 30060 9764 30064 9820
rect 30000 9760 30064 9764
rect 30080 9820 30144 9824
rect 30080 9764 30084 9820
rect 30084 9764 30140 9820
rect 30140 9764 30144 9820
rect 30080 9760 30144 9764
rect 44284 9820 44348 9824
rect 44284 9764 44288 9820
rect 44288 9764 44344 9820
rect 44344 9764 44348 9820
rect 44284 9760 44348 9764
rect 44364 9820 44428 9824
rect 44364 9764 44368 9820
rect 44368 9764 44424 9820
rect 44424 9764 44428 9820
rect 44364 9760 44428 9764
rect 44444 9820 44508 9824
rect 44444 9764 44448 9820
rect 44448 9764 44504 9820
rect 44504 9764 44508 9820
rect 44444 9760 44508 9764
rect 44524 9820 44588 9824
rect 44524 9764 44528 9820
rect 44528 9764 44584 9820
rect 44584 9764 44588 9820
rect 44524 9760 44588 9764
rect 58728 9820 58792 9824
rect 58728 9764 58732 9820
rect 58732 9764 58788 9820
rect 58788 9764 58792 9820
rect 58728 9760 58792 9764
rect 58808 9820 58872 9824
rect 58808 9764 58812 9820
rect 58812 9764 58868 9820
rect 58868 9764 58872 9820
rect 58808 9760 58872 9764
rect 58888 9820 58952 9824
rect 58888 9764 58892 9820
rect 58892 9764 58948 9820
rect 58948 9764 58952 9820
rect 58888 9760 58952 9764
rect 58968 9820 59032 9824
rect 58968 9764 58972 9820
rect 58972 9764 59028 9820
rect 59028 9764 59032 9820
rect 58968 9760 59032 9764
rect 34284 9556 34348 9620
rect 9812 9420 9876 9484
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 22618 9276 22682 9280
rect 22618 9220 22622 9276
rect 22622 9220 22678 9276
rect 22678 9220 22682 9276
rect 22618 9216 22682 9220
rect 22698 9276 22762 9280
rect 22698 9220 22702 9276
rect 22702 9220 22758 9276
rect 22758 9220 22762 9276
rect 22698 9216 22762 9220
rect 22778 9276 22842 9280
rect 22778 9220 22782 9276
rect 22782 9220 22838 9276
rect 22838 9220 22842 9276
rect 22778 9216 22842 9220
rect 22858 9276 22922 9280
rect 22858 9220 22862 9276
rect 22862 9220 22918 9276
rect 22918 9220 22922 9276
rect 22858 9216 22922 9220
rect 37062 9276 37126 9280
rect 37062 9220 37066 9276
rect 37066 9220 37122 9276
rect 37122 9220 37126 9276
rect 37062 9216 37126 9220
rect 37142 9276 37206 9280
rect 37142 9220 37146 9276
rect 37146 9220 37202 9276
rect 37202 9220 37206 9276
rect 37142 9216 37206 9220
rect 37222 9276 37286 9280
rect 37222 9220 37226 9276
rect 37226 9220 37282 9276
rect 37282 9220 37286 9276
rect 37222 9216 37286 9220
rect 37302 9276 37366 9280
rect 37302 9220 37306 9276
rect 37306 9220 37362 9276
rect 37362 9220 37366 9276
rect 37302 9216 37366 9220
rect 51506 9276 51570 9280
rect 51506 9220 51510 9276
rect 51510 9220 51566 9276
rect 51566 9220 51570 9276
rect 51506 9216 51570 9220
rect 51586 9276 51650 9280
rect 51586 9220 51590 9276
rect 51590 9220 51646 9276
rect 51646 9220 51650 9276
rect 51586 9216 51650 9220
rect 51666 9276 51730 9280
rect 51666 9220 51670 9276
rect 51670 9220 51726 9276
rect 51726 9220 51730 9276
rect 51666 9216 51730 9220
rect 51746 9276 51810 9280
rect 51746 9220 51750 9276
rect 51750 9220 51806 9276
rect 51806 9220 51810 9276
rect 51746 9216 51810 9220
rect 15396 8732 15460 8736
rect 15396 8676 15400 8732
rect 15400 8676 15456 8732
rect 15456 8676 15460 8732
rect 15396 8672 15460 8676
rect 15476 8732 15540 8736
rect 15476 8676 15480 8732
rect 15480 8676 15536 8732
rect 15536 8676 15540 8732
rect 15476 8672 15540 8676
rect 15556 8732 15620 8736
rect 15556 8676 15560 8732
rect 15560 8676 15616 8732
rect 15616 8676 15620 8732
rect 15556 8672 15620 8676
rect 15636 8732 15700 8736
rect 15636 8676 15640 8732
rect 15640 8676 15696 8732
rect 15696 8676 15700 8732
rect 15636 8672 15700 8676
rect 29840 8732 29904 8736
rect 29840 8676 29844 8732
rect 29844 8676 29900 8732
rect 29900 8676 29904 8732
rect 29840 8672 29904 8676
rect 29920 8732 29984 8736
rect 29920 8676 29924 8732
rect 29924 8676 29980 8732
rect 29980 8676 29984 8732
rect 29920 8672 29984 8676
rect 30000 8732 30064 8736
rect 30000 8676 30004 8732
rect 30004 8676 30060 8732
rect 30060 8676 30064 8732
rect 30000 8672 30064 8676
rect 30080 8732 30144 8736
rect 30080 8676 30084 8732
rect 30084 8676 30140 8732
rect 30140 8676 30144 8732
rect 30080 8672 30144 8676
rect 44284 8732 44348 8736
rect 44284 8676 44288 8732
rect 44288 8676 44344 8732
rect 44344 8676 44348 8732
rect 44284 8672 44348 8676
rect 44364 8732 44428 8736
rect 44364 8676 44368 8732
rect 44368 8676 44424 8732
rect 44424 8676 44428 8732
rect 44364 8672 44428 8676
rect 44444 8732 44508 8736
rect 44444 8676 44448 8732
rect 44448 8676 44504 8732
rect 44504 8676 44508 8732
rect 44444 8672 44508 8676
rect 44524 8732 44588 8736
rect 44524 8676 44528 8732
rect 44528 8676 44584 8732
rect 44584 8676 44588 8732
rect 44524 8672 44588 8676
rect 58728 8732 58792 8736
rect 58728 8676 58732 8732
rect 58732 8676 58788 8732
rect 58788 8676 58792 8732
rect 58728 8672 58792 8676
rect 58808 8732 58872 8736
rect 58808 8676 58812 8732
rect 58812 8676 58868 8732
rect 58868 8676 58872 8732
rect 58808 8672 58872 8676
rect 58888 8732 58952 8736
rect 58888 8676 58892 8732
rect 58892 8676 58948 8732
rect 58948 8676 58952 8732
rect 58888 8672 58952 8676
rect 58968 8732 59032 8736
rect 58968 8676 58972 8732
rect 58972 8676 59028 8732
rect 59028 8676 59032 8732
rect 58968 8672 59032 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 22618 8188 22682 8192
rect 22618 8132 22622 8188
rect 22622 8132 22678 8188
rect 22678 8132 22682 8188
rect 22618 8128 22682 8132
rect 22698 8188 22762 8192
rect 22698 8132 22702 8188
rect 22702 8132 22758 8188
rect 22758 8132 22762 8188
rect 22698 8128 22762 8132
rect 22778 8188 22842 8192
rect 22778 8132 22782 8188
rect 22782 8132 22838 8188
rect 22838 8132 22842 8188
rect 22778 8128 22842 8132
rect 22858 8188 22922 8192
rect 22858 8132 22862 8188
rect 22862 8132 22918 8188
rect 22918 8132 22922 8188
rect 22858 8128 22922 8132
rect 37062 8188 37126 8192
rect 37062 8132 37066 8188
rect 37066 8132 37122 8188
rect 37122 8132 37126 8188
rect 37062 8128 37126 8132
rect 37142 8188 37206 8192
rect 37142 8132 37146 8188
rect 37146 8132 37202 8188
rect 37202 8132 37206 8188
rect 37142 8128 37206 8132
rect 37222 8188 37286 8192
rect 37222 8132 37226 8188
rect 37226 8132 37282 8188
rect 37282 8132 37286 8188
rect 37222 8128 37286 8132
rect 37302 8188 37366 8192
rect 37302 8132 37306 8188
rect 37306 8132 37362 8188
rect 37362 8132 37366 8188
rect 37302 8128 37366 8132
rect 51506 8188 51570 8192
rect 51506 8132 51510 8188
rect 51510 8132 51566 8188
rect 51566 8132 51570 8188
rect 51506 8128 51570 8132
rect 51586 8188 51650 8192
rect 51586 8132 51590 8188
rect 51590 8132 51646 8188
rect 51646 8132 51650 8188
rect 51586 8128 51650 8132
rect 51666 8188 51730 8192
rect 51666 8132 51670 8188
rect 51670 8132 51726 8188
rect 51726 8132 51730 8188
rect 51666 8128 51730 8132
rect 51746 8188 51810 8192
rect 51746 8132 51750 8188
rect 51750 8132 51806 8188
rect 51806 8132 51810 8188
rect 51746 8128 51810 8132
rect 15396 7644 15460 7648
rect 15396 7588 15400 7644
rect 15400 7588 15456 7644
rect 15456 7588 15460 7644
rect 15396 7584 15460 7588
rect 15476 7644 15540 7648
rect 15476 7588 15480 7644
rect 15480 7588 15536 7644
rect 15536 7588 15540 7644
rect 15476 7584 15540 7588
rect 15556 7644 15620 7648
rect 15556 7588 15560 7644
rect 15560 7588 15616 7644
rect 15616 7588 15620 7644
rect 15556 7584 15620 7588
rect 15636 7644 15700 7648
rect 15636 7588 15640 7644
rect 15640 7588 15696 7644
rect 15696 7588 15700 7644
rect 15636 7584 15700 7588
rect 29840 7644 29904 7648
rect 29840 7588 29844 7644
rect 29844 7588 29900 7644
rect 29900 7588 29904 7644
rect 29840 7584 29904 7588
rect 29920 7644 29984 7648
rect 29920 7588 29924 7644
rect 29924 7588 29980 7644
rect 29980 7588 29984 7644
rect 29920 7584 29984 7588
rect 30000 7644 30064 7648
rect 30000 7588 30004 7644
rect 30004 7588 30060 7644
rect 30060 7588 30064 7644
rect 30000 7584 30064 7588
rect 30080 7644 30144 7648
rect 30080 7588 30084 7644
rect 30084 7588 30140 7644
rect 30140 7588 30144 7644
rect 30080 7584 30144 7588
rect 44284 7644 44348 7648
rect 44284 7588 44288 7644
rect 44288 7588 44344 7644
rect 44344 7588 44348 7644
rect 44284 7584 44348 7588
rect 44364 7644 44428 7648
rect 44364 7588 44368 7644
rect 44368 7588 44424 7644
rect 44424 7588 44428 7644
rect 44364 7584 44428 7588
rect 44444 7644 44508 7648
rect 44444 7588 44448 7644
rect 44448 7588 44504 7644
rect 44504 7588 44508 7644
rect 44444 7584 44508 7588
rect 44524 7644 44588 7648
rect 44524 7588 44528 7644
rect 44528 7588 44584 7644
rect 44584 7588 44588 7644
rect 44524 7584 44588 7588
rect 58728 7644 58792 7648
rect 58728 7588 58732 7644
rect 58732 7588 58788 7644
rect 58788 7588 58792 7644
rect 58728 7584 58792 7588
rect 58808 7644 58872 7648
rect 58808 7588 58812 7644
rect 58812 7588 58868 7644
rect 58868 7588 58872 7644
rect 58808 7584 58872 7588
rect 58888 7644 58952 7648
rect 58888 7588 58892 7644
rect 58892 7588 58948 7644
rect 58948 7588 58952 7644
rect 58888 7584 58952 7588
rect 58968 7644 59032 7648
rect 58968 7588 58972 7644
rect 58972 7588 59028 7644
rect 59028 7588 59032 7644
rect 58968 7584 59032 7588
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 22618 7100 22682 7104
rect 22618 7044 22622 7100
rect 22622 7044 22678 7100
rect 22678 7044 22682 7100
rect 22618 7040 22682 7044
rect 22698 7100 22762 7104
rect 22698 7044 22702 7100
rect 22702 7044 22758 7100
rect 22758 7044 22762 7100
rect 22698 7040 22762 7044
rect 22778 7100 22842 7104
rect 22778 7044 22782 7100
rect 22782 7044 22838 7100
rect 22838 7044 22842 7100
rect 22778 7040 22842 7044
rect 22858 7100 22922 7104
rect 22858 7044 22862 7100
rect 22862 7044 22918 7100
rect 22918 7044 22922 7100
rect 22858 7040 22922 7044
rect 37062 7100 37126 7104
rect 37062 7044 37066 7100
rect 37066 7044 37122 7100
rect 37122 7044 37126 7100
rect 37062 7040 37126 7044
rect 37142 7100 37206 7104
rect 37142 7044 37146 7100
rect 37146 7044 37202 7100
rect 37202 7044 37206 7100
rect 37142 7040 37206 7044
rect 37222 7100 37286 7104
rect 37222 7044 37226 7100
rect 37226 7044 37282 7100
rect 37282 7044 37286 7100
rect 37222 7040 37286 7044
rect 37302 7100 37366 7104
rect 37302 7044 37306 7100
rect 37306 7044 37362 7100
rect 37362 7044 37366 7100
rect 37302 7040 37366 7044
rect 51506 7100 51570 7104
rect 51506 7044 51510 7100
rect 51510 7044 51566 7100
rect 51566 7044 51570 7100
rect 51506 7040 51570 7044
rect 51586 7100 51650 7104
rect 51586 7044 51590 7100
rect 51590 7044 51646 7100
rect 51646 7044 51650 7100
rect 51586 7040 51650 7044
rect 51666 7100 51730 7104
rect 51666 7044 51670 7100
rect 51670 7044 51726 7100
rect 51726 7044 51730 7100
rect 51666 7040 51730 7044
rect 51746 7100 51810 7104
rect 51746 7044 51750 7100
rect 51750 7044 51806 7100
rect 51806 7044 51810 7100
rect 51746 7040 51810 7044
rect 15396 6556 15460 6560
rect 15396 6500 15400 6556
rect 15400 6500 15456 6556
rect 15456 6500 15460 6556
rect 15396 6496 15460 6500
rect 15476 6556 15540 6560
rect 15476 6500 15480 6556
rect 15480 6500 15536 6556
rect 15536 6500 15540 6556
rect 15476 6496 15540 6500
rect 15556 6556 15620 6560
rect 15556 6500 15560 6556
rect 15560 6500 15616 6556
rect 15616 6500 15620 6556
rect 15556 6496 15620 6500
rect 15636 6556 15700 6560
rect 15636 6500 15640 6556
rect 15640 6500 15696 6556
rect 15696 6500 15700 6556
rect 15636 6496 15700 6500
rect 29840 6556 29904 6560
rect 29840 6500 29844 6556
rect 29844 6500 29900 6556
rect 29900 6500 29904 6556
rect 29840 6496 29904 6500
rect 29920 6556 29984 6560
rect 29920 6500 29924 6556
rect 29924 6500 29980 6556
rect 29980 6500 29984 6556
rect 29920 6496 29984 6500
rect 30000 6556 30064 6560
rect 30000 6500 30004 6556
rect 30004 6500 30060 6556
rect 30060 6500 30064 6556
rect 30000 6496 30064 6500
rect 30080 6556 30144 6560
rect 30080 6500 30084 6556
rect 30084 6500 30140 6556
rect 30140 6500 30144 6556
rect 30080 6496 30144 6500
rect 44284 6556 44348 6560
rect 44284 6500 44288 6556
rect 44288 6500 44344 6556
rect 44344 6500 44348 6556
rect 44284 6496 44348 6500
rect 44364 6556 44428 6560
rect 44364 6500 44368 6556
rect 44368 6500 44424 6556
rect 44424 6500 44428 6556
rect 44364 6496 44428 6500
rect 44444 6556 44508 6560
rect 44444 6500 44448 6556
rect 44448 6500 44504 6556
rect 44504 6500 44508 6556
rect 44444 6496 44508 6500
rect 44524 6556 44588 6560
rect 44524 6500 44528 6556
rect 44528 6500 44584 6556
rect 44584 6500 44588 6556
rect 44524 6496 44588 6500
rect 58728 6556 58792 6560
rect 58728 6500 58732 6556
rect 58732 6500 58788 6556
rect 58788 6500 58792 6556
rect 58728 6496 58792 6500
rect 58808 6556 58872 6560
rect 58808 6500 58812 6556
rect 58812 6500 58868 6556
rect 58868 6500 58872 6556
rect 58808 6496 58872 6500
rect 58888 6556 58952 6560
rect 58888 6500 58892 6556
rect 58892 6500 58948 6556
rect 58948 6500 58952 6556
rect 58888 6496 58952 6500
rect 58968 6556 59032 6560
rect 58968 6500 58972 6556
rect 58972 6500 59028 6556
rect 59028 6500 59032 6556
rect 58968 6496 59032 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 22618 6012 22682 6016
rect 22618 5956 22622 6012
rect 22622 5956 22678 6012
rect 22678 5956 22682 6012
rect 22618 5952 22682 5956
rect 22698 6012 22762 6016
rect 22698 5956 22702 6012
rect 22702 5956 22758 6012
rect 22758 5956 22762 6012
rect 22698 5952 22762 5956
rect 22778 6012 22842 6016
rect 22778 5956 22782 6012
rect 22782 5956 22838 6012
rect 22838 5956 22842 6012
rect 22778 5952 22842 5956
rect 22858 6012 22922 6016
rect 22858 5956 22862 6012
rect 22862 5956 22918 6012
rect 22918 5956 22922 6012
rect 22858 5952 22922 5956
rect 37062 6012 37126 6016
rect 37062 5956 37066 6012
rect 37066 5956 37122 6012
rect 37122 5956 37126 6012
rect 37062 5952 37126 5956
rect 37142 6012 37206 6016
rect 37142 5956 37146 6012
rect 37146 5956 37202 6012
rect 37202 5956 37206 6012
rect 37142 5952 37206 5956
rect 37222 6012 37286 6016
rect 37222 5956 37226 6012
rect 37226 5956 37282 6012
rect 37282 5956 37286 6012
rect 37222 5952 37286 5956
rect 37302 6012 37366 6016
rect 37302 5956 37306 6012
rect 37306 5956 37362 6012
rect 37362 5956 37366 6012
rect 37302 5952 37366 5956
rect 51506 6012 51570 6016
rect 51506 5956 51510 6012
rect 51510 5956 51566 6012
rect 51566 5956 51570 6012
rect 51506 5952 51570 5956
rect 51586 6012 51650 6016
rect 51586 5956 51590 6012
rect 51590 5956 51646 6012
rect 51646 5956 51650 6012
rect 51586 5952 51650 5956
rect 51666 6012 51730 6016
rect 51666 5956 51670 6012
rect 51670 5956 51726 6012
rect 51726 5956 51730 6012
rect 51666 5952 51730 5956
rect 51746 6012 51810 6016
rect 51746 5956 51750 6012
rect 51750 5956 51806 6012
rect 51806 5956 51810 6012
rect 51746 5952 51810 5956
rect 15396 5468 15460 5472
rect 15396 5412 15400 5468
rect 15400 5412 15456 5468
rect 15456 5412 15460 5468
rect 15396 5408 15460 5412
rect 15476 5468 15540 5472
rect 15476 5412 15480 5468
rect 15480 5412 15536 5468
rect 15536 5412 15540 5468
rect 15476 5408 15540 5412
rect 15556 5468 15620 5472
rect 15556 5412 15560 5468
rect 15560 5412 15616 5468
rect 15616 5412 15620 5468
rect 15556 5408 15620 5412
rect 15636 5468 15700 5472
rect 15636 5412 15640 5468
rect 15640 5412 15696 5468
rect 15696 5412 15700 5468
rect 15636 5408 15700 5412
rect 29840 5468 29904 5472
rect 29840 5412 29844 5468
rect 29844 5412 29900 5468
rect 29900 5412 29904 5468
rect 29840 5408 29904 5412
rect 29920 5468 29984 5472
rect 29920 5412 29924 5468
rect 29924 5412 29980 5468
rect 29980 5412 29984 5468
rect 29920 5408 29984 5412
rect 30000 5468 30064 5472
rect 30000 5412 30004 5468
rect 30004 5412 30060 5468
rect 30060 5412 30064 5468
rect 30000 5408 30064 5412
rect 30080 5468 30144 5472
rect 30080 5412 30084 5468
rect 30084 5412 30140 5468
rect 30140 5412 30144 5468
rect 30080 5408 30144 5412
rect 44284 5468 44348 5472
rect 44284 5412 44288 5468
rect 44288 5412 44344 5468
rect 44344 5412 44348 5468
rect 44284 5408 44348 5412
rect 44364 5468 44428 5472
rect 44364 5412 44368 5468
rect 44368 5412 44424 5468
rect 44424 5412 44428 5468
rect 44364 5408 44428 5412
rect 44444 5468 44508 5472
rect 44444 5412 44448 5468
rect 44448 5412 44504 5468
rect 44504 5412 44508 5468
rect 44444 5408 44508 5412
rect 44524 5468 44588 5472
rect 44524 5412 44528 5468
rect 44528 5412 44584 5468
rect 44584 5412 44588 5468
rect 44524 5408 44588 5412
rect 58728 5468 58792 5472
rect 58728 5412 58732 5468
rect 58732 5412 58788 5468
rect 58788 5412 58792 5468
rect 58728 5408 58792 5412
rect 58808 5468 58872 5472
rect 58808 5412 58812 5468
rect 58812 5412 58868 5468
rect 58868 5412 58872 5468
rect 58808 5408 58872 5412
rect 58888 5468 58952 5472
rect 58888 5412 58892 5468
rect 58892 5412 58948 5468
rect 58948 5412 58952 5468
rect 58888 5408 58952 5412
rect 58968 5468 59032 5472
rect 58968 5412 58972 5468
rect 58972 5412 59028 5468
rect 59028 5412 59032 5468
rect 58968 5408 59032 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 22618 4924 22682 4928
rect 22618 4868 22622 4924
rect 22622 4868 22678 4924
rect 22678 4868 22682 4924
rect 22618 4864 22682 4868
rect 22698 4924 22762 4928
rect 22698 4868 22702 4924
rect 22702 4868 22758 4924
rect 22758 4868 22762 4924
rect 22698 4864 22762 4868
rect 22778 4924 22842 4928
rect 22778 4868 22782 4924
rect 22782 4868 22838 4924
rect 22838 4868 22842 4924
rect 22778 4864 22842 4868
rect 22858 4924 22922 4928
rect 22858 4868 22862 4924
rect 22862 4868 22918 4924
rect 22918 4868 22922 4924
rect 22858 4864 22922 4868
rect 37062 4924 37126 4928
rect 37062 4868 37066 4924
rect 37066 4868 37122 4924
rect 37122 4868 37126 4924
rect 37062 4864 37126 4868
rect 37142 4924 37206 4928
rect 37142 4868 37146 4924
rect 37146 4868 37202 4924
rect 37202 4868 37206 4924
rect 37142 4864 37206 4868
rect 37222 4924 37286 4928
rect 37222 4868 37226 4924
rect 37226 4868 37282 4924
rect 37282 4868 37286 4924
rect 37222 4864 37286 4868
rect 37302 4924 37366 4928
rect 37302 4868 37306 4924
rect 37306 4868 37362 4924
rect 37362 4868 37366 4924
rect 37302 4864 37366 4868
rect 51506 4924 51570 4928
rect 51506 4868 51510 4924
rect 51510 4868 51566 4924
rect 51566 4868 51570 4924
rect 51506 4864 51570 4868
rect 51586 4924 51650 4928
rect 51586 4868 51590 4924
rect 51590 4868 51646 4924
rect 51646 4868 51650 4924
rect 51586 4864 51650 4868
rect 51666 4924 51730 4928
rect 51666 4868 51670 4924
rect 51670 4868 51726 4924
rect 51726 4868 51730 4924
rect 51666 4864 51730 4868
rect 51746 4924 51810 4928
rect 51746 4868 51750 4924
rect 51750 4868 51806 4924
rect 51806 4868 51810 4924
rect 51746 4864 51810 4868
rect 15396 4380 15460 4384
rect 15396 4324 15400 4380
rect 15400 4324 15456 4380
rect 15456 4324 15460 4380
rect 15396 4320 15460 4324
rect 15476 4380 15540 4384
rect 15476 4324 15480 4380
rect 15480 4324 15536 4380
rect 15536 4324 15540 4380
rect 15476 4320 15540 4324
rect 15556 4380 15620 4384
rect 15556 4324 15560 4380
rect 15560 4324 15616 4380
rect 15616 4324 15620 4380
rect 15556 4320 15620 4324
rect 15636 4380 15700 4384
rect 15636 4324 15640 4380
rect 15640 4324 15696 4380
rect 15696 4324 15700 4380
rect 15636 4320 15700 4324
rect 29840 4380 29904 4384
rect 29840 4324 29844 4380
rect 29844 4324 29900 4380
rect 29900 4324 29904 4380
rect 29840 4320 29904 4324
rect 29920 4380 29984 4384
rect 29920 4324 29924 4380
rect 29924 4324 29980 4380
rect 29980 4324 29984 4380
rect 29920 4320 29984 4324
rect 30000 4380 30064 4384
rect 30000 4324 30004 4380
rect 30004 4324 30060 4380
rect 30060 4324 30064 4380
rect 30000 4320 30064 4324
rect 30080 4380 30144 4384
rect 30080 4324 30084 4380
rect 30084 4324 30140 4380
rect 30140 4324 30144 4380
rect 30080 4320 30144 4324
rect 44284 4380 44348 4384
rect 44284 4324 44288 4380
rect 44288 4324 44344 4380
rect 44344 4324 44348 4380
rect 44284 4320 44348 4324
rect 44364 4380 44428 4384
rect 44364 4324 44368 4380
rect 44368 4324 44424 4380
rect 44424 4324 44428 4380
rect 44364 4320 44428 4324
rect 44444 4380 44508 4384
rect 44444 4324 44448 4380
rect 44448 4324 44504 4380
rect 44504 4324 44508 4380
rect 44444 4320 44508 4324
rect 44524 4380 44588 4384
rect 44524 4324 44528 4380
rect 44528 4324 44584 4380
rect 44584 4324 44588 4380
rect 44524 4320 44588 4324
rect 58728 4380 58792 4384
rect 58728 4324 58732 4380
rect 58732 4324 58788 4380
rect 58788 4324 58792 4380
rect 58728 4320 58792 4324
rect 58808 4380 58872 4384
rect 58808 4324 58812 4380
rect 58812 4324 58868 4380
rect 58868 4324 58872 4380
rect 58808 4320 58872 4324
rect 58888 4380 58952 4384
rect 58888 4324 58892 4380
rect 58892 4324 58948 4380
rect 58948 4324 58952 4380
rect 58888 4320 58952 4324
rect 58968 4380 59032 4384
rect 58968 4324 58972 4380
rect 58972 4324 59028 4380
rect 59028 4324 59032 4380
rect 58968 4320 59032 4324
rect 10548 4040 10612 4044
rect 10548 3984 10562 4040
rect 10562 3984 10612 4040
rect 10548 3980 10612 3984
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 22618 3836 22682 3840
rect 22618 3780 22622 3836
rect 22622 3780 22678 3836
rect 22678 3780 22682 3836
rect 22618 3776 22682 3780
rect 22698 3836 22762 3840
rect 22698 3780 22702 3836
rect 22702 3780 22758 3836
rect 22758 3780 22762 3836
rect 22698 3776 22762 3780
rect 22778 3836 22842 3840
rect 22778 3780 22782 3836
rect 22782 3780 22838 3836
rect 22838 3780 22842 3836
rect 22778 3776 22842 3780
rect 22858 3836 22922 3840
rect 22858 3780 22862 3836
rect 22862 3780 22918 3836
rect 22918 3780 22922 3836
rect 22858 3776 22922 3780
rect 37062 3836 37126 3840
rect 37062 3780 37066 3836
rect 37066 3780 37122 3836
rect 37122 3780 37126 3836
rect 37062 3776 37126 3780
rect 37142 3836 37206 3840
rect 37142 3780 37146 3836
rect 37146 3780 37202 3836
rect 37202 3780 37206 3836
rect 37142 3776 37206 3780
rect 37222 3836 37286 3840
rect 37222 3780 37226 3836
rect 37226 3780 37282 3836
rect 37282 3780 37286 3836
rect 37222 3776 37286 3780
rect 37302 3836 37366 3840
rect 37302 3780 37306 3836
rect 37306 3780 37362 3836
rect 37362 3780 37366 3836
rect 37302 3776 37366 3780
rect 51506 3836 51570 3840
rect 51506 3780 51510 3836
rect 51510 3780 51566 3836
rect 51566 3780 51570 3836
rect 51506 3776 51570 3780
rect 51586 3836 51650 3840
rect 51586 3780 51590 3836
rect 51590 3780 51646 3836
rect 51646 3780 51650 3836
rect 51586 3776 51650 3780
rect 51666 3836 51730 3840
rect 51666 3780 51670 3836
rect 51670 3780 51726 3836
rect 51726 3780 51730 3836
rect 51666 3776 51730 3780
rect 51746 3836 51810 3840
rect 51746 3780 51750 3836
rect 51750 3780 51806 3836
rect 51806 3780 51810 3836
rect 51746 3776 51810 3780
rect 37596 3436 37660 3500
rect 15396 3292 15460 3296
rect 15396 3236 15400 3292
rect 15400 3236 15456 3292
rect 15456 3236 15460 3292
rect 15396 3232 15460 3236
rect 15476 3292 15540 3296
rect 15476 3236 15480 3292
rect 15480 3236 15536 3292
rect 15536 3236 15540 3292
rect 15476 3232 15540 3236
rect 15556 3292 15620 3296
rect 15556 3236 15560 3292
rect 15560 3236 15616 3292
rect 15616 3236 15620 3292
rect 15556 3232 15620 3236
rect 15636 3292 15700 3296
rect 15636 3236 15640 3292
rect 15640 3236 15696 3292
rect 15696 3236 15700 3292
rect 15636 3232 15700 3236
rect 29840 3292 29904 3296
rect 29840 3236 29844 3292
rect 29844 3236 29900 3292
rect 29900 3236 29904 3292
rect 29840 3232 29904 3236
rect 29920 3292 29984 3296
rect 29920 3236 29924 3292
rect 29924 3236 29980 3292
rect 29980 3236 29984 3292
rect 29920 3232 29984 3236
rect 30000 3292 30064 3296
rect 30000 3236 30004 3292
rect 30004 3236 30060 3292
rect 30060 3236 30064 3292
rect 30000 3232 30064 3236
rect 30080 3292 30144 3296
rect 30080 3236 30084 3292
rect 30084 3236 30140 3292
rect 30140 3236 30144 3292
rect 30080 3232 30144 3236
rect 44284 3292 44348 3296
rect 44284 3236 44288 3292
rect 44288 3236 44344 3292
rect 44344 3236 44348 3292
rect 44284 3232 44348 3236
rect 44364 3292 44428 3296
rect 44364 3236 44368 3292
rect 44368 3236 44424 3292
rect 44424 3236 44428 3292
rect 44364 3232 44428 3236
rect 44444 3292 44508 3296
rect 44444 3236 44448 3292
rect 44448 3236 44504 3292
rect 44504 3236 44508 3292
rect 44444 3232 44508 3236
rect 44524 3292 44588 3296
rect 44524 3236 44528 3292
rect 44528 3236 44584 3292
rect 44584 3236 44588 3292
rect 44524 3232 44588 3236
rect 58728 3292 58792 3296
rect 58728 3236 58732 3292
rect 58732 3236 58788 3292
rect 58788 3236 58792 3292
rect 58728 3232 58792 3236
rect 58808 3292 58872 3296
rect 58808 3236 58812 3292
rect 58812 3236 58868 3292
rect 58868 3236 58872 3292
rect 58808 3232 58872 3236
rect 58888 3292 58952 3296
rect 58888 3236 58892 3292
rect 58892 3236 58948 3292
rect 58948 3236 58952 3292
rect 58888 3232 58952 3236
rect 58968 3292 59032 3296
rect 58968 3236 58972 3292
rect 58972 3236 59028 3292
rect 59028 3236 59032 3292
rect 58968 3232 59032 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 22618 2748 22682 2752
rect 22618 2692 22622 2748
rect 22622 2692 22678 2748
rect 22678 2692 22682 2748
rect 22618 2688 22682 2692
rect 22698 2748 22762 2752
rect 22698 2692 22702 2748
rect 22702 2692 22758 2748
rect 22758 2692 22762 2748
rect 22698 2688 22762 2692
rect 22778 2748 22842 2752
rect 22778 2692 22782 2748
rect 22782 2692 22838 2748
rect 22838 2692 22842 2748
rect 22778 2688 22842 2692
rect 22858 2748 22922 2752
rect 22858 2692 22862 2748
rect 22862 2692 22918 2748
rect 22918 2692 22922 2748
rect 22858 2688 22922 2692
rect 37062 2748 37126 2752
rect 37062 2692 37066 2748
rect 37066 2692 37122 2748
rect 37122 2692 37126 2748
rect 37062 2688 37126 2692
rect 37142 2748 37206 2752
rect 37142 2692 37146 2748
rect 37146 2692 37202 2748
rect 37202 2692 37206 2748
rect 37142 2688 37206 2692
rect 37222 2748 37286 2752
rect 37222 2692 37226 2748
rect 37226 2692 37282 2748
rect 37282 2692 37286 2748
rect 37222 2688 37286 2692
rect 37302 2748 37366 2752
rect 37302 2692 37306 2748
rect 37306 2692 37362 2748
rect 37362 2692 37366 2748
rect 37302 2688 37366 2692
rect 51506 2748 51570 2752
rect 51506 2692 51510 2748
rect 51510 2692 51566 2748
rect 51566 2692 51570 2748
rect 51506 2688 51570 2692
rect 51586 2748 51650 2752
rect 51586 2692 51590 2748
rect 51590 2692 51646 2748
rect 51646 2692 51650 2748
rect 51586 2688 51650 2692
rect 51666 2748 51730 2752
rect 51666 2692 51670 2748
rect 51670 2692 51726 2748
rect 51726 2692 51730 2748
rect 51666 2688 51730 2692
rect 51746 2748 51810 2752
rect 51746 2692 51750 2748
rect 51750 2692 51806 2748
rect 51806 2692 51810 2748
rect 51746 2688 51810 2692
rect 15396 2204 15460 2208
rect 15396 2148 15400 2204
rect 15400 2148 15456 2204
rect 15456 2148 15460 2204
rect 15396 2144 15460 2148
rect 15476 2204 15540 2208
rect 15476 2148 15480 2204
rect 15480 2148 15536 2204
rect 15536 2148 15540 2204
rect 15476 2144 15540 2148
rect 15556 2204 15620 2208
rect 15556 2148 15560 2204
rect 15560 2148 15616 2204
rect 15616 2148 15620 2204
rect 15556 2144 15620 2148
rect 15636 2204 15700 2208
rect 15636 2148 15640 2204
rect 15640 2148 15696 2204
rect 15696 2148 15700 2204
rect 15636 2144 15700 2148
rect 29840 2204 29904 2208
rect 29840 2148 29844 2204
rect 29844 2148 29900 2204
rect 29900 2148 29904 2204
rect 29840 2144 29904 2148
rect 29920 2204 29984 2208
rect 29920 2148 29924 2204
rect 29924 2148 29980 2204
rect 29980 2148 29984 2204
rect 29920 2144 29984 2148
rect 30000 2204 30064 2208
rect 30000 2148 30004 2204
rect 30004 2148 30060 2204
rect 30060 2148 30064 2204
rect 30000 2144 30064 2148
rect 30080 2204 30144 2208
rect 30080 2148 30084 2204
rect 30084 2148 30140 2204
rect 30140 2148 30144 2204
rect 30080 2144 30144 2148
rect 44284 2204 44348 2208
rect 44284 2148 44288 2204
rect 44288 2148 44344 2204
rect 44344 2148 44348 2204
rect 44284 2144 44348 2148
rect 44364 2204 44428 2208
rect 44364 2148 44368 2204
rect 44368 2148 44424 2204
rect 44424 2148 44428 2204
rect 44364 2144 44428 2148
rect 44444 2204 44508 2208
rect 44444 2148 44448 2204
rect 44448 2148 44504 2204
rect 44504 2148 44508 2204
rect 44444 2144 44508 2148
rect 44524 2204 44588 2208
rect 44524 2148 44528 2204
rect 44528 2148 44584 2204
rect 44584 2148 44588 2204
rect 44524 2144 44588 2148
rect 58728 2204 58792 2208
rect 58728 2148 58732 2204
rect 58732 2148 58788 2204
rect 58788 2148 58792 2204
rect 58728 2144 58792 2148
rect 58808 2204 58872 2208
rect 58808 2148 58812 2204
rect 58812 2148 58868 2204
rect 58868 2148 58872 2204
rect 58808 2144 58872 2148
rect 58888 2204 58952 2208
rect 58888 2148 58892 2204
rect 58892 2148 58948 2204
rect 58948 2148 58952 2204
rect 58888 2144 58952 2148
rect 58968 2204 59032 2208
rect 58968 2148 58972 2204
rect 58972 2148 59028 2204
rect 59028 2148 59032 2204
rect 58968 2144 59032 2148
<< metal4 >>
rect 8166 27776 8486 27792
rect 8166 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8486 27776
rect 8166 26688 8486 27712
rect 8166 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8486 26688
rect 8166 25600 8486 26624
rect 8166 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8486 25600
rect 8166 24512 8486 25536
rect 8166 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8486 24512
rect 8166 23424 8486 24448
rect 8166 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8486 23424
rect 8166 22336 8486 23360
rect 8166 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8486 22336
rect 8166 21248 8486 22272
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 15388 27232 15708 27792
rect 15388 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15708 27232
rect 15388 26144 15708 27168
rect 15388 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15708 26144
rect 15388 25056 15708 26080
rect 15388 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15708 25056
rect 15388 23968 15708 24992
rect 15388 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15708 23968
rect 15388 22880 15708 23904
rect 15388 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15708 22880
rect 15388 21792 15708 22816
rect 15388 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15708 21792
rect 15388 20704 15708 21728
rect 15388 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15708 20704
rect 15388 19616 15708 20640
rect 15388 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15708 19616
rect 10179 19412 10245 19413
rect 10179 19348 10180 19412
rect 10244 19348 10245 19412
rect 10179 19347 10245 19348
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 9811 16692 9877 16693
rect 9811 16628 9812 16692
rect 9876 16628 9877 16692
rect 9811 16627 9877 16628
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 9814 9485 9874 16627
rect 10182 12450 10242 19347
rect 15388 18528 15708 19552
rect 15388 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15708 18528
rect 15388 17440 15708 18464
rect 15388 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15708 17440
rect 15388 16352 15708 17376
rect 15388 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15708 16352
rect 15388 15264 15708 16288
rect 15388 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15708 15264
rect 15388 14176 15708 15200
rect 15388 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15708 14176
rect 15388 13088 15708 14112
rect 15388 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15708 13088
rect 10182 12390 10610 12450
rect 10550 11117 10610 12390
rect 15388 12000 15708 13024
rect 15388 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15708 12000
rect 10547 11116 10613 11117
rect 10547 11052 10548 11116
rect 10612 11052 10613 11116
rect 10547 11051 10613 11052
rect 9811 9484 9877 9485
rect 9811 9420 9812 9484
rect 9876 9420 9877 9484
rect 9811 9419 9877 9420
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 10550 4045 10610 11051
rect 15388 10912 15708 11936
rect 15388 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15708 10912
rect 15388 9824 15708 10848
rect 15388 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15708 9824
rect 15388 8736 15708 9760
rect 15388 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15708 8736
rect 15388 7648 15708 8672
rect 15388 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15708 7648
rect 15388 6560 15708 7584
rect 15388 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15708 6560
rect 15388 5472 15708 6496
rect 15388 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15708 5472
rect 15388 4384 15708 5408
rect 15388 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15708 4384
rect 10547 4044 10613 4045
rect 10547 3980 10548 4044
rect 10612 3980 10613 4044
rect 10547 3979 10613 3980
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 2128 8486 2688
rect 15388 3296 15708 4320
rect 15388 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15708 3296
rect 15388 2208 15708 3232
rect 15388 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15708 2208
rect 15388 2128 15708 2144
rect 22610 27776 22930 27792
rect 22610 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22930 27776
rect 22610 26688 22930 27712
rect 22610 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22930 26688
rect 22610 25600 22930 26624
rect 22610 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22930 25600
rect 22610 24512 22930 25536
rect 22610 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22930 24512
rect 22610 23424 22930 24448
rect 22610 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22930 23424
rect 22610 22336 22930 23360
rect 22610 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22930 22336
rect 22610 21248 22930 22272
rect 22610 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22930 21248
rect 22610 20160 22930 21184
rect 22610 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22930 20160
rect 22610 19072 22930 20096
rect 22610 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22930 19072
rect 22610 17984 22930 19008
rect 22610 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22930 17984
rect 22610 16896 22930 17920
rect 22610 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22930 16896
rect 22610 15808 22930 16832
rect 22610 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22930 15808
rect 22610 14720 22930 15744
rect 22610 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22930 14720
rect 22610 13632 22930 14656
rect 22610 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22930 13632
rect 22610 12544 22930 13568
rect 22610 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22930 12544
rect 22610 11456 22930 12480
rect 22610 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22930 11456
rect 22610 10368 22930 11392
rect 22610 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22930 10368
rect 22610 9280 22930 10304
rect 22610 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22930 9280
rect 22610 8192 22930 9216
rect 22610 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22930 8192
rect 22610 7104 22930 8128
rect 22610 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22930 7104
rect 22610 6016 22930 7040
rect 22610 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22930 6016
rect 22610 4928 22930 5952
rect 22610 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22930 4928
rect 22610 3840 22930 4864
rect 22610 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22930 3840
rect 22610 2752 22930 3776
rect 22610 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22930 2752
rect 22610 2128 22930 2688
rect 29832 27232 30152 27792
rect 29832 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30152 27232
rect 29832 26144 30152 27168
rect 29832 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30152 26144
rect 29832 25056 30152 26080
rect 29832 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30152 25056
rect 29832 23968 30152 24992
rect 29832 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30152 23968
rect 29832 22880 30152 23904
rect 29832 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30152 22880
rect 29832 21792 30152 22816
rect 29832 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30152 21792
rect 29832 20704 30152 21728
rect 29832 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30152 20704
rect 29832 19616 30152 20640
rect 29832 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30152 19616
rect 29832 18528 30152 19552
rect 29832 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30152 18528
rect 29832 17440 30152 18464
rect 29832 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30152 17440
rect 29832 16352 30152 17376
rect 37054 27776 37374 27792
rect 37054 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37374 27776
rect 37054 26688 37374 27712
rect 37054 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37374 26688
rect 37054 25600 37374 26624
rect 37054 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37374 25600
rect 37054 24512 37374 25536
rect 37054 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37374 24512
rect 37054 23424 37374 24448
rect 37054 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37374 23424
rect 37054 22336 37374 23360
rect 37054 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37374 22336
rect 37054 21248 37374 22272
rect 37054 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37374 21248
rect 37054 20160 37374 21184
rect 37054 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37374 20160
rect 37054 19072 37374 20096
rect 37054 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37374 19072
rect 37054 17984 37374 19008
rect 37054 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37374 17984
rect 37054 16896 37374 17920
rect 37054 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37374 16896
rect 34283 16692 34349 16693
rect 34283 16628 34284 16692
rect 34348 16628 34349 16692
rect 34283 16627 34349 16628
rect 29832 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30152 16352
rect 29832 15264 30152 16288
rect 29832 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30152 15264
rect 29832 14176 30152 15200
rect 29832 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30152 14176
rect 29832 13088 30152 14112
rect 29832 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30152 13088
rect 29832 12000 30152 13024
rect 29832 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30152 12000
rect 29832 10912 30152 11936
rect 29832 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30152 10912
rect 29832 9824 30152 10848
rect 29832 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30152 9824
rect 29832 8736 30152 9760
rect 34286 9621 34346 16627
rect 37054 15808 37374 16832
rect 37054 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37374 15808
rect 37054 14720 37374 15744
rect 37054 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37374 14720
rect 37054 13632 37374 14656
rect 37054 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37374 13632
rect 37054 12544 37374 13568
rect 37054 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37374 12544
rect 37054 11456 37374 12480
rect 37054 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37374 11456
rect 37054 10368 37374 11392
rect 44276 27232 44596 27792
rect 44276 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44596 27232
rect 44276 26144 44596 27168
rect 44276 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44596 26144
rect 44276 25056 44596 26080
rect 44276 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44596 25056
rect 44276 23968 44596 24992
rect 44276 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44596 23968
rect 44276 22880 44596 23904
rect 44276 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44596 22880
rect 44276 21792 44596 22816
rect 44276 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44596 21792
rect 44276 20704 44596 21728
rect 44276 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44596 20704
rect 44276 19616 44596 20640
rect 44276 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44596 19616
rect 44276 18528 44596 19552
rect 44276 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44596 18528
rect 44276 17440 44596 18464
rect 44276 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44596 17440
rect 44276 16352 44596 17376
rect 44276 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44596 16352
rect 44276 15264 44596 16288
rect 44276 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44596 15264
rect 44276 14176 44596 15200
rect 44276 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44596 14176
rect 44276 13088 44596 14112
rect 44276 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44596 13088
rect 44276 12000 44596 13024
rect 44276 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44596 12000
rect 37595 11116 37661 11117
rect 37595 11052 37596 11116
rect 37660 11052 37661 11116
rect 37595 11051 37661 11052
rect 37054 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37374 10368
rect 34283 9620 34349 9621
rect 34283 9556 34284 9620
rect 34348 9556 34349 9620
rect 34283 9555 34349 9556
rect 29832 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30152 8736
rect 29832 7648 30152 8672
rect 29832 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30152 7648
rect 29832 6560 30152 7584
rect 29832 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30152 6560
rect 29832 5472 30152 6496
rect 29832 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30152 5472
rect 29832 4384 30152 5408
rect 29832 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30152 4384
rect 29832 3296 30152 4320
rect 29832 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30152 3296
rect 29832 2208 30152 3232
rect 29832 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30152 2208
rect 29832 2128 30152 2144
rect 37054 9280 37374 10304
rect 37054 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37374 9280
rect 37054 8192 37374 9216
rect 37054 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37374 8192
rect 37054 7104 37374 8128
rect 37054 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37374 7104
rect 37054 6016 37374 7040
rect 37054 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37374 6016
rect 37054 4928 37374 5952
rect 37054 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37374 4928
rect 37054 3840 37374 4864
rect 37054 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37374 3840
rect 37054 2752 37374 3776
rect 37598 3501 37658 11051
rect 44276 10912 44596 11936
rect 44276 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44596 10912
rect 44276 9824 44596 10848
rect 44276 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44596 9824
rect 44276 8736 44596 9760
rect 44276 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44596 8736
rect 44276 7648 44596 8672
rect 44276 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44596 7648
rect 44276 6560 44596 7584
rect 44276 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44596 6560
rect 44276 5472 44596 6496
rect 44276 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44596 5472
rect 44276 4384 44596 5408
rect 44276 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44596 4384
rect 37595 3500 37661 3501
rect 37595 3436 37596 3500
rect 37660 3436 37661 3500
rect 37595 3435 37661 3436
rect 37054 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37374 2752
rect 37054 2128 37374 2688
rect 44276 3296 44596 4320
rect 44276 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44596 3296
rect 44276 2208 44596 3232
rect 44276 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44596 2208
rect 44276 2128 44596 2144
rect 51498 27776 51818 27792
rect 51498 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51818 27776
rect 51498 26688 51818 27712
rect 51498 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51818 26688
rect 51498 25600 51818 26624
rect 51498 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51818 25600
rect 51498 24512 51818 25536
rect 51498 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51818 24512
rect 51498 23424 51818 24448
rect 51498 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51818 23424
rect 51498 22336 51818 23360
rect 51498 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51818 22336
rect 51498 21248 51818 22272
rect 51498 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51818 21248
rect 51498 20160 51818 21184
rect 51498 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51818 20160
rect 51498 19072 51818 20096
rect 51498 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51818 19072
rect 51498 17984 51818 19008
rect 51498 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51818 17984
rect 51498 16896 51818 17920
rect 51498 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51818 16896
rect 51498 15808 51818 16832
rect 51498 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51818 15808
rect 51498 14720 51818 15744
rect 51498 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51818 14720
rect 51498 13632 51818 14656
rect 51498 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51818 13632
rect 51498 12544 51818 13568
rect 51498 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51818 12544
rect 51498 11456 51818 12480
rect 51498 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51818 11456
rect 51498 10368 51818 11392
rect 51498 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51818 10368
rect 51498 9280 51818 10304
rect 51498 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51818 9280
rect 51498 8192 51818 9216
rect 51498 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51818 8192
rect 51498 7104 51818 8128
rect 51498 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51818 7104
rect 51498 6016 51818 7040
rect 51498 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51818 6016
rect 51498 4928 51818 5952
rect 51498 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51818 4928
rect 51498 3840 51818 4864
rect 51498 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51818 3840
rect 51498 2752 51818 3776
rect 51498 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51818 2752
rect 51498 2128 51818 2688
rect 58720 27232 59040 27792
rect 58720 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59040 27232
rect 58720 26144 59040 27168
rect 58720 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59040 26144
rect 58720 25056 59040 26080
rect 58720 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59040 25056
rect 58720 23968 59040 24992
rect 58720 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59040 23968
rect 58720 22880 59040 23904
rect 58720 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59040 22880
rect 58720 21792 59040 22816
rect 58720 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59040 21792
rect 58720 20704 59040 21728
rect 58720 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59040 20704
rect 58720 19616 59040 20640
rect 58720 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59040 19616
rect 58720 18528 59040 19552
rect 58720 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59040 18528
rect 58720 17440 59040 18464
rect 58720 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59040 17440
rect 58720 16352 59040 17376
rect 58720 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59040 16352
rect 58720 15264 59040 16288
rect 58720 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59040 15264
rect 58720 14176 59040 15200
rect 58720 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59040 14176
rect 58720 13088 59040 14112
rect 58720 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59040 13088
rect 58720 12000 59040 13024
rect 58720 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59040 12000
rect 58720 10912 59040 11936
rect 58720 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59040 10912
rect 58720 9824 59040 10848
rect 58720 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59040 9824
rect 58720 8736 59040 9760
rect 58720 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59040 8736
rect 58720 7648 59040 8672
rect 58720 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59040 7648
rect 58720 6560 59040 7584
rect 58720 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59040 6560
rect 58720 5472 59040 6496
rect 58720 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59040 5472
rect 58720 4384 59040 5408
rect 58720 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59040 4384
rect 58720 3296 59040 4320
rect 58720 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59040 3296
rect 58720 2208 59040 3232
rect 58720 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59040 2208
rect 58720 2128 59040 2144
use sky130_fd_sc_hd__inv_2  _0517_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1688980957
transform -1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0519_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_4  _0520_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0521_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 45816 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0522_
timestamp 1688980957
transform 1 0 48668 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1688980957
transform -1 0 52440 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0524_
timestamp 1688980957
transform -1 0 52440 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0526_
timestamp 1688980957
transform -1 0 57408 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1688980957
transform 1 0 56212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1688980957
transform 1 0 57132 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0529_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3864 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0530_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0531_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0532_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0533_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0534_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0535_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0536_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0537_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0538_
timestamp 1688980957
transform -1 0 5612 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0539_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0540_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0541_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0542_
timestamp 1688980957
transform -1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0543_
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0545_
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0546_
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0547_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0548_
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0549_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0550_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1688980957
transform 1 0 3404 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0553_
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1688980957
transform 1 0 10580 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0555_
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0557_
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1688980957
transform 1 0 20240 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1688980957
transform 1 0 23552 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1688980957
transform 1 0 27784 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1688980957
transform 1 0 28980 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1688980957
transform 1 0 32384 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1688980957
transform 1 0 35328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1688980957
transform 1 0 35880 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1688980957
transform 1 0 40020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 1688980957
transform -1 0 46460 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1688980957
transform 1 0 50324 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0577_
timestamp 1688980957
transform 1 0 47840 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1688980957
transform -1 0 54740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1688980957
transform 1 0 53636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 1688980957
transform 1 0 53820 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _0582_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1688980957
transform 1 0 3680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1688980957
transform 1 0 6716 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1688980957
transform 1 0 13800 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1688980957
transform 1 0 19412 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1688980957
transform -1 0 21712 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1688980957
transform -1 0 26588 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1688980957
transform -1 0 26496 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform 1 0 30176 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1688980957
transform -1 0 26864 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1688980957
transform 1 0 33304 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1688980957
transform 1 0 30176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform -1 0 35512 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform -1 0 36892 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1688980957
transform -1 0 40204 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1688980957
transform -1 0 43240 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1688980957
transform 1 0 44344 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform -1 0 43332 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1688980957
transform 1 0 46460 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform -1 0 54096 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1688980957
transform 1 0 51612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1688980957
transform 1 0 50968 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1688980957
transform 1 0 56488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1688980957
transform -1 0 57224 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1688980957
transform 1 0 57224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_4  _0615_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1688980957
transform -1 0 6992 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1688980957
transform -1 0 12788 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1688980957
transform -1 0 7176 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 7912 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1688980957
transform -1 0 14168 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform -1 0 18308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1688980957
transform -1 0 22632 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform -1 0 22816 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1688980957
transform -1 0 26680 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform 1 0 27048 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1688980957
transform -1 0 32016 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform -1 0 28888 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1688980957
transform -1 0 33304 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform -1 0 32568 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1688980957
transform 1 0 35328 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform -1 0 40756 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform -1 0 38548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform -1 0 41032 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1688980957
transform -1 0 43240 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform -1 0 49128 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1688980957
transform -1 0 46000 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform -1 0 45080 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1688980957
transform -1 0 48760 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 54188 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform -1 0 52256 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform -1 0 53268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1688980957
transform 1 0 57776 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1688980957
transform 1 0 56580 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1688980957
transform 1 0 56580 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0648_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__mux4_1  _0649_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0650_
timestamp 1688980957
transform -1 0 8832 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0651_
timestamp 1688980957
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0653_
timestamp 1688980957
transform -1 0 13248 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0654_
timestamp 1688980957
transform -1 0 12328 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0656_
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0657_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0658_
timestamp 1688980957
transform -1 0 10212 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1688980957
transform 1 0 10212 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0660_
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0661_
timestamp 1688980957
transform -1 0 8188 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0662_
timestamp 1688980957
transform -1 0 8280 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 1688980957
transform -1 0 8832 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0664_
timestamp 1688980957
transform 1 0 9568 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0665_
timestamp 1688980957
transform -1 0 13800 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0666_
timestamp 1688980957
transform -1 0 13984 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0668_
timestamp 1688980957
transform -1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0669_
timestamp 1688980957
transform -1 0 18584 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0670_
timestamp 1688980957
transform 1 0 16192 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1688980957
transform 1 0 17204 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0673_
timestamp 1688980957
transform -1 0 16008 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0674_
timestamp 1688980957
transform -1 0 16008 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1688980957
transform -1 0 15732 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0677_
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0678_
timestamp 1688980957
transform -1 0 17756 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1688980957
transform -1 0 18584 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1688980957
transform 1 0 17664 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0681_
timestamp 1688980957
transform -1 0 21160 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0682_
timestamp 1688980957
transform -1 0 21160 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform -1 0 20700 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform -1 0 19964 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0685_
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0686_
timestamp 1688980957
transform -1 0 22448 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1688980957
transform 1 0 21804 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0689_
timestamp 1688980957
transform -1 0 22908 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0690_
timestamp 1688980957
transform -1 0 23460 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0693_
timestamp 1688980957
transform -1 0 26404 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0694_
timestamp 1688980957
transform -1 0 26404 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform 1 0 25576 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform 1 0 24932 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0697_
timestamp 1688980957
transform -1 0 27048 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0698_
timestamp 1688980957
transform -1 0 27508 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1688980957
transform -1 0 27784 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0701_
timestamp 1688980957
transform -1 0 31188 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0702_
timestamp 1688980957
transform -1 0 31188 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform 1 0 30176 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1688980957
transform 1 0 30084 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0705_
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0706_
timestamp 1688980957
transform -1 0 28796 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform -1 0 28980 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform 1 0 28244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0709_
timestamp 1688980957
transform -1 0 33396 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0710_
timestamp 1688980957
transform -1 0 33396 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1688980957
transform -1 0 33396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1688980957
transform -1 0 32752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0713_
timestamp 1688980957
transform 1 0 30084 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0714_
timestamp 1688980957
transform 1 0 30820 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1688980957
transform -1 0 33028 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1688980957
transform 1 0 32844 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0717_
timestamp 1688980957
transform -1 0 35328 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0718_
timestamp 1688980957
transform -1 0 34592 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1688980957
transform 1 0 35052 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform -1 0 34776 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0721_
timestamp 1688980957
transform -1 0 39744 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0722_
timestamp 1688980957
transform -1 0 39652 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1688980957
transform 1 0 37260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0725_
timestamp 1688980957
transform 1 0 36248 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0726_
timestamp 1688980957
transform -1 0 38180 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1688980957
transform -1 0 38456 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform -1 0 38548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0729_
timestamp 1688980957
transform -1 0 39744 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0730_
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1688980957
transform -1 0 40020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform 1 0 40020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0733_
timestamp 1688980957
transform -1 0 43148 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0734_
timestamp 1688980957
transform -1 0 43148 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1688980957
transform 1 0 43240 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0737_
timestamp 1688980957
transform -1 0 48024 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0738_
timestamp 1688980957
transform -1 0 48392 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1688980957
transform 1 0 48024 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform 1 0 45632 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0741_
timestamp 1688980957
transform -1 0 45448 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0742_
timestamp 1688980957
transform 1 0 42872 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform -1 0 45816 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform 1 0 45816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0745_
timestamp 1688980957
transform 1 0 42688 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0746_
timestamp 1688980957
transform -1 0 44896 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1688980957
transform -1 0 45264 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 46000 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0749_
timestamp 1688980957
transform -1 0 48024 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0750_
timestamp 1688980957
transform -1 0 49496 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1688980957
transform -1 0 48576 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform 1 0 47748 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0753_
timestamp 1688980957
transform -1 0 53268 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0754_
timestamp 1688980957
transform -1 0 52624 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 50140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0757_
timestamp 1688980957
transform -1 0 51428 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0758_
timestamp 1688980957
transform -1 0 52072 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 1688980957
transform -1 0 51612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform 1 0 50692 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0761_
timestamp 1688980957
transform -1 0 52624 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0762_
timestamp 1688980957
transform -1 0 52992 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1688980957
transform -1 0 52624 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0765_
timestamp 1688980957
transform -1 0 57316 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0766_
timestamp 1688980957
transform -1 0 57316 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 1688980957
transform 1 0 56304 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform 1 0 55384 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0769_
timestamp 1688980957
transform -1 0 57132 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0770_
timestamp 1688980957
transform -1 0 57224 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1688980957
transform 1 0 57224 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform -1 0 57040 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0773_
timestamp 1688980957
transform -1 0 57224 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0774_
timestamp 1688980957
transform -1 0 56672 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1688980957
transform -1 0 57224 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1688980957
transform 1 0 56672 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _0777_
timestamp 1688980957
transform 1 0 6164 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1688980957
transform -1 0 10764 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1688980957
transform -1 0 8004 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1688980957
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform 1 0 14628 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1688980957
transform 1 0 20884 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 23552 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1688980957
transform 1 0 24748 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1688980957
transform 1 0 28612 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1688980957
transform 1 0 25852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform 1 0 30084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1688980957
transform 1 0 30084 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1688980957
transform 1 0 32016 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1688980957
transform -1 0 38088 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1688980957
transform 1 0 36156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1688980957
transform 1 0 36064 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1688980957
transform 1 0 40204 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1688980957
transform 1 0 46092 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1688980957
transform 1 0 42688 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1688980957
transform -1 0 43056 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1688980957
transform 1 0 46460 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1688980957
transform 1 0 50416 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1688980957
transform -1 0 48668 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1688980957
transform 1 0 50232 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1688980957
transform -1 0 55108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1688980957
transform 1 0 54464 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1688980957
transform 1 0 53544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0810_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0811_
timestamp 1688980957
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0812_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0813_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0814_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3496 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0816_
timestamp 1688980957
transform -1 0 6440 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0817_
timestamp 1688980957
transform -1 0 5980 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1688980957
transform -1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0819_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3496 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0820_
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0821_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1688980957
transform -1 0 3588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0823_
timestamp 1688980957
transform -1 0 3312 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0824_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3956 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0825_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0826_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1688980957
transform 1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0828_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 1688980957
transform -1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0830_
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0831_
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0832_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43424 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0833_
timestamp 1688980957
transform -1 0 40112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0834_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 49956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0835_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 55200 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0836_
timestamp 1688980957
transform -1 0 44436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0837_
timestamp 1688980957
transform -1 0 18492 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0838_
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0839_
timestamp 1688980957
transform -1 0 24656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0840_
timestamp 1688980957
transform -1 0 30728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1688980957
transform -1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1688980957
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0843_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5520 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1688980957
transform 1 0 6256 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0847_
timestamp 1688980957
transform -1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_1  _0848_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0849_
timestamp 1688980957
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0850_
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0851_
timestamp 1688980957
transform -1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0852_
timestamp 1688980957
transform 1 0 10488 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0853_
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0854_
timestamp 1688980957
transform -1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0855_
timestamp 1688980957
transform -1 0 14168 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0856_
timestamp 1688980957
transform -1 0 15732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1688980957
transform -1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0858_
timestamp 1688980957
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0859_
timestamp 1688980957
transform -1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0860_
timestamp 1688980957
transform 1 0 18124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1688980957
transform -1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0862_
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1688980957
transform -1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0864_
timestamp 1688980957
transform -1 0 21712 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1688980957
transform -1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0866_
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1688980957
transform -1 0 21712 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0868_
timestamp 1688980957
transform -1 0 25392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform -1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0870_
timestamp 1688980957
transform -1 0 27508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1688980957
transform -1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0872_
timestamp 1688980957
transform -1 0 28796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0873_
timestamp 1688980957
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0874_
timestamp 1688980957
transform -1 0 30176 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0875_
timestamp 1688980957
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0876_
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0877_
timestamp 1688980957
transform -1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0878_
timestamp 1688980957
transform 1 0 35420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1688980957
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0880_
timestamp 1688980957
transform 1 0 35512 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1688980957
transform -1 0 34960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0882_
timestamp 1688980957
transform -1 0 38548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0883_
timestamp 1688980957
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0884_
timestamp 1688980957
transform 1 0 40112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1688980957
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0886_
timestamp 1688980957
transform -1 0 39928 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1688980957
transform -1 0 39744 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0888_
timestamp 1688980957
transform -1 0 42320 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1688980957
transform 1 0 43056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0890_
timestamp 1688980957
transform -1 0 45724 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0891_
timestamp 1688980957
transform -1 0 43608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0892_
timestamp 1688980957
transform -1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1688980957
transform -1 0 46000 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0894_
timestamp 1688980957
transform 1 0 46920 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1688980957
transform -1 0 47104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0896_
timestamp 1688980957
transform 1 0 48300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1688980957
transform -1 0 48300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0898_
timestamp 1688980957
transform 1 0 50876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1688980957
transform -1 0 49956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0900_
timestamp 1688980957
transform 1 0 51428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1688980957
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0902_
timestamp 1688980957
transform 1 0 53452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1688980957
transform 1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0904_
timestamp 1688980957
transform 1 0 56304 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0905_
timestamp 1688980957
transform -1 0 55476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0906_
timestamp 1688980957
transform -1 0 58420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1688980957
transform -1 0 56120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0908_
timestamp 1688980957
transform -1 0 57408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1688980957
transform -1 0 58604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0910_
timestamp 1688980957
transform 1 0 1840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0911_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0913_
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 1688980957
transform -1 0 2208 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0915_
timestamp 1688980957
transform 1 0 5428 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 1688980957
transform 1 0 12512 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0919_
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0921_
timestamp 1688980957
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0923_
timestamp 1688980957
transform 1 0 23092 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 1688980957
transform 1 0 24380 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 1688980957
transform 1 0 28612 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp 1688980957
transform 1 0 26128 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp 1688980957
transform -1 0 31556 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1688980957
transform 1 0 33396 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 1688980957
transform -1 0 37996 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0931_
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 1688980957
transform -1 0 37720 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp 1688980957
transform 1 0 41032 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 1688980957
transform 1 0 45632 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1688980957
transform -1 0 43240 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1688980957
transform 1 0 42228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0937_
timestamp 1688980957
transform 1 0 44988 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1688980957
transform -1 0 52072 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1688980957
transform 1 0 48668 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1688980957
transform 1 0 50140 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 1688980957
transform 1 0 54280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1688980957
transform -1 0 54740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp 1688980957
transform -1 0 55476 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0944_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1688980957
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1688980957
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 1688980957
transform 1 0 12144 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1688980957
transform 1 0 15272 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1688980957
transform 1 0 17756 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1688980957
transform -1 0 19136 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1688980957
transform 1 0 20056 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp 1688980957
transform 1 0 25392 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 1688980957
transform 1 0 28428 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0959_
timestamp 1688980957
transform 1 0 25760 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 1688980957
transform -1 0 31372 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1688980957
transform 1 0 28612 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0963_
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 1688980957
transform 1 0 35236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp 1688980957
transform 1 0 35328 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 1688980957
transform 1 0 40848 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0967_
timestamp 1688980957
transform 1 0 45172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 1688980957
transform 1 0 41860 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 1688980957
transform 1 0 46000 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1688980957
transform -1 0 50968 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 1688980957
transform 1 0 48852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1688980957
transform -1 0 51980 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp 1688980957
transform 1 0 54096 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 1688980957
transform 1 0 53636 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 1688980957
transform -1 0 55108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0977_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 1688980957
transform 1 0 11408 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 1688980957
transform -1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1688980957
transform 1 0 13156 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0983_
timestamp 1688980957
transform -1 0 16560 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp 1688980957
transform -1 0 17480 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 1688980957
transform -1 0 23368 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 1688980957
transform 1 0 25392 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1688980957
transform -1 0 26864 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 1688980957
transform 1 0 31188 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1688980957
transform 1 0 33580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1688980957
transform -1 0 30820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1688980957
transform -1 0 34316 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1688980957
transform -1 0 38916 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1688980957
transform 1 0 37536 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1688980957
transform -1 0 37720 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform -1 0 43240 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1688980957
transform -1 0 48392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1688980957
transform -1 0 43792 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1688980957
transform -1 0 44712 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 1688980957
transform -1 0 48392 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1688980957
transform -1 0 52348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1688980957
transform -1 0 50692 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1688980957
transform 1 0 52440 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1007_
timestamp 1688980957
transform 1 0 56580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1688980957
transform -1 0 57316 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1688980957
transform 1 0 57592 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1688980957
transform -1 0 9660 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 1688980957
transform -1 0 7728 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 1688980957
transform -1 0 17756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1688980957
transform 1 0 15732 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1688980957
transform -1 0 18584 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp 1688980957
transform -1 0 21252 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1688980957
transform -1 0 22724 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1020_
timestamp 1688980957
transform -1 0 24288 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1688980957
transform -1 0 27784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1022_
timestamp 1688980957
transform 1 0 27416 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 1688980957
transform 1 0 29624 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1024_
timestamp 1688980957
transform 1 0 28612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1688980957
transform -1 0 34224 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1688980957
transform -1 0 33580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1688980957
transform -1 0 35512 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1688980957
transform 1 0 40204 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1688980957
transform -1 0 39008 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp 1688980957
transform 1 0 40388 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp 1688980957
transform -1 0 43976 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1688980957
transform -1 0 49220 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1033_
timestamp 1688980957
transform -1 0 45816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1034_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 46460 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1688980957
transform 1 0 47196 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1688980957
transform -1 0 52624 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1688980957
transform -1 0 52164 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1688980957
transform 1 0 51152 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1688980957
transform 1 0 56212 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1688980957
transform 1 0 56120 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1688980957
transform 1 0 55660 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1688980957
transform 1 0 2392 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1043_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1044_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1688980957
transform 1 0 7268 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1688980957
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1688980957
transform 1 0 8372 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1688980957
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1688980957
transform -1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1688980957
transform 1 0 3956 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1688980957
transform 1 0 9844 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1688980957
transform 1 0 16744 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1688980957
transform 1 0 18768 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 22356 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform 1 0 22816 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform 1 0 27508 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform -1 0 25944 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform 1 0 29808 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 27968 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 31924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform 1 0 36340 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform 1 0 34776 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform 1 0 35420 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform 1 0 39376 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform 1 0 44160 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1688980957
transform 1 0 41676 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1688980957
transform 1 0 40848 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1688980957
transform -1 0 45632 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1688980957
transform 1 0 49220 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1688980957
transform 1 0 53544 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform 1 0 53084 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform 1 0 53452 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1688980957
transform 1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform 1 0 2208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 6348 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 12328 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform -1 0 18768 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform -1 0 15916 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1688980957
transform -1 0 22356 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform 1 0 25392 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform -1 0 26588 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1688980957
transform 1 0 29808 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1688980957
transform 1 0 24748 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1688980957
transform 1 0 32384 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1688980957
transform 1 0 29624 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1688980957
transform 1 0 38456 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1688980957
transform -1 0 37720 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1688980957
transform -1 0 41308 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1688980957
transform 1 0 41860 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1688980957
transform 1 0 46000 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1688980957
transform 1 0 43424 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1688980957
transform 1 0 42412 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1688980957
transform 1 0 46460 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1688980957
transform 1 0 52164 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1688980957
transform 1 0 50508 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1688980957
transform 1 0 56304 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1688980957
transform 1 0 56120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1688980957
transform 1 0 56212 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1688980957
transform -1 0 7820 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1688980957
transform 1 0 11592 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1688980957
transform 1 0 5704 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform 1 0 7544 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1688980957
transform -1 0 18400 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1688980957
transform -1 0 23276 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1688980957
transform -1 0 27876 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1688980957
transform 1 0 25392 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1688980957
transform -1 0 31648 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1688980957
transform -1 0 29072 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1688980957
transform -1 0 33580 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1688980957
transform 1 0 34224 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1688980957
transform 1 0 38824 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1688980957
transform -1 0 39192 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1688980957
transform 1 0 39100 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1688980957
transform 1 0 41952 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1688980957
transform -1 0 49036 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1688980957
transform -1 0 44712 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1688980957
transform 1 0 52716 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1688980957
transform 1 0 50416 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1688980957
transform -1 0 54188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1688980957
transform 1 0 56396 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1688980957
transform 1 0 56304 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1688980957
transform 1 0 56304 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1688980957
transform -1 0 7820 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1688980957
transform 1 0 8924 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1688980957
transform 1 0 9384 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1688980957
transform 1 0 12420 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1688980957
transform 1 0 14168 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1688980957
transform -1 0 19964 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1688980957
transform 1 0 21896 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1688980957
transform 1 0 24288 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1688980957
transform -1 0 30084 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1688980957
transform 1 0 27876 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1688980957
transform -1 0 33580 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1688980957
transform 1 0 32568 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1688980957
transform -1 0 34868 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1688980957
transform 1 0 37352 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1688980957
transform 1 0 38916 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1688980957
transform 1 0 40848 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1688980957
transform -1 0 45632 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1688980957
transform 1 0 45264 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1688980957
transform 1 0 45816 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1688980957
transform 1 0 47564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1688980957
transform 1 0 50140 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1688980957
transform 1 0 50232 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1688980957
transform 1 0 52164 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1688980957
transform 1 0 56764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1688980957
transform 1 0 56212 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1688980957
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp 1688980957
transform 1 0 6440 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1688980957
transform 1 0 4784 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1688980957
transform 1 0 10212 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1688980957
transform 1 0 20240 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1688980957
transform 1 0 24104 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1688980957
transform 1 0 27784 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1688980957
transform 1 0 25208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1688980957
transform 1 0 29992 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1688980957
transform 1 0 29532 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1688980957
transform 1 0 36248 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1688980957
transform 1 0 34684 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1688980957
transform 1 0 34592 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1688980957
transform 1 0 45264 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1688980957
transform 1 0 41676 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1688980957
transform 1 0 45908 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1688980957
transform 1 0 50140 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 1688980957
transform -1 0 51152 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1688980957
transform 1 0 53728 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1688980957
transform 1 0 53084 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1688980957
transform 1 0 52900 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 1688980957
transform -1 0 3036 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 1688980957
transform 1 0 2668 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 1688980957
transform 1 0 4784 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1688980957
transform -1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 1688980957
transform 1 0 14536 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1688980957
transform 1 0 15272 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp 1688980957
transform -1 0 20700 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1220_
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1221_
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp 1688980957
transform 1 0 24472 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp 1688980957
transform 1 0 25944 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1224_
timestamp 1688980957
transform 1 0 27876 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1225_
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp 1688980957
transform 1 0 31464 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp 1688980957
transform 1 0 33120 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp 1688980957
transform 1 0 34500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp 1688980957
transform 1 0 36248 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp 1688980957
transform 1 0 37904 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 1688980957
transform -1 0 42780 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1688980957
transform 1 0 43424 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1688980957
transform 1 0 45264 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1688980957
transform 1 0 46552 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1688980957
transform 1 0 47748 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1688980957
transform -1 0 53084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1688980957
transform -1 0 54556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1688980957
transform 1 0 56304 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1688980957
transform -1 0 58328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1688980957
transform -1 0 3036 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1688980957
transform 1 0 2024 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1688980957
transform 1 0 9844 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1688980957
transform -1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1688980957
transform 1 0 9936 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1688980957
transform 1 0 15364 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1688980957
transform 1 0 11960 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1688980957
transform 1 0 17296 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1688980957
transform 1 0 18768 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1688980957
transform 1 0 22448 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1688980957
transform 1 0 27876 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1688980957
transform 1 0 24656 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1688980957
transform -1 0 31464 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1688980957
transform 1 0 28428 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1688980957
transform 1 0 35236 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1688980957
transform 1 0 35696 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1688980957
transform 1 0 39560 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1688980957
transform 1 0 44804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1688980957
transform 1 0 42412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1688980957
transform 1 0 41216 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1688980957
transform 1 0 44988 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1688980957
transform 1 0 47288 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1688980957
transform 1 0 49036 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1688980957
transform 1 0 53728 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1688980957
transform 1 0 53360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1688980957
transform 1 0 53636 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1688980957
transform 1 0 5520 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1688980957
transform -1 0 5980 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1688980957
transform 1 0 15088 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1688980957
transform 1 0 13800 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1688980957
transform -1 0 19964 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1688980957
transform 1 0 19412 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1688980957
transform 1 0 23920 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1688980957
transform 1 0 27784 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1688980957
transform 1 0 29808 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1688980957
transform -1 0 29992 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1688980957
transform 1 0 31096 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1688980957
transform 1 0 36064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1688980957
transform 1 0 39376 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1688980957
transform 1 0 40848 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1688980957
transform 1 0 41400 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1688980957
transform 1 0 45448 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1688980957
transform 1 0 50140 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1688980957
transform 1 0 47380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1688980957
transform 1 0 53728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1688980957
transform 1 0 53084 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1688980957
transform 1 0 52808 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1688980957
transform -1 0 9936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1688980957
transform 1 0 9016 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1688980957
transform -1 0 8832 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1688980957
transform 1 0 12512 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1688980957
transform -1 0 17388 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1688980957
transform 1 0 13524 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1688980957
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1688980957
transform 1 0 24840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1688980957
transform -1 0 28980 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1688980957
transform 1 0 29808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1688980957
transform 1 0 27140 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1688980957
transform 1 0 29992 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1688980957
transform -1 0 35052 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1688980957
transform 1 0 38732 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1688980957
transform 1 0 36064 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1688980957
transform 1 0 36340 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1688980957
transform -1 0 49036 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1688980957
transform -1 0 44620 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1688980957
transform 1 0 42596 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1688980957
transform 1 0 47104 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1688980957
transform -1 0 53084 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1688980957
transform 1 0 49404 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1688980957
transform 1 0 50968 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1688980957
transform 1 0 56396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1688980957
transform 1 0 56304 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1688980957
transform 1 0 56120 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1688980957
transform -1 0 10396 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1688980957
transform 1 0 9200 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1688980957
transform 1 0 6348 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1688980957
transform -1 0 17940 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1688980957
transform -1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1688980957
transform 1 0 19872 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1688980957
transform 1 0 22448 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1688980957
transform -1 0 23828 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1688980957
transform 1 0 26036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1688980957
transform 1 0 27600 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1688980957
transform -1 0 33672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1688980957
transform -1 0 34224 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1688980957
transform 1 0 33764 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1688980957
transform 1 0 38916 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1688980957
transform 1 0 37444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1688980957
transform 1 0 37904 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1688980957
transform 1 0 47288 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1688980957
transform 1 0 45724 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__S
timestamp 1688980957
transform -1 0 44436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__S
timestamp 1688980957
transform 1 0 49680 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S
timestamp 1688980957
transform 1 0 51428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__S
timestamp 1688980957
transform 1 0 52256 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__S
timestamp 1688980957
transform 1 0 53176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__S
timestamp 1688980957
transform 1 0 56396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S
timestamp 1688980957
transform 1 0 57224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__S
timestamp 1688980957
transform -1 0 58328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__D
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A1
timestamp 1688980957
transform -1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1688980957
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__S
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S
timestamp 1688980957
transform 1 0 5152 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__S
timestamp 1688980957
transform 1 0 5520 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__S
timestamp 1688980957
transform 1 0 10396 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__S
timestamp 1688980957
transform 1 0 14996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__S
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__S
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__S
timestamp 1688980957
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__S
timestamp 1688980957
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__S
timestamp 1688980957
transform -1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__S
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__S
timestamp 1688980957
transform 1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__S
timestamp 1688980957
transform 1 0 27232 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__S
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__S
timestamp 1688980957
transform 1 0 29808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__S
timestamp 1688980957
transform 1 0 29808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1688980957
transform 1 0 32292 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__S
timestamp 1688980957
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1688980957
transform 1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__S
timestamp 1688980957
transform 1 0 35696 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1688980957
transform -1 0 39744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__S
timestamp 1688980957
transform 1 0 44344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__S
timestamp 1688980957
transform 1 0 42228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1688980957
transform 1 0 41308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__S
timestamp 1688980957
transform -1 0 44896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1688980957
transform 1 0 49864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__S
timestamp 1688980957
transform 1 0 47656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__S
timestamp 1688980957
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__S
timestamp 1688980957
transform 1 0 53728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1688980957
transform 1 0 53452 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__S
timestamp 1688980957
transform -1 0 53820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__S
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__S
timestamp 1688980957
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1688980957
transform 1 0 9200 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__S
timestamp 1688980957
transform 1 0 15364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1688980957
transform -1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__S
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1688980957
transform -1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__S
timestamp 1688980957
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1688980957
transform 1 0 20700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__S
timestamp 1688980957
transform 1 0 23184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1688980957
transform 1 0 24748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1688980957
transform 1 0 31188 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1688980957
transform 1 0 24656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__S
timestamp 1688980957
transform -1 0 35328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1688980957
transform 1 0 31004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1688980957
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1688980957
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__S
timestamp 1688980957
transform 1 0 36800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1688980957
transform 1 0 39192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__S
timestamp 1688980957
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1688980957
transform 1 0 47380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__S
timestamp 1688980957
transform 1 0 44988 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1688980957
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__S
timestamp 1688980957
transform 1 0 46828 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1688980957
transform 1 0 53084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__S
timestamp 1688980957
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__S
timestamp 1688980957
transform -1 0 51612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__S
timestamp 1688980957
transform 1 0 56304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__S
timestamp 1688980957
transform -1 0 56396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__S
timestamp 1688980957
transform -1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__S
timestamp 1688980957
transform -1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1688980957
transform 1 0 7912 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__S
timestamp 1688980957
transform 1 0 8832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1688980957
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__S
timestamp 1688980957
transform -1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1688980957
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__S
timestamp 1688980957
transform -1 0 17112 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1688980957
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__S
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__S
timestamp 1688980957
transform 1 0 24932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__S
timestamp 1688980957
transform 1 0 27140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1688980957
transform -1 0 31280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1688980957
transform 1 0 27140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__S
timestamp 1688980957
transform -1 0 32108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1688980957
transform 1 0 34224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__S
timestamp 1688980957
transform 1 0 35144 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1688980957
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__S
timestamp 1688980957
transform 1 0 38916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1688980957
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1688980957
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__S
timestamp 1688980957
transform 1 0 47932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1688980957
transform 1 0 45356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__S
timestamp 1688980957
transform 1 0 45172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__S
timestamp 1688980957
transform -1 0 48668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__S
timestamp 1688980957
transform 1 0 55200 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__S
timestamp 1688980957
transform 1 0 51244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__S
timestamp 1688980957
transform 1 0 52256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__S
timestamp 1688980957
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__S
timestamp 1688980957
transform 1 0 56396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__S
timestamp 1688980957
transform 1 0 56396 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__S0
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__S1
timestamp 1688980957
transform 1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__S0
timestamp 1688980957
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__S1
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__S
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__S
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__S0
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__S1
timestamp 1688980957
transform -1 0 11316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__S0
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__S1
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__S
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__S
timestamp 1688980957
transform -1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__S0
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__S1
timestamp 1688980957
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__S0
timestamp 1688980957
transform 1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__S1
timestamp 1688980957
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__S
timestamp 1688980957
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__S
timestamp 1688980957
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__S0
timestamp 1688980957
transform 1 0 8372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__S1
timestamp 1688980957
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__S0
timestamp 1688980957
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__S1
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__S
timestamp 1688980957
transform -1 0 9292 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__S
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__S0
timestamp 1688980957
transform -1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__S1
timestamp 1688980957
transform -1 0 11868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__S0
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__S1
timestamp 1688980957
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__S
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__S
timestamp 1688980957
transform -1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__S0
timestamp 1688980957
transform -1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__S1
timestamp 1688980957
transform -1 0 19136 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__S0
timestamp 1688980957
transform 1 0 16008 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__S1
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__S
timestamp 1688980957
transform 1 0 17020 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__S
timestamp 1688980957
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__S0
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__S1
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__S0
timestamp 1688980957
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__S1
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__S
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__S
timestamp 1688980957
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S0
timestamp 1688980957
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S1
timestamp 1688980957
transform -1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__S0
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__S1
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__S
timestamp 1688980957
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S0
timestamp 1688980957
transform 1 0 17112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S1
timestamp 1688980957
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S0
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S1
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__S
timestamp 1688980957
transform 1 0 19688 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__S
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S0
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S1
timestamp 1688980957
transform 1 0 22632 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S0
timestamp 1688980957
transform 1 0 20240 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S1
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__S
timestamp 1688980957
transform 1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__S
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S0
timestamp 1688980957
transform -1 0 21712 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S1
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S0
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S1
timestamp 1688980957
transform 1 0 21988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__S
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__S
timestamp 1688980957
transform 1 0 22172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S0
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S1
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S0
timestamp 1688980957
transform 1 0 24380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S1
timestamp 1688980957
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__S
timestamp 1688980957
transform 1 0 25392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__S
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S0
timestamp 1688980957
transform 1 0 25300 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S1
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S0
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S1
timestamp 1688980957
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__S
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__S
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__S0
timestamp 1688980957
transform -1 0 32384 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__S1
timestamp 1688980957
transform -1 0 31648 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S0
timestamp 1688980957
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S1
timestamp 1688980957
transform 1 0 31188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__S
timestamp 1688980957
transform 1 0 29992 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__S
timestamp 1688980957
transform 1 0 29900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S0
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S1
timestamp 1688980957
transform 1 0 26404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S0
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S1
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__S
timestamp 1688980957
transform -1 0 28152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__S
timestamp 1688980957
transform 1 0 28060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S0
timestamp 1688980957
transform -1 0 35052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S1
timestamp 1688980957
transform 1 0 34316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S0
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S1
timestamp 1688980957
transform 1 0 33580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__S
timestamp 1688980957
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__S
timestamp 1688980957
transform 1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S0
timestamp 1688980957
transform 1 0 32292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S1
timestamp 1688980957
transform 1 0 32292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S0
timestamp 1688980957
transform 1 0 33120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S1
timestamp 1688980957
transform 1 0 32752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__S
timestamp 1688980957
transform 1 0 33028 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__S
timestamp 1688980957
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S0
timestamp 1688980957
transform 1 0 35512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S1
timestamp 1688980957
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S0
timestamp 1688980957
transform 1 0 34776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S1
timestamp 1688980957
transform 1 0 34868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__S
timestamp 1688980957
transform 1 0 35604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__S
timestamp 1688980957
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S0
timestamp 1688980957
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S1
timestamp 1688980957
transform 1 0 36616 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S0
timestamp 1688980957
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S1
timestamp 1688980957
transform 1 0 38272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__S
timestamp 1688980957
transform 1 0 40020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__S
timestamp 1688980957
transform 1 0 37444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S0
timestamp 1688980957
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S1
timestamp 1688980957
transform -1 0 36248 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S0
timestamp 1688980957
transform 1 0 36892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S1
timestamp 1688980957
transform 1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__S
timestamp 1688980957
transform 1 0 38640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S0
timestamp 1688980957
transform 1 0 37444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S1
timestamp 1688980957
transform 1 0 37812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S0
timestamp 1688980957
transform 1 0 38640 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S1
timestamp 1688980957
transform 1 0 37076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1688980957
transform 1 0 39008 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__S
timestamp 1688980957
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S0
timestamp 1688980957
transform -1 0 41032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S1
timestamp 1688980957
transform 1 0 41216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S0
timestamp 1688980957
transform 1 0 41124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S1
timestamp 1688980957
transform 1 0 41492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__S
timestamp 1688980957
transform 1 0 43332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__S
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S0
timestamp 1688980957
transform 1 0 49036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S1
timestamp 1688980957
transform 1 0 48208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S0
timestamp 1688980957
transform 1 0 49312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S1
timestamp 1688980957
transform 1 0 48944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__S
timestamp 1688980957
transform 1 0 47840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__S
timestamp 1688980957
transform 1 0 46644 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S0
timestamp 1688980957
transform 1 0 44160 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S1
timestamp 1688980957
transform 1 0 44528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S0
timestamp 1688980957
transform 1 0 44988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S1
timestamp 1688980957
transform 1 0 44988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__S
timestamp 1688980957
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1688980957
transform 1 0 45908 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S0
timestamp 1688980957
transform 1 0 45264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S1
timestamp 1688980957
transform 1 0 44896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S0
timestamp 1688980957
transform 1 0 45540 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S1
timestamp 1688980957
transform 1 0 45172 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S
timestamp 1688980957
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1688980957
transform 1 0 45816 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__S0
timestamp 1688980957
transform 1 0 48576 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__S1
timestamp 1688980957
transform -1 0 48392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S0
timestamp 1688980957
transform 1 0 45724 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S1
timestamp 1688980957
transform 1 0 49680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S
timestamp 1688980957
transform 1 0 47564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__S
timestamp 1688980957
transform -1 0 47472 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S0
timestamp 1688980957
transform 1 0 50232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S1
timestamp 1688980957
transform -1 0 52440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S0
timestamp 1688980957
transform 1 0 50324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S1
timestamp 1688980957
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S
timestamp 1688980957
transform 1 0 52624 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1688980957
transform 1 0 49956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S0
timestamp 1688980957
transform 1 0 49220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S1
timestamp 1688980957
transform 1 0 49680 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S0
timestamp 1688980957
transform 1 0 50324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S1
timestamp 1688980957
transform 1 0 50692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S
timestamp 1688980957
transform 1 0 50600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__S
timestamp 1688980957
transform 1 0 50508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S0
timestamp 1688980957
transform -1 0 50508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S1
timestamp 1688980957
transform 1 0 49864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S0
timestamp 1688980957
transform 1 0 50692 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S1
timestamp 1688980957
transform 1 0 52164 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__S
timestamp 1688980957
transform -1 0 52348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp 1688980957
transform 1 0 52440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S0
timestamp 1688980957
transform 1 0 55200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S1
timestamp 1688980957
transform 1 0 55476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S0
timestamp 1688980957
transform 1 0 55016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S1
timestamp 1688980957
transform 1 0 55384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__S
timestamp 1688980957
transform 1 0 56120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp 1688980957
transform 1 0 55200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S0
timestamp 1688980957
transform 1 0 54832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S1
timestamp 1688980957
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S0
timestamp 1688980957
transform 1 0 54924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S1
timestamp 1688980957
transform 1 0 55476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp 1688980957
transform -1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp 1688980957
transform 1 0 55292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S0
timestamp 1688980957
transform 1 0 54924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S1
timestamp 1688980957
transform 1 0 55476 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S0
timestamp 1688980957
transform 1 0 54372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S1
timestamp 1688980957
transform 1 0 54740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S
timestamp 1688980957
transform 1 0 56212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__S
timestamp 1688980957
transform -1 0 56120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S
timestamp 1688980957
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__S
timestamp 1688980957
transform 1 0 8464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__S
timestamp 1688980957
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S
timestamp 1688980957
transform 1 0 11684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S
timestamp 1688980957
transform 1 0 14720 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp 1688980957
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S
timestamp 1688980957
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S
timestamp 1688980957
transform 1 0 18124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1688980957
transform -1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp 1688980957
transform 1 0 23368 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S
timestamp 1688980957
transform 1 0 23920 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S
timestamp 1688980957
transform -1 0 28612 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S
timestamp 1688980957
transform 1 0 31832 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp 1688980957
transform 1 0 31832 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__S
timestamp 1688980957
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__S
timestamp 1688980957
transform -1 0 36340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S
timestamp 1688980957
transform 1 0 35880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__S
timestamp 1688980957
transform 1 0 40020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__S
timestamp 1688980957
transform 1 0 47104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__S
timestamp 1688980957
transform 1 0 42596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__S
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__S
timestamp 1688980957
transform 1 0 46276 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__S
timestamp 1688980957
transform -1 0 50416 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__S
timestamp 1688980957
transform 1 0 47656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__S
timestamp 1688980957
transform 1 0 49128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__S
timestamp 1688980957
transform 1 0 54096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__S
timestamp 1688980957
transform 1 0 54740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__S
timestamp 1688980957
transform -1 0 54740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A_N
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A_N
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A_N
timestamp 1688980957
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A1
timestamp 1688980957
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__D
timestamp 1688980957
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A2
timestamp 1688980957
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B1
timestamp 1688980957
transform 1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B1
timestamp 1688980957
transform -1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2
timestamp 1688980957
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B1
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1688980957
transform 1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1
timestamp 1688980957
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A2
timestamp 1688980957
transform 1 0 14996 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A2
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B1
timestamp 1688980957
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1688980957
transform 1 0 16744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1688980957
transform -1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1688980957
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A2
timestamp 1688980957
transform -1 0 19596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B1
timestamp 1688980957
transform -1 0 19964 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1688980957
transform 1 0 20516 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A2
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B1
timestamp 1688980957
transform -1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A2
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B1
timestamp 1688980957
transform 1 0 21528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1688980957
transform 1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A2
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B1
timestamp 1688980957
transform 1 0 24840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1688980957
transform 1 0 26772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1688980957
transform 1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A2
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1688980957
transform 1 0 27416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1688980957
transform 1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1688980957
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1688980957
transform -1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1688980957
transform -1 0 32016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B1
timestamp 1688980957
transform 1 0 31004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1688980957
transform 1 0 31556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1688980957
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1688980957
transform -1 0 39744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1688980957
transform 1 0 40296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A2
timestamp 1688980957
transform 1 0 36156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B1
timestamp 1688980957
transform 1 0 37536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1688980957
transform 1 0 35512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A2
timestamp 1688980957
transform 1 0 40848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B1
timestamp 1688980957
transform 1 0 41216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1688980957
transform 1 0 39008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A2
timestamp 1688980957
transform 1 0 41308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B1
timestamp 1688980957
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1688980957
transform 1 0 40664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A2
timestamp 1688980957
transform 1 0 43700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B1
timestamp 1688980957
transform -1 0 39376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1688980957
transform -1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A2
timestamp 1688980957
transform 1 0 45172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B1
timestamp 1688980957
transform 1 0 45540 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1688980957
transform 1 0 44620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A2
timestamp 1688980957
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B1
timestamp 1688980957
transform 1 0 45172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1688980957
transform 1 0 45908 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A2
timestamp 1688980957
transform 1 0 46460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B1
timestamp 1688980957
transform 1 0 46828 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1688980957
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A2
timestamp 1688980957
transform 1 0 47380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1
timestamp 1688980957
transform 1 0 48484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1688980957
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1688980957
transform 1 0 48852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1688980957
transform 1 0 48576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1688980957
transform 1 0 48208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1688980957
transform 1 0 52900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1688980957
transform 1 0 50324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1688980957
transform 1 0 49496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1688980957
transform 1 0 51796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1688980957
transform 1 0 49588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1688980957
transform 1 0 52164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A2
timestamp 1688980957
transform 1 0 53728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B1
timestamp 1688980957
transform 1 0 54556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1688980957
transform 1 0 55016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A2
timestamp 1688980957
transform 1 0 55016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B1
timestamp 1688980957
transform 1 0 54464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1688980957
transform 1 0 55016 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1688980957
transform -1 0 57408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B1
timestamp 1688980957
transform 1 0 56488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1688980957
transform 1 0 54832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A2
timestamp 1688980957
transform -1 0 54280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B1
timestamp 1688980957
transform 1 0 54648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1688980957
transform -1 0 55108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__S
timestamp 1688980957
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__S
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__S
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__S
timestamp 1688980957
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__S
timestamp 1688980957
transform 1 0 11684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__S
timestamp 1688980957
transform 1 0 14996 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__S
timestamp 1688980957
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__S
timestamp 1688980957
transform -1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__S
timestamp 1688980957
transform 1 0 17848 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__S
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__S
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__S
timestamp 1688980957
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__S
timestamp 1688980957
transform 1 0 23920 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__S
timestamp 1688980957
transform 1 0 27600 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__S
timestamp 1688980957
transform -1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__S
timestamp 1688980957
transform 1 0 31740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__S
timestamp 1688980957
transform 1 0 29992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__S
timestamp 1688980957
transform 1 0 33764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__S
timestamp 1688980957
transform 1 0 36984 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__S
timestamp 1688980957
transform 1 0 39192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__S
timestamp 1688980957
transform 1 0 36892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__S
timestamp 1688980957
transform 1 0 41032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__S
timestamp 1688980957
transform 1 0 45356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__S
timestamp 1688980957
transform 1 0 41860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__S
timestamp 1688980957
transform 1 0 42044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__S
timestamp 1688980957
transform 1 0 44712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__S
timestamp 1688980957
transform -1 0 51980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__S
timestamp 1688980957
transform 1 0 49680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__S
timestamp 1688980957
transform -1 0 50140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__S
timestamp 1688980957
transform 1 0 54096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__S
timestamp 1688980957
transform 1 0 53728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__S
timestamp 1688980957
transform -1 0 54924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__S
timestamp 1688980957
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__S
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__S
timestamp 1688980957
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__S
timestamp 1688980957
transform -1 0 5336 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__S
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__S
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__S
timestamp 1688980957
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__S
timestamp 1688980957
transform -1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__S
timestamp 1688980957
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__S
timestamp 1688980957
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__S
timestamp 1688980957
transform 1 0 19688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__S
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__S
timestamp 1688980957
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__S
timestamp 1688980957
transform 1 0 28244 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__S
timestamp 1688980957
transform 1 0 24840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__S
timestamp 1688980957
transform 1 0 31556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__S
timestamp 1688980957
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__S
timestamp 1688980957
transform 1 0 31924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__S
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__S
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__S
timestamp 1688980957
transform 1 0 35144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__S
timestamp 1688980957
transform 1 0 41860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__S
timestamp 1688980957
transform 1 0 46184 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__S
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__S
timestamp 1688980957
transform 1 0 41400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__S
timestamp 1688980957
transform -1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__S
timestamp 1688980957
transform 1 0 50324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__S
timestamp 1688980957
transform 1 0 49220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__S
timestamp 1688980957
transform -1 0 51152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__S
timestamp 1688980957
transform 1 0 53912 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__S
timestamp 1688980957
transform 1 0 53452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__S
timestamp 1688980957
transform -1 0 55660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__C
timestamp 1688980957
transform -1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__S
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__S
timestamp 1688980957
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__S
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__S
timestamp 1688980957
transform 1 0 9936 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__S
timestamp 1688980957
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__S
timestamp 1688980957
transform 1 0 15548 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__S
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__S
timestamp 1688980957
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__S
timestamp 1688980957
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__S
timestamp 1688980957
transform 1 0 20700 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__S
timestamp 1688980957
transform -1 0 22540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__S
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__S
timestamp 1688980957
transform 1 0 25852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__S
timestamp 1688980957
transform 1 0 31280 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__S
timestamp 1688980957
transform -1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__S
timestamp 1688980957
transform -1 0 34592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__S
timestamp 1688980957
transform 1 0 29808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__S
timestamp 1688980957
transform 1 0 33304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__S
timestamp 1688980957
transform 1 0 38640 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__S
timestamp 1688980957
transform 1 0 37444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__S
timestamp 1688980957
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__S
timestamp 1688980957
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__S
timestamp 1688980957
transform 1 0 47932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__S
timestamp 1688980957
transform 1 0 42136 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__S
timestamp 1688980957
transform 1 0 43700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__S
timestamp 1688980957
transform -1 0 47932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__S
timestamp 1688980957
transform 1 0 49864 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__S
timestamp 1688980957
transform 1 0 49680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__S
timestamp 1688980957
transform 1 0 53452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__S
timestamp 1688980957
transform -1 0 57776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__S
timestamp 1688980957
transform 1 0 56304 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__S
timestamp 1688980957
transform -1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__S
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__S
timestamp 1688980957
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__S
timestamp 1688980957
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__S
timestamp 1688980957
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__S
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__S
timestamp 1688980957
transform 1 0 17020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__S
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__S
timestamp 1688980957
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__S
timestamp 1688980957
transform 1 0 20240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__S
timestamp 1688980957
transform -1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__S
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__S
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__S
timestamp 1688980957
transform 1 0 27140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__S
timestamp 1688980957
transform 1 0 29440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__S
timestamp 1688980957
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__S
timestamp 1688980957
transform -1 0 34500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__S
timestamp 1688980957
transform 1 0 33764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__S
timestamp 1688980957
transform 1 0 35696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__S
timestamp 1688980957
transform 1 0 40020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__S
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__S
timestamp 1688980957
transform 1 0 41768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__S
timestamp 1688980957
transform -1 0 43148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__S
timestamp 1688980957
transform 1 0 48576 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__S
timestamp 1688980957
transform 1 0 45540 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__CLK
timestamp 1688980957
transform 1 0 55936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__CLK
timestamp 1688980957
transform -1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__CLK
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__CLK
timestamp 1688980957
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__CLK
timestamp 1688980957
transform 1 0 29716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1688980957
transform 1 0 27508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1688980957
transform 1 0 31280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__CLK
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1688980957
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1688980957
transform -1 0 33764 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1688980957
transform 1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1688980957
transform 1 0 25944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1688980957
transform 1 0 32660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1688980957
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1688980957
transform -1 0 45540 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1688980957
transform 1 0 50048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1688980957
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1688980957
transform 1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1688980957
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1688980957
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1688980957
transform -1 0 36432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1688980957
transform 1 0 41308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1688980957
transform -1 0 45264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1688980957
transform 1 0 43332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1688980957
transform 1 0 52900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1688980957
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1688980957
transform 1 0 29992 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__CLK
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__CLK
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__CLK
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__CLK
timestamp 1688980957
transform -1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 1688980957
transform -1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 1688980957
transform 1 0 29716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 1688980957
transform 1 0 34868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 1688980957
transform 1 0 36892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__CLK
timestamp 1688980957
transform 1 0 39284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__CLK
timestamp 1688980957
transform -1 0 46920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__CLK
timestamp 1688980957
transform 1 0 42596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 1688980957
transform 1 0 47196 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 1688980957
transform 1 0 52900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 1688980957
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__CLK
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__CLK
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 1688980957
transform 1 0 23736 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__CLK
timestamp 1688980957
transform 1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__CLK
timestamp 1688980957
transform 1 0 32660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__CLK
timestamp 1688980957
transform 1 0 35880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__CLK
timestamp 1688980957
transform 1 0 38456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1688980957
transform 1 0 44068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__CLK
timestamp 1688980957
transform 1 0 46736 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1688980957
transform 1 0 45172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1688980957
transform 1 0 49864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1688980957
transform -1 0 10948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1688980957
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__CLK
timestamp 1688980957
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1688980957
transform 1 0 30084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1688980957
transform 1 0 39100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1688980957
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1688980957
transform 1 0 44436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1688980957
transform 1 0 46828 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1688980957
transform 1 0 46276 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_wb_clk_i_A
timestamp 1688980957
transform -1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_wb_clk_i_A
timestamp 1688980957
transform -1 0 41584 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1688980957
transform 1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1688980957
transform -1 0 25208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1688980957
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1688980957
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1688980957
transform 1 0 41492 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1688980957
transform 1 0 50600 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1688980957
transform 1 0 52900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1688980957
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1688980957
transform 1 0 43700 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1688980957
transform 1 0 53176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1688980957
transform 1 0 49128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1688980957
transform 1 0 41584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1688980957
transform 1 0 36616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1688980957
transform 1 0 27140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform -1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform -1 0 8832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform -1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1688980957
transform -1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1688980957
transform 1 0 29808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 1688980957
transform -1 0 34500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 1688980957
transform -1 0 11960 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 1688980957
transform 1 0 32292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_A
timestamp 1688980957
transform -1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 1688980957
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 1688980957
transform -1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1688980957
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp 1688980957
transform -1 0 8372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 1688980957
transform -1 0 35788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_A
timestamp 1688980957
transform -1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1688980957
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1688980957
transform 1 0 47104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1688980957
transform 1 0 32568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout130_A
timestamp 1688980957
transform -1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout131_A
timestamp 1688980957
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout132_A
timestamp 1688980957
transform 1 0 46276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout133_A
timestamp 1688980957
transform 1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout135_A
timestamp 1688980957
transform -1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout136_A
timestamp 1688980957
transform 1 0 37168 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout137_A
timestamp 1688980957
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout138_A
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout139_A
timestamp 1688980957
transform 1 0 31372 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 20056 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1688980957
transform -1 0 8832 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1688980957
transform 1 0 25208 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1688980957
transform 1 0 25576 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1688980957
transform 1 0 35144 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1688980957
transform -1 0 52624 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1688980957
transform 1 0 52808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1688980957
transform 1 0 43884 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1688980957
transform 1 0 53360 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1688980957
transform -1 0 51980 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1688980957
transform 1 0 39284 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1688980957
transform -1 0 36616 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1688980957
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1688980957
transform -1 0 23920 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1688980957
transform 1 0 9292 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout102 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout103
timestamp 1688980957
transform 1 0 11684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout104
timestamp 1688980957
transform 1 0 32752 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout105
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout106 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13800 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout107
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout108
timestamp 1688980957
transform 1 0 8648 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout109
timestamp 1688980957
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout110 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout111
timestamp 1688980957
transform 1 0 36064 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout113
timestamp 1688980957
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout114
timestamp 1688980957
transform -1 0 7912 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout115
timestamp 1688980957
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout116
timestamp 1688980957
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout117
timestamp 1688980957
transform 1 0 33396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout118
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout119
timestamp 1688980957
transform 1 0 30820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout120
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout121
timestamp 1688980957
transform 1 0 33672 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout122
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout123
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout124
timestamp 1688980957
transform 1 0 33580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout125 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout126
timestamp 1688980957
transform 1 0 16744 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout127
timestamp 1688980957
transform 1 0 47288 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout128
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout129
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout130
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout131
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout132
timestamp 1688980957
transform 1 0 46368 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout133
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout134
timestamp 1688980957
transform -1 0 9016 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout135
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout136
timestamp 1688980957
transform 1 0 34592 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout137
timestamp 1688980957
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout138
timestamp 1688980957
transform 1 0 4784 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout139
timestamp 1688980957
transform -1 0 33488 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_340
timestamp 1688980957
transform 1 0 32384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_536
timestamp 1688980957
transform 1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_558
timestamp 1688980957
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_609
timestamp 1688980957
transform 1 0 57132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_80 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_213
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_233
timestamp 1688980957
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_275
timestamp 1688980957
transform 1 0 26404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_321
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_355
timestamp 1688980957
transform 1 0 33764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_370
timestamp 1688980957
transform 1 0 35144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_379
timestamp 1688980957
transform 1 0 35972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_386
timestamp 1688980957
transform 1 0 36616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_411
timestamp 1688980957
transform 1 0 38916 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_415
timestamp 1688980957
transform 1 0 39284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_430
timestamp 1688980957
transform 1 0 40664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_497
timestamp 1688980957
transform 1 0 46828 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_519
timestamp 1688980957
transform 1 0 48852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_545
timestamp 1688980957
transform 1 0 51244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_553
timestamp 1688980957
transform 1 0 51980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1688980957
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_599
timestamp 1688980957
transform 1 0 56212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_101
timestamp 1688980957
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_148
timestamp 1688980957
transform 1 0 14720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_152
timestamp 1688980957
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_170
timestamp 1688980957
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_216
timestamp 1688980957
transform 1 0 20976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_286
timestamp 1688980957
transform 1 0 27416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_325
timestamp 1688980957
transform 1 0 31004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_346
timestamp 1688980957
transform 1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_398
timestamp 1688980957
transform 1 0 37720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_416
timestamp 1688980957
transform 1 0 39376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_453
timestamp 1688980957
transform 1 0 42780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_496
timestamp 1688980957
transform 1 0 46736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_501
timestamp 1688980957
transform 1 0 47196 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_505
timestamp 1688980957
transform 1 0 47564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1688980957
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_605
timestamp 1688980957
transform 1 0 56764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_30
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_71
timestamp 1688980957
transform 1 0 7636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_92
timestamp 1688980957
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_108
timestamp 1688980957
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_121
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_183
timestamp 1688980957
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_199
timestamp 1688980957
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_208
timestamp 1688980957
transform 1 0 20240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_256
timestamp 1688980957
transform 1 0 24656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_284
timestamp 1688980957
transform 1 0 27232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_288
timestamp 1688980957
transform 1 0 27600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_309
timestamp 1688980957
transform 1 0 29532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_325
timestamp 1688980957
transform 1 0 31004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_379
timestamp 1688980957
transform 1 0 35972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_389
timestamp 1688980957
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_430
timestamp 1688980957
transform 1 0 40664 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_434
timestamp 1688980957
transform 1 0 41032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_457
timestamp 1688980957
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_496
timestamp 1688980957
transform 1 0 46736 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_505
timestamp 1688980957
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_509
timestamp 1688980957
transform 1 0 47932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_513
timestamp 1688980957
transform 1 0 48300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_517
timestamp 1688980957
transform 1 0 48668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_521
timestamp 1688980957
transform 1 0 49036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_531
timestamp 1688980957
transform 1 0 49956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_547
timestamp 1688980957
transform 1 0 51428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_561
timestamp 1688980957
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_565
timestamp 1688980957
transform 1 0 53084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_584
timestamp 1688980957
transform 1 0 54832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_591
timestamp 1688980957
transform 1 0 55476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_13
timestamp 1688980957
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_17
timestamp 1688980957
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_44
timestamp 1688980957
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_55
timestamp 1688980957
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_60
timestamp 1688980957
transform 1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_64
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_68
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_72
timestamp 1688980957
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_95
timestamp 1688980957
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_106
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_111
timestamp 1688980957
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_115
timestamp 1688980957
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_131
timestamp 1688980957
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_136
timestamp 1688980957
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_149
timestamp 1688980957
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_164
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_168
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_172
timestamp 1688980957
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_201
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_205
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_216
timestamp 1688980957
transform 1 0 20976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_220
timestamp 1688980957
transform 1 0 21344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_224
timestamp 1688980957
transform 1 0 21712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_248
timestamp 1688980957
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_256
timestamp 1688980957
transform 1 0 24656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_260
timestamp 1688980957
transform 1 0 25024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_264
timestamp 1688980957
transform 1 0 25392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_281
timestamp 1688980957
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_287
timestamp 1688980957
transform 1 0 27508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_291
timestamp 1688980957
transform 1 0 27876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_304
timestamp 1688980957
transform 1 0 29072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_319 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_327
timestamp 1688980957
transform 1 0 31188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_331
timestamp 1688980957
transform 1 0 31556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_386
timestamp 1688980957
transform 1 0 36616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_390
timestamp 1688980957
transform 1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_394
timestamp 1688980957
transform 1 0 37352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_407
timestamp 1688980957
transform 1 0 38548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_416
timestamp 1688980957
transform 1 0 39376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_424
timestamp 1688980957
transform 1 0 40112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_428
timestamp 1688980957
transform 1 0 40480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_465
timestamp 1688980957
transform 1 0 43884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_481
timestamp 1688980957
transform 1 0 45356 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_485
timestamp 1688980957
transform 1 0 45724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_489
timestamp 1688980957
transform 1 0 46092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_493
timestamp 1688980957
transform 1 0 46460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_510
timestamp 1688980957
transform 1 0 48024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_514
timestamp 1688980957
transform 1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_518
timestamp 1688980957
transform 1 0 48760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_524
timestamp 1688980957
transform 1 0 49312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1688980957
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_553
timestamp 1688980957
transform 1 0 51980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_579
timestamp 1688980957
transform 1 0 54372 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_583
timestamp 1688980957
transform 1 0 54740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_589
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_598
timestamp 1688980957
transform 1 0 56120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_608
timestamp 1688980957
transform 1 0 57040 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_38
timestamp 1688980957
transform 1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_43
timestamp 1688980957
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_47
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_150
timestamp 1688980957
transform 1 0 14904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_201
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_211
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 1688980957
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_240
timestamp 1688980957
transform 1 0 23184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_244
timestamp 1688980957
transform 1 0 23552 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_248
timestamp 1688980957
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_260
timestamp 1688980957
transform 1 0 25024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_274
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_289
timestamp 1688980957
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_307
timestamp 1688980957
transform 1 0 29348 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_333
timestamp 1688980957
transform 1 0 31740 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_368
timestamp 1688980957
transform 1 0 34960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_372
timestamp 1688980957
transform 1 0 35328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_376
timestamp 1688980957
transform 1 0 35696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_382
timestamp 1688980957
transform 1 0 36248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_388
timestamp 1688980957
transform 1 0 36800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_410
timestamp 1688980957
transform 1 0 38824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_414
timestamp 1688980957
transform 1 0 39192 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_435
timestamp 1688980957
transform 1 0 41124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_439
timestamp 1688980957
transform 1 0 41492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_458
timestamp 1688980957
transform 1 0 43240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_493
timestamp 1688980957
transform 1 0 46460 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_500
timestamp 1688980957
transform 1 0 47104 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_513
timestamp 1688980957
transform 1 0 48300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_525
timestamp 1688980957
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_529
timestamp 1688980957
transform 1 0 49772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_533
timestamp 1688980957
transform 1 0 50140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_545
timestamp 1688980957
transform 1 0 51244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_549
timestamp 1688980957
transform 1 0 51612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_556
timestamp 1688980957
transform 1 0 52256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_570
timestamp 1688980957
transform 1 0 53544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_574
timestamp 1688980957
transform 1 0 53912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_578
timestamp 1688980957
transform 1 0 54280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_582
timestamp 1688980957
transform 1 0 54648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_586
timestamp 1688980957
transform 1 0 55016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_599
timestamp 1688980957
transform 1 0 56212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_19
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_49
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_59
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_76
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_136
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_188
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_201
timestamp 1688980957
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_229
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_238
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_242
timestamp 1688980957
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1688980957
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303
timestamp 1688980957
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_317
timestamp 1688980957
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_328
timestamp 1688980957
transform 1 0 31280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_334
timestamp 1688980957
transform 1 0 31832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_337
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_359
timestamp 1688980957
transform 1 0 34132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_369
timestamp 1688980957
transform 1 0 35052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_411
timestamp 1688980957
transform 1 0 38916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_415
timestamp 1688980957
transform 1 0 39284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_429
timestamp 1688980957
transform 1 0 40572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_434
timestamp 1688980957
transform 1 0 41032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_438
timestamp 1688980957
transform 1 0 41400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_442
timestamp 1688980957
transform 1 0 41768 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_467
timestamp 1688980957
transform 1 0 44068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_471
timestamp 1688980957
transform 1 0 44436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_481
timestamp 1688980957
transform 1 0 45356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_491
timestamp 1688980957
transform 1 0 46276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_495
timestamp 1688980957
transform 1 0 46644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_499
timestamp 1688980957
transform 1 0 47012 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_505
timestamp 1688980957
transform 1 0 47564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_517
timestamp 1688980957
transform 1 0 48668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_523
timestamp 1688980957
transform 1 0 49220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_551
timestamp 1688980957
transform 1 0 51796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_557
timestamp 1688980957
transform 1 0 52348 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_568
timestamp 1688980957
transform 1 0 53360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_580
timestamp 1688980957
transform 1 0 54464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_584
timestamp 1688980957
transform 1 0 54832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_621
timestamp 1688980957
transform 1 0 58236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_24
timestamp 1688980957
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_64
timestamp 1688980957
transform 1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_89
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_140
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_194
timestamp 1688980957
transform 1 0 18952 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1688980957
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_289
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_294
timestamp 1688980957
transform 1 0 28152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_298
timestamp 1688980957
transform 1 0 28520 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_303
timestamp 1688980957
transform 1 0 28980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_315
timestamp 1688980957
transform 1 0 30084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_321
timestamp 1688980957
transform 1 0 30636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_331
timestamp 1688980957
transform 1 0 31556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_364
timestamp 1688980957
transform 1 0 34592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_386
timestamp 1688980957
transform 1 0 36616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_390
timestamp 1688980957
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_402
timestamp 1688980957
transform 1 0 38088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_412
timestamp 1688980957
transform 1 0 39008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_444
timestamp 1688980957
transform 1 0 41952 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_466
timestamp 1688980957
transform 1 0 43976 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_478
timestamp 1688980957
transform 1 0 45080 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_486
timestamp 1688980957
transform 1 0 45816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_514
timestamp 1688980957
transform 1 0 48392 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_520
timestamp 1688980957
transform 1 0 48944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_553
timestamp 1688980957
transform 1 0 51980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_557
timestamp 1688980957
transform 1 0 52348 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_573
timestamp 1688980957
transform 1 0 53820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_578
timestamp 1688980957
transform 1 0 54280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_584
timestamp 1688980957
transform 1 0 54832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_587
timestamp 1688980957
transform 1 0 55108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_89
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_94
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_127
timestamp 1688980957
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_131
timestamp 1688980957
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_154
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_213
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_246
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_270
timestamp 1688980957
transform 1 0 25944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_303
timestamp 1688980957
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_313
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_373
timestamp 1688980957
transform 1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_381
timestamp 1688980957
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_403
timestamp 1688980957
transform 1 0 38180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_407
timestamp 1688980957
transform 1 0 38548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_417
timestamp 1688980957
transform 1 0 39468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_432
timestamp 1688980957
transform 1 0 40848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_465
timestamp 1688980957
transform 1 0 43884 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1688980957
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_495
timestamp 1688980957
transform 1 0 46644 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_499
timestamp 1688980957
transform 1 0 47012 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_524
timestamp 1688980957
transform 1 0 49312 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_537
timestamp 1688980957
transform 1 0 50508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_576
timestamp 1688980957
transform 1 0 54096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_585
timestamp 1688980957
transform 1 0 54924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_600
timestamp 1688980957
transform 1 0 56304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_608
timestamp 1688980957
transform 1 0 57040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_616
timestamp 1688980957
transform 1 0 57776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_623
timestamp 1688980957
transform 1 0 58420 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_63
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_92
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_98
timestamp 1688980957
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_163
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_188
timestamp 1688980957
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_192
timestamp 1688980957
transform 1 0 18768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_212
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_250
timestamp 1688980957
transform 1 0 24104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_285
timestamp 1688980957
transform 1 0 27324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_377
timestamp 1688980957
transform 1 0 35788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_389
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_406
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_410
timestamp 1688980957
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_416
timestamp 1688980957
transform 1 0 39376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_443
timestamp 1688980957
transform 1 0 41860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_467
timestamp 1688980957
transform 1 0 44068 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_501
timestamp 1688980957
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_505
timestamp 1688980957
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_510
timestamp 1688980957
transform 1 0 48024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_514
timestamp 1688980957
transform 1 0 48392 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_522
timestamp 1688980957
transform 1 0 49128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_539
timestamp 1688980957
transform 1 0 50692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_549
timestamp 1688980957
transform 1 0 51612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_577
timestamp 1688980957
transform 1 0 54188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_595
timestamp 1688980957
transform 1 0 55844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_609
timestamp 1688980957
transform 1 0 57132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_613
timestamp 1688980957
transform 1 0 57500 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_34
timestamp 1688980957
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_38
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_50
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_63
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_166
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_218
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_224
timestamp 1688980957
transform 1 0 21712 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_236
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_280
timestamp 1688980957
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_302
timestamp 1688980957
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_414
timestamp 1688980957
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_418
timestamp 1688980957
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_427
timestamp 1688980957
transform 1 0 40388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_468
timestamp 1688980957
transform 1 0 44160 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_486
timestamp 1688980957
transform 1 0 45816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_519
timestamp 1688980957
transform 1 0 48852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_523
timestamp 1688980957
transform 1 0 49220 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_529
timestamp 1688980957
transform 1 0 49772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_567
timestamp 1688980957
transform 1 0 53268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_571
timestamp 1688980957
transform 1 0 53636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_597
timestamp 1688980957
transform 1 0 56028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_31
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_35
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_67
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_95
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_142
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_146
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_150
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_158
timestamp 1688980957
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_213
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_244
timestamp 1688980957
transform 1 0 23552 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_274
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_289
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_297
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_331
timestamp 1688980957
transform 1 0 31556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_341
timestamp 1688980957
transform 1 0 32476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_355
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_371
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_397
timestamp 1688980957
transform 1 0 37628 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_423
timestamp 1688980957
transform 1 0 40020 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_435
timestamp 1688980957
transform 1 0 41124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_491
timestamp 1688980957
transform 1 0 46276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_521
timestamp 1688980957
transform 1 0 49036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_529
timestamp 1688980957
transform 1 0 49772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_538
timestamp 1688980957
transform 1 0 50600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_544
timestamp 1688980957
transform 1 0 51152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_548
timestamp 1688980957
transform 1 0 51520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_553
timestamp 1688980957
transform 1 0 51980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_558
timestamp 1688980957
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_586
timestamp 1688980957
transform 1 0 55016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_611
timestamp 1688980957
transform 1 0 57316 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_35
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_39
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_66
timestamp 1688980957
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_75
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_94
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_164
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_176
timestamp 1688980957
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_186
timestamp 1688980957
transform 1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_212
timestamp 1688980957
transform 1 0 20608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_225
timestamp 1688980957
transform 1 0 21804 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_242
timestamp 1688980957
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_246
timestamp 1688980957
transform 1 0 23736 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1688980957
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_313
timestamp 1688980957
transform 1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_317
timestamp 1688980957
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_329
timestamp 1688980957
transform 1 0 31372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_341
timestamp 1688980957
transform 1 0 32476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_351
timestamp 1688980957
transform 1 0 33396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_355
timestamp 1688980957
transform 1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_359
timestamp 1688980957
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_369
timestamp 1688980957
transform 1 0 35052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_379
timestamp 1688980957
transform 1 0 35972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_391
timestamp 1688980957
transform 1 0 37076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_400
timestamp 1688980957
transform 1 0 37904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_404
timestamp 1688980957
transform 1 0 38272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_409
timestamp 1688980957
transform 1 0 38732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_453
timestamp 1688980957
transform 1 0 42780 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_501
timestamp 1688980957
transform 1 0 47196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_530
timestamp 1688980957
transform 1 0 49864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_557
timestamp 1688980957
transform 1 0 52348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_565
timestamp 1688980957
transform 1 0 53084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_589
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_133
timestamp 1688980957
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_163
timestamp 1688980957
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_185
timestamp 1688980957
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_229
timestamp 1688980957
transform 1 0 22172 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_255
timestamp 1688980957
transform 1 0 24564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_259
timestamp 1688980957
transform 1 0 24932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_276
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_285
timestamp 1688980957
transform 1 0 27324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_345
timestamp 1688980957
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_397
timestamp 1688980957
transform 1 0 37628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_415
timestamp 1688980957
transform 1 0 39284 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_423
timestamp 1688980957
transform 1 0 40020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_433
timestamp 1688980957
transform 1 0 40940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_437
timestamp 1688980957
transform 1 0 41308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_441
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_445
timestamp 1688980957
transform 1 0 42044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_458
timestamp 1688980957
transform 1 0 43240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_467
timestamp 1688980957
transform 1 0 44068 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_475
timestamp 1688980957
transform 1 0 44804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_480
timestamp 1688980957
transform 1 0 45264 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_494
timestamp 1688980957
transform 1 0 46552 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_498
timestamp 1688980957
transform 1 0 46920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_502
timestamp 1688980957
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_519
timestamp 1688980957
transform 1 0 48852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_527
timestamp 1688980957
transform 1 0 49588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_553
timestamp 1688980957
transform 1 0 51980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_557
timestamp 1688980957
transform 1 0 52348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_569
timestamp 1688980957
transform 1 0 53452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_599
timestamp 1688980957
transform 1 0 56212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_611
timestamp 1688980957
transform 1 0 57316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_38
timestamp 1688980957
transform 1 0 4600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_44
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_58
timestamp 1688980957
transform 1 0 6440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_70
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1688980957
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_190
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_215
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_219
timestamp 1688980957
transform 1 0 21252 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_261
timestamp 1688980957
transform 1 0 25116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_278
timestamp 1688980957
transform 1 0 26680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_305
timestamp 1688980957
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_360
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_381
timestamp 1688980957
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_434
timestamp 1688980957
transform 1 0 41032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_474
timestamp 1688980957
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_477
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_496
timestamp 1688980957
transform 1 0 46736 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_507
timestamp 1688980957
transform 1 0 47748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_511
timestamp 1688980957
transform 1 0 48116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_519
timestamp 1688980957
transform 1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_533
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_564
timestamp 1688980957
transform 1 0 52992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_568
timestamp 1688980957
transform 1 0 53360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_578
timestamp 1688980957
transform 1 0 54280 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_586
timestamp 1688980957
transform 1 0 55016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_589
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_597
timestamp 1688980957
transform 1 0 56028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_602
timestamp 1688980957
transform 1 0 56488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_606
timestamp 1688980957
transform 1 0 56856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_615
timestamp 1688980957
transform 1 0 57684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_623
timestamp 1688980957
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_73
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_91
timestamp 1688980957
transform 1 0 9476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_129
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_140
timestamp 1688980957
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_144
timestamp 1688980957
transform 1 0 14352 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_156
timestamp 1688980957
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_244
timestamp 1688980957
transform 1 0 23552 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_248
timestamp 1688980957
transform 1 0 23920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_252
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_260
timestamp 1688980957
transform 1 0 25024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1688980957
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_319
timestamp 1688980957
transform 1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_362
timestamp 1688980957
transform 1 0 34408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_411
timestamp 1688980957
transform 1 0 38916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_415
timestamp 1688980957
transform 1 0 39284 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_441
timestamp 1688980957
transform 1 0 41676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_445
timestamp 1688980957
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_498
timestamp 1688980957
transform 1 0 46920 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_502
timestamp 1688980957
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_514
timestamp 1688980957
transform 1 0 48392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_518
timestamp 1688980957
transform 1 0 48760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_522
timestamp 1688980957
transform 1 0 49128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_526
timestamp 1688980957
transform 1 0 49496 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_531
timestamp 1688980957
transform 1 0 49956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_541
timestamp 1688980957
transform 1 0 50876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_595
timestamp 1688980957
transform 1 0 55844 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_612
timestamp 1688980957
transform 1 0 57408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_11
timestamp 1688980957
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1688980957
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_39
timestamp 1688980957
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_51
timestamp 1688980957
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_59
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_71
timestamp 1688980957
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_134
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_154
timestamp 1688980957
transform 1 0 15272 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_166
timestamp 1688980957
transform 1 0 16376 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_186
timestamp 1688980957
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1688980957
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_211
timestamp 1688980957
transform 1 0 20516 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_236
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1688980957
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_259
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_269
timestamp 1688980957
transform 1 0 25852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_281
timestamp 1688980957
transform 1 0 26956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_336
timestamp 1688980957
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_369
timestamp 1688980957
transform 1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_413
timestamp 1688980957
transform 1 0 39100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_417
timestamp 1688980957
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_469
timestamp 1688980957
transform 1 0 44252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_473
timestamp 1688980957
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_477
timestamp 1688980957
transform 1 0 44988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_488
timestamp 1688980957
transform 1 0 46000 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_492
timestamp 1688980957
transform 1 0 46368 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 1688980957
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_533
timestamp 1688980957
transform 1 0 50140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_541
timestamp 1688980957
transform 1 0 50876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_567
timestamp 1688980957
transform 1 0 53268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_571
timestamp 1688980957
transform 1 0 53636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_597
timestamp 1688980957
transform 1 0 56028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_623
timestamp 1688980957
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_11
timestamp 1688980957
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_28
timestamp 1688980957
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_32
timestamp 1688980957
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_73
timestamp 1688980957
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_94
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_104
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_138
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_142
timestamp 1688980957
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 1688980957
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_184
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_187
timestamp 1688980957
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_197
timestamp 1688980957
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_247
timestamp 1688980957
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_251
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_268
timestamp 1688980957
transform 1 0 25760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_295
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_299
timestamp 1688980957
transform 1 0 28612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_306
timestamp 1688980957
transform 1 0 29256 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_314
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_324
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_333
timestamp 1688980957
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_341
timestamp 1688980957
transform 1 0 32476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_345
timestamp 1688980957
transform 1 0 32844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_363
timestamp 1688980957
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_371
timestamp 1688980957
transform 1 0 35236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_417
timestamp 1688980957
transform 1 0 39468 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_425
timestamp 1688980957
transform 1 0 40204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_434
timestamp 1688980957
transform 1 0 41032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_439
timestamp 1688980957
transform 1 0 41492 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_457
timestamp 1688980957
transform 1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_465
timestamp 1688980957
transform 1 0 43884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_469
timestamp 1688980957
transform 1 0 44252 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_477
timestamp 1688980957
transform 1 0 44988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_494
timestamp 1688980957
transform 1 0 46552 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_502
timestamp 1688980957
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_529
timestamp 1688980957
transform 1 0 49772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_533
timestamp 1688980957
transform 1 0 50140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_537
timestamp 1688980957
transform 1 0 50508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_541
timestamp 1688980957
transform 1 0 50876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_545
timestamp 1688980957
transform 1 0 51244 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_551
timestamp 1688980957
transform 1 0 51796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_569
timestamp 1688980957
transform 1 0 53452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_588
timestamp 1688980957
transform 1 0 55200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_611
timestamp 1688980957
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1688980957
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_617
timestamp 1688980957
transform 1 0 57868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_621
timestamp 1688980957
transform 1 0 58236 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_57
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_66
timestamp 1688980957
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_78
timestamp 1688980957
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_96
timestamp 1688980957
transform 1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_162
timestamp 1688980957
transform 1 0 16008 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_170
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_178
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1688980957
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_213
timestamp 1688980957
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_218
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_238
timestamp 1688980957
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1688980957
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_285
timestamp 1688980957
transform 1 0 27324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_313
timestamp 1688980957
transform 1 0 29900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_323
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_327
timestamp 1688980957
transform 1 0 31188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_339
timestamp 1688980957
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_351
timestamp 1688980957
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_380
timestamp 1688980957
transform 1 0 36064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_388
timestamp 1688980957
transform 1 0 36800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_393
timestamp 1688980957
transform 1 0 37260 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_397
timestamp 1688980957
transform 1 0 37628 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_409
timestamp 1688980957
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_417
timestamp 1688980957
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_437
timestamp 1688980957
transform 1 0 41308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_464
timestamp 1688980957
transform 1 0 43792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_481
timestamp 1688980957
transform 1 0 45356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_485
timestamp 1688980957
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_489
timestamp 1688980957
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_493
timestamp 1688980957
transform 1 0 46460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_526
timestamp 1688980957
transform 1 0 49496 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_533
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_548
timestamp 1688980957
transform 1 0 51520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_556
timestamp 1688980957
transform 1 0 52256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_568
timestamp 1688980957
transform 1 0 53360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_585
timestamp 1688980957
transform 1 0 54924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_597
timestamp 1688980957
transform 1 0 56028 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_41
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_47
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_68
timestamp 1688980957
transform 1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_72
timestamp 1688980957
transform 1 0 7728 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_76
timestamp 1688980957
transform 1 0 8096 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_88
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_98
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1688980957
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_123
timestamp 1688980957
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_131
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_135
timestamp 1688980957
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1688980957
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_289
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_302
timestamp 1688980957
transform 1 0 28888 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_312
timestamp 1688980957
transform 1 0 29808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_333
timestamp 1688980957
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_341
timestamp 1688980957
transform 1 0 32476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_354
timestamp 1688980957
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_358
timestamp 1688980957
transform 1 0 34040 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_378
timestamp 1688980957
transform 1 0 35880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_387
timestamp 1688980957
transform 1 0 36708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_404
timestamp 1688980957
transform 1 0 38272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_408
timestamp 1688980957
transform 1 0 38640 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_436
timestamp 1688980957
transform 1 0 41216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_440
timestamp 1688980957
transform 1 0 41584 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_444
timestamp 1688980957
transform 1 0 41952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_453
timestamp 1688980957
transform 1 0 42780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_464
timestamp 1688980957
transform 1 0 43792 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_515
timestamp 1688980957
transform 1 0 48484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_527
timestamp 1688980957
transform 1 0 49588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_531
timestamp 1688980957
transform 1 0 49956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_550
timestamp 1688980957
transform 1 0 51704 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_558
timestamp 1688980957
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_573
timestamp 1688980957
transform 1 0 53820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_584
timestamp 1688980957
transform 1 0 54832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_588
timestamp 1688980957
transform 1 0 55200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_592
timestamp 1688980957
transform 1 0 55568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_612
timestamp 1688980957
transform 1 0 57408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_617
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_19
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_35
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_47
timestamp 1688980957
transform 1 0 5428 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_106
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_118
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_122
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_131
timestamp 1688980957
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_135
timestamp 1688980957
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_150
timestamp 1688980957
transform 1 0 14904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_154
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_168
timestamp 1688980957
transform 1 0 16560 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_192
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_231
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_248
timestamp 1688980957
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_326
timestamp 1688980957
transform 1 0 31096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_330
timestamp 1688980957
transform 1 0 31464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_358
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_362
timestamp 1688980957
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_381
timestamp 1688980957
transform 1 0 36156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_399
timestamp 1688980957
transform 1 0 37812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_416
timestamp 1688980957
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_473
timestamp 1688980957
transform 1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_511
timestamp 1688980957
transform 1 0 48116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_519
timestamp 1688980957
transform 1 0 48852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_529
timestamp 1688980957
transform 1 0 49772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_533
timestamp 1688980957
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_537
timestamp 1688980957
transform 1 0 50508 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_541
timestamp 1688980957
transform 1 0 50876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_553
timestamp 1688980957
transform 1 0 51980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_565
timestamp 1688980957
transform 1 0 53084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_577
timestamp 1688980957
transform 1 0 54188 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_585
timestamp 1688980957
transform 1 0 54924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_589
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_593
timestamp 1688980957
transform 1 0 55660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_598
timestamp 1688980957
transform 1 0 56120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_608
timestamp 1688980957
transform 1 0 57040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_612
timestamp 1688980957
transform 1 0 57408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_616
timestamp 1688980957
transform 1 0 57776 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_72
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_76
timestamp 1688980957
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_109
timestamp 1688980957
transform 1 0 11132 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_129
timestamp 1688980957
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_151
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_175
timestamp 1688980957
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_197
timestamp 1688980957
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_256
timestamp 1688980957
transform 1 0 24656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 1688980957
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_291
timestamp 1688980957
transform 1 0 27876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_295
timestamp 1688980957
transform 1 0 28244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_313
timestamp 1688980957
transform 1 0 29900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_389
timestamp 1688980957
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_453
timestamp 1688980957
transform 1 0 42780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_475
timestamp 1688980957
transform 1 0 44804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_479
timestamp 1688980957
transform 1 0 45172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_505
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_521
timestamp 1688980957
transform 1 0 49036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_557
timestamp 1688980957
transform 1 0 52348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_561
timestamp 1688980957
transform 1 0 52716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_581
timestamp 1688980957
transform 1 0 54556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_587
timestamp 1688980957
transform 1 0 55108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_614
timestamp 1688980957
transform 1 0 57592 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_38
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_42
timestamp 1688980957
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_46
timestamp 1688980957
transform 1 0 5336 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_110
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_174
timestamp 1688980957
transform 1 0 17112 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_184
timestamp 1688980957
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1688980957
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_239
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_248
timestamp 1688980957
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_261
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_283
timestamp 1688980957
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_295
timestamp 1688980957
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_299
timestamp 1688980957
transform 1 0 28612 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_318
timestamp 1688980957
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_337
timestamp 1688980957
transform 1 0 32108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_369
timestamp 1688980957
transform 1 0 35052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_406
timestamp 1688980957
transform 1 0 38456 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_410
timestamp 1688980957
transform 1 0 38824 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_414
timestamp 1688980957
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_473
timestamp 1688980957
transform 1 0 44620 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_486
timestamp 1688980957
transform 1 0 45816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_498
timestamp 1688980957
transform 1 0 46920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_528
timestamp 1688980957
transform 1 0 49680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_554
timestamp 1688980957
transform 1 0 52072 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_562
timestamp 1688980957
transform 1 0 52808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_581
timestamp 1688980957
transform 1 0 54556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_585
timestamp 1688980957
transform 1 0 54924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_619
timestamp 1688980957
transform 1 0 58052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_623
timestamp 1688980957
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_82
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_129
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_139
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_143
timestamp 1688980957
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_195
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_207
timestamp 1688980957
transform 1 0 20148 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_219
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_251
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_255
timestamp 1688980957
transform 1 0 24564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_267
timestamp 1688980957
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_299
timestamp 1688980957
transform 1 0 28612 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_308
timestamp 1688980957
transform 1 0 29440 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_341
timestamp 1688980957
transform 1 0 32476 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_355
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_367
timestamp 1688980957
transform 1 0 34868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_375
timestamp 1688980957
transform 1 0 35604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_380
timestamp 1688980957
transform 1 0 36064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_384
timestamp 1688980957
transform 1 0 36432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_389
timestamp 1688980957
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_401
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_413
timestamp 1688980957
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_425
timestamp 1688980957
transform 1 0 40204 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_437
timestamp 1688980957
transform 1 0 41308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_443
timestamp 1688980957
transform 1 0 41860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_471
timestamp 1688980957
transform 1 0 44436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_479
timestamp 1688980957
transform 1 0 45172 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_483
timestamp 1688980957
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_495
timestamp 1688980957
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 1688980957
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_529
timestamp 1688980957
transform 1 0 49772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_555
timestamp 1688980957
transform 1 0 52164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 1688980957
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_561
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_597
timestamp 1688980957
transform 1 0 56028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_51
timestamp 1688980957
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_73
timestamp 1688980957
transform 1 0 7820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_95
timestamp 1688980957
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_99
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_111
timestamp 1688980957
transform 1 0 11316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_117
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_126
timestamp 1688980957
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1688980957
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_160
timestamp 1688980957
transform 1 0 15824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_168
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_178
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_190
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_201
timestamp 1688980957
transform 1 0 19596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_213
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_225
timestamp 1688980957
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_269
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_295
timestamp 1688980957
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_299
timestamp 1688980957
transform 1 0 28612 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_332
timestamp 1688980957
transform 1 0 31648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_336
timestamp 1688980957
transform 1 0 32016 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_348
timestamp 1688980957
transform 1 0 33120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_360
timestamp 1688980957
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_397
timestamp 1688980957
transform 1 0 37628 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_433
timestamp 1688980957
transform 1 0 40940 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_441
timestamp 1688980957
transform 1 0 41676 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_445
timestamp 1688980957
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_466
timestamp 1688980957
transform 1 0 43976 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_470
timestamp 1688980957
transform 1 0 44344 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_474
timestamp 1688980957
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_489
timestamp 1688980957
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_501
timestamp 1688980957
transform 1 0 47196 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_505
timestamp 1688980957
transform 1 0 47564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_525
timestamp 1688980957
transform 1 0 49404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_530
timestamp 1688980957
transform 1 0 49864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_537
timestamp 1688980957
transform 1 0 50508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_566
timestamp 1688980957
transform 1 0 53176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_586
timestamp 1688980957
transform 1 0 55016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_597
timestamp 1688980957
transform 1 0 56028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_619
timestamp 1688980957
transform 1 0 58052 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_26
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_45
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_135
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_144
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_189
timestamp 1688980957
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_220
timestamp 1688980957
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_234
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_252
timestamp 1688980957
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_275
timestamp 1688980957
transform 1 0 26404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_330
timestamp 1688980957
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_343
timestamp 1688980957
transform 1 0 32660 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_346
timestamp 1688980957
transform 1 0 32936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_350
timestamp 1688980957
transform 1 0 33304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_367
timestamp 1688980957
transform 1 0 34868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_375
timestamp 1688980957
transform 1 0 35604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_409
timestamp 1688980957
transform 1 0 38732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_437
timestamp 1688980957
transform 1 0 41308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_458
timestamp 1688980957
transform 1 0 43240 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_482
timestamp 1688980957
transform 1 0 45448 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_494
timestamp 1688980957
transform 1 0 46552 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_502
timestamp 1688980957
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_513
timestamp 1688980957
transform 1 0 48300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_519
timestamp 1688980957
transform 1 0 48852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_544
timestamp 1688980957
transform 1 0 51152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_554
timestamp 1688980957
transform 1 0 52072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_558
timestamp 1688980957
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_561
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_569
timestamp 1688980957
transform 1 0 53452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_591
timestamp 1688980957
transform 1 0 55476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_610
timestamp 1688980957
transform 1 0 57224 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_19
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_46
timestamp 1688980957
transform 1 0 5336 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_54
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_64
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_72
timestamp 1688980957
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_98
timestamp 1688980957
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_102
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_116
timestamp 1688980957
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_137
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_170
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_176
timestamp 1688980957
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_257
timestamp 1688980957
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_274
timestamp 1688980957
transform 1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_293
timestamp 1688980957
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_360
timestamp 1688980957
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_398
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_437
timestamp 1688980957
transform 1 0 41308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_457
timestamp 1688980957
transform 1 0 43148 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_493
timestamp 1688980957
transform 1 0 46460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_501
timestamp 1688980957
transform 1 0 47196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_526
timestamp 1688980957
transform 1 0 49496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_530
timestamp 1688980957
transform 1 0 49864 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_555
timestamp 1688980957
transform 1 0 52164 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_567
timestamp 1688980957
transform 1 0 53268 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_584
timestamp 1688980957
transform 1 0 54832 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_597
timestamp 1688980957
transform 1 0 56028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_622
timestamp 1688980957
transform 1 0 58328 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_33
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_37
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_40
timestamp 1688980957
transform 1 0 4784 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_44
timestamp 1688980957
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_78
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_143
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_163
timestamp 1688980957
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_178
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_219
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_241
timestamp 1688980957
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_277
timestamp 1688980957
transform 1 0 26588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_290
timestamp 1688980957
transform 1 0 27784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_298
timestamp 1688980957
transform 1 0 28520 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_333
timestamp 1688980957
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_343
timestamp 1688980957
transform 1 0 32660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_353
timestamp 1688980957
transform 1 0 33580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_366
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_374
timestamp 1688980957
transform 1 0 35512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_387
timestamp 1688980957
transform 1 0 36708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_409
timestamp 1688980957
transform 1 0 38732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_413
timestamp 1688980957
transform 1 0 39100 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_442
timestamp 1688980957
transform 1 0 41768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_469
timestamp 1688980957
transform 1 0 44252 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_521
timestamp 1688980957
transform 1 0 49036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_525
timestamp 1688980957
transform 1 0 49404 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_556
timestamp 1688980957
transform 1 0 52256 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_561
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_581
timestamp 1688980957
transform 1 0 54556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_586
timestamp 1688980957
transform 1 0 55016 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 1688980957
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 1688980957
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_617
timestamp 1688980957
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_45
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_112
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_120
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_161
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_172
timestamp 1688980957
transform 1 0 16928 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_225
timestamp 1688980957
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_237
timestamp 1688980957
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_241
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_244
timestamp 1688980957
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_279
timestamp 1688980957
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_291
timestamp 1688980957
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_303
timestamp 1688980957
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_313
timestamp 1688980957
transform 1 0 29900 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_330
timestamp 1688980957
transform 1 0 31464 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_342
timestamp 1688980957
transform 1 0 32568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_346
timestamp 1688980957
transform 1 0 32936 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_402
timestamp 1688980957
transform 1 0 38088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_414
timestamp 1688980957
transform 1 0 39192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_473
timestamp 1688980957
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_485
timestamp 1688980957
transform 1 0 45724 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_497
timestamp 1688980957
transform 1 0 46828 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_505
timestamp 1688980957
transform 1 0 47564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_526
timestamp 1688980957
transform 1 0 49496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_530
timestamp 1688980957
transform 1 0 49864 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_566
timestamp 1688980957
transform 1 0 53176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_589
timestamp 1688980957
transform 1 0 55292 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_597
timestamp 1688980957
transform 1 0 56028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_616
timestamp 1688980957
transform 1 0 57776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_624
timestamp 1688980957
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_25
timestamp 1688980957
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_36
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_40
timestamp 1688980957
transform 1 0 4784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1688980957
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_74
timestamp 1688980957
transform 1 0 7912 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_139
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_159
timestamp 1688980957
transform 1 0 15732 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_210
timestamp 1688980957
transform 1 0 20424 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_266
timestamp 1688980957
transform 1 0 25576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_363
timestamp 1688980957
transform 1 0 34500 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_368
timestamp 1688980957
transform 1 0 34960 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_380
timestamp 1688980957
transform 1 0 36064 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_397
timestamp 1688980957
transform 1 0 37628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1688980957
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 1688980957
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 1688980957
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 1688980957
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_465
timestamp 1688980957
transform 1 0 43884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_475
timestamp 1688980957
transform 1 0 44804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_479
timestamp 1688980957
transform 1 0 45172 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_483
timestamp 1688980957
transform 1 0 45540 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_488
timestamp 1688980957
transform 1 0 46000 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_500
timestamp 1688980957
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_505
timestamp 1688980957
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_516
timestamp 1688980957
transform 1 0 48576 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_525
timestamp 1688980957
transform 1 0 49404 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_533
timestamp 1688980957
transform 1 0 50140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_561
timestamp 1688980957
transform 1 0 52716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_565
timestamp 1688980957
transform 1 0 53084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_569
timestamp 1688980957
transform 1 0 53452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_578
timestamp 1688980957
transform 1 0 54280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_590
timestamp 1688980957
transform 1 0 55384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_598
timestamp 1688980957
transform 1 0 56120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_612
timestamp 1688980957
transform 1 0 57408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_110
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_122
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_134
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_159
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_175
timestamp 1688980957
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_187
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_205
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_217
timestamp 1688980957
transform 1 0 21068 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_234
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_246
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_263
timestamp 1688980957
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_303
timestamp 1688980957
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_315
timestamp 1688980957
transform 1 0 30084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_327
timestamp 1688980957
transform 1 0 31188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_349
timestamp 1688980957
transform 1 0 33212 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_361
timestamp 1688980957
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_373
timestamp 1688980957
transform 1 0 35420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_381
timestamp 1688980957
transform 1 0 36156 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_414
timestamp 1688980957
transform 1 0 39192 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_425
timestamp 1688980957
transform 1 0 40204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_437
timestamp 1688980957
transform 1 0 41308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_449
timestamp 1688980957
transform 1 0 42412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1688980957
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_485
timestamp 1688980957
transform 1 0 45724 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_497
timestamp 1688980957
transform 1 0 46828 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_509
timestamp 1688980957
transform 1 0 47932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_521
timestamp 1688980957
transform 1 0 49036 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_529
timestamp 1688980957
transform 1 0 49772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_533
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_541
timestamp 1688980957
transform 1 0 50876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_560
timestamp 1688980957
transform 1 0 52624 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_582
timestamp 1688980957
transform 1 0 54648 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_601
timestamp 1688980957
transform 1 0 56396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_619
timestamp 1688980957
transform 1 0 58052 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_42
timestamp 1688980957
transform 1 0 4968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_46
timestamp 1688980957
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_52
timestamp 1688980957
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_74
timestamp 1688980957
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_78
timestamp 1688980957
transform 1 0 8280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_82
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_147
timestamp 1688980957
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_151
timestamp 1688980957
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_187
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_206
timestamp 1688980957
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_210
timestamp 1688980957
transform 1 0 20424 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_241
timestamp 1688980957
transform 1 0 23276 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_247
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_266
timestamp 1688980957
transform 1 0 25576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_297
timestamp 1688980957
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_324
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_386
timestamp 1688980957
transform 1 0 36616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_402
timestamp 1688980957
transform 1 0 38088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_406
timestamp 1688980957
transform 1 0 38456 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_434
timestamp 1688980957
transform 1 0 41032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_446
timestamp 1688980957
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_474
timestamp 1688980957
transform 1 0 44712 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_502
timestamp 1688980957
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_521
timestamp 1688980957
transform 1 0 49036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_529
timestamp 1688980957
transform 1 0 49772 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_542
timestamp 1688980957
transform 1 0 50968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_546
timestamp 1688980957
transform 1 0 51336 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_549
timestamp 1688980957
transform 1 0 51612 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_557
timestamp 1688980957
transform 1 0 52348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_595
timestamp 1688980957
transform 1 0 55844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 1688980957
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_37
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_55
timestamp 1688980957
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_72
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_76
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_91
timestamp 1688980957
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_101
timestamp 1688980957
transform 1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_158
timestamp 1688980957
transform 1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_166
timestamp 1688980957
transform 1 0 16376 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_183
timestamp 1688980957
transform 1 0 17940 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_206
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_248
timestamp 1688980957
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_303
timestamp 1688980957
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_325
timestamp 1688980957
transform 1 0 31004 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_342
timestamp 1688980957
transform 1 0 32568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_374
timestamp 1688980957
transform 1 0 35512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_378
timestamp 1688980957
transform 1 0 35880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_396
timestamp 1688980957
transform 1 0 37536 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1688980957
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_454
timestamp 1688980957
transform 1 0 42872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_526
timestamp 1688980957
transform 1 0 49496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_530
timestamp 1688980957
transform 1 0 49864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_558
timestamp 1688980957
transform 1 0 52440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 1688980957
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_589
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_618
timestamp 1688980957
transform 1 0 57960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_622
timestamp 1688980957
transform 1 0 58328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_20
timestamp 1688980957
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_32
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_48
timestamp 1688980957
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_80
timestamp 1688980957
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_84
timestamp 1688980957
transform 1 0 8832 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_106
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_145
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_188
timestamp 1688980957
transform 1 0 18400 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_213
timestamp 1688980957
transform 1 0 20700 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_235
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_239
timestamp 1688980957
transform 1 0 23092 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_277
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_298
timestamp 1688980957
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_306
timestamp 1688980957
transform 1 0 29256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_319
timestamp 1688980957
transform 1 0 30452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_354
timestamp 1688980957
transform 1 0 33672 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_387
timestamp 1688980957
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_435
timestamp 1688980957
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_466
timestamp 1688980957
transform 1 0 43976 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_496
timestamp 1688980957
transform 1 0 46736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_505
timestamp 1688980957
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_524
timestamp 1688980957
transform 1 0 49312 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_536
timestamp 1688980957
transform 1 0 50416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_569
timestamp 1688980957
transform 1 0 53452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_579
timestamp 1688980957
transform 1 0 54372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_613
timestamp 1688980957
transform 1 0 57500 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_89
timestamp 1688980957
transform 1 0 9292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_125
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_176
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_188
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_206
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_218
timestamp 1688980957
transform 1 0 21160 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_226
timestamp 1688980957
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_246
timestamp 1688980957
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_279
timestamp 1688980957
transform 1 0 26772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_303
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_319
timestamp 1688980957
transform 1 0 30452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_331
timestamp 1688980957
transform 1 0 31556 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_337
timestamp 1688980957
transform 1 0 32108 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_349
timestamp 1688980957
transform 1 0 33212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_361
timestamp 1688980957
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_369
timestamp 1688980957
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_406
timestamp 1688980957
transform 1 0 38456 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_410
timestamp 1688980957
transform 1 0 38824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_472
timestamp 1688980957
transform 1 0 44528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_481
timestamp 1688980957
transform 1 0 45356 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_485
timestamp 1688980957
transform 1 0 45724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_497
timestamp 1688980957
transform 1 0 46828 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_509
timestamp 1688980957
transform 1 0 47932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_521
timestamp 1688980957
transform 1 0 49036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_529
timestamp 1688980957
transform 1 0 49772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_533
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_537
timestamp 1688980957
transform 1 0 50508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_557
timestamp 1688980957
transform 1 0 52348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_565
timestamp 1688980957
transform 1 0 53084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_576
timestamp 1688980957
transform 1 0 54096 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_585
timestamp 1688980957
transform 1 0 54924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_589
timestamp 1688980957
transform 1 0 55292 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_595
timestamp 1688980957
transform 1 0 55844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_623
timestamp 1688980957
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_31
timestamp 1688980957
transform 1 0 3956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_86
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_202
timestamp 1688980957
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_214
timestamp 1688980957
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_264
timestamp 1688980957
transform 1 0 25392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_276
timestamp 1688980957
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_314
timestamp 1688980957
transform 1 0 29992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_326
timestamp 1688980957
transform 1 0 31096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_330
timestamp 1688980957
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_341
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_353
timestamp 1688980957
transform 1 0 33580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_365
timestamp 1688980957
transform 1 0 34684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_369
timestamp 1688980957
transform 1 0 35052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_372
timestamp 1688980957
transform 1 0 35328 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_376
timestamp 1688980957
transform 1 0 35696 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_388
timestamp 1688980957
transform 1 0 36800 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_397
timestamp 1688980957
transform 1 0 37628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_409
timestamp 1688980957
transform 1 0 38732 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_421
timestamp 1688980957
transform 1 0 39836 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_433
timestamp 1688980957
transform 1 0 40940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 1688980957
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_459
timestamp 1688980957
transform 1 0 43332 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_471
timestamp 1688980957
transform 1 0 44436 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_483
timestamp 1688980957
transform 1 0 45540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_491
timestamp 1688980957
transform 1 0 46276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_500
timestamp 1688980957
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_513
timestamp 1688980957
transform 1 0 48300 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_530
timestamp 1688980957
transform 1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_558
timestamp 1688980957
transform 1 0 52440 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_573
timestamp 1688980957
transform 1 0 53820 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_581
timestamp 1688980957
transform 1 0 54556 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 1688980957
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_597
timestamp 1688980957
transform 1 0 56028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_610
timestamp 1688980957
transform 1 0 57224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_614
timestamp 1688980957
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_66
timestamp 1688980957
transform 1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_94
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_98
timestamp 1688980957
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_145
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_150
timestamp 1688980957
transform 1 0 14904 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_156
timestamp 1688980957
transform 1 0 15456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_159
timestamp 1688980957
transform 1 0 15732 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_185
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_239
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_261
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_328
timestamp 1688980957
transform 1 0 31280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_338
timestamp 1688980957
transform 1 0 32200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_347
timestamp 1688980957
transform 1 0 33028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_356
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_360
timestamp 1688980957
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_382
timestamp 1688980957
transform 1 0 36248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_417
timestamp 1688980957
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_464
timestamp 1688980957
transform 1 0 43792 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 1688980957
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_489
timestamp 1688980957
transform 1 0 46092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_502
timestamp 1688980957
transform 1 0 47288 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_516
timestamp 1688980957
transform 1 0 48576 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_528
timestamp 1688980957
transform 1 0 49680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_549
timestamp 1688980957
transform 1 0 51612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_558
timestamp 1688980957
transform 1 0 52440 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_562
timestamp 1688980957
transform 1 0 52808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_574
timestamp 1688980957
transform 1 0 53912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_582
timestamp 1688980957
transform 1 0 54648 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 1688980957
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_589
timestamp 1688980957
transform 1 0 55292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_593
timestamp 1688980957
transform 1 0 55660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_620
timestamp 1688980957
transform 1 0 58144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_624
timestamp 1688980957
transform 1 0 58512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_43
timestamp 1688980957
transform 1 0 5060 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_61
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_73
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_92
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_208
timestamp 1688980957
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_212
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_241
timestamp 1688980957
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_276
timestamp 1688980957
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_285
timestamp 1688980957
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_289
timestamp 1688980957
transform 1 0 27692 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_389
timestamp 1688980957
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_409
timestamp 1688980957
transform 1 0 38732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_426
timestamp 1688980957
transform 1 0 40296 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_474
timestamp 1688980957
transform 1 0 44712 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_478
timestamp 1688980957
transform 1 0 45080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_482
timestamp 1688980957
transform 1 0 45448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_503
timestamp 1688980957
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_526
timestamp 1688980957
transform 1 0 49496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_530
timestamp 1688980957
transform 1 0 49864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_534
timestamp 1688980957
transform 1 0 50232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_537
timestamp 1688980957
transform 1 0 50508 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_570
timestamp 1688980957
transform 1 0 53544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_595
timestamp 1688980957
transform 1 0 55844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 1688980957
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_45
timestamp 1688980957
transform 1 0 5244 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_50
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_62
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_74
timestamp 1688980957
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_89
timestamp 1688980957
transform 1 0 9292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_101
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 1688980957
transform 1 0 11500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_122
timestamp 1688980957
transform 1 0 12328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_126
timestamp 1688980957
transform 1 0 12696 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_185
timestamp 1688980957
transform 1 0 18124 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_208
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_313
timestamp 1688980957
transform 1 0 29900 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_360
timestamp 1688980957
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_381
timestamp 1688980957
transform 1 0 36156 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_430
timestamp 1688980957
transform 1 0 40664 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_434
timestamp 1688980957
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_473
timestamp 1688980957
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_477
timestamp 1688980957
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_481
timestamp 1688980957
transform 1 0 45356 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_498
timestamp 1688980957
transform 1 0 46920 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_516
timestamp 1688980957
transform 1 0 48576 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_528
timestamp 1688980957
transform 1 0 49680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_565
timestamp 1688980957
transform 1 0 53084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_585
timestamp 1688980957
transform 1 0 54924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_619
timestamp 1688980957
transform 1 0 58052 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_623
timestamp 1688980957
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_61
timestamp 1688980957
transform 1 0 6716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_73
timestamp 1688980957
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_79
timestamp 1688980957
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_91
timestamp 1688980957
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_103
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_142
timestamp 1688980957
transform 1 0 14168 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_146
timestamp 1688980957
transform 1 0 14536 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_179
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_187
timestamp 1688980957
transform 1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_242
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_262
timestamp 1688980957
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_289
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_299
timestamp 1688980957
transform 1 0 28612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_319
timestamp 1688980957
transform 1 0 30452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_333
timestamp 1688980957
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_353
timestamp 1688980957
transform 1 0 33580 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_357
timestamp 1688980957
transform 1 0 33948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_384
timestamp 1688980957
transform 1 0 36432 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_388
timestamp 1688980957
transform 1 0 36800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_402
timestamp 1688980957
transform 1 0 38088 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_486
timestamp 1688980957
transform 1 0 45816 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_497
timestamp 1688980957
transform 1 0 46828 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_501
timestamp 1688980957
transform 1 0 47196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_522
timestamp 1688980957
transform 1 0 49128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_532
timestamp 1688980957
transform 1 0 50048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_545
timestamp 1688980957
transform 1 0 51244 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_557
timestamp 1688980957
transform 1 0 52348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_561
timestamp 1688980957
transform 1 0 52716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_571
timestamp 1688980957
transform 1 0 53636 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_599
timestamp 1688980957
transform 1 0 56212 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_169
timestamp 1688980957
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_181
timestamp 1688980957
transform 1 0 17756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1688980957
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_223
timestamp 1688980957
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_227
timestamp 1688980957
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_236
timestamp 1688980957
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_290
timestamp 1688980957
transform 1 0 27784 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_302
timestamp 1688980957
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_381
timestamp 1688980957
transform 1 0 36156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_406
timestamp 1688980957
transform 1 0 38456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_437
timestamp 1688980957
transform 1 0 41308 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_465
timestamp 1688980957
transform 1 0 43884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_474
timestamp 1688980957
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_477
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_485
timestamp 1688980957
transform 1 0 45724 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_503
timestamp 1688980957
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_512
timestamp 1688980957
transform 1 0 48208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_524
timestamp 1688980957
transform 1 0 49312 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_544
timestamp 1688980957
transform 1 0 51152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_569
timestamp 1688980957
transform 1 0 53452 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_585
timestamp 1688980957
transform 1 0 54924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_597
timestamp 1688980957
transform 1 0 56028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_619
timestamp 1688980957
transform 1 0 58052 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_86
timestamp 1688980957
transform 1 0 9016 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_90
timestamp 1688980957
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_94
timestamp 1688980957
transform 1 0 9752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_153
timestamp 1688980957
transform 1 0 15180 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_157
timestamp 1688980957
transform 1 0 15548 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_177
timestamp 1688980957
transform 1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_185
timestamp 1688980957
transform 1 0 18124 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_194
timestamp 1688980957
transform 1 0 18952 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_208
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_245
timestamp 1688980957
transform 1 0 23644 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_258
timestamp 1688980957
transform 1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_289
timestamp 1688980957
transform 1 0 27692 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_313
timestamp 1688980957
transform 1 0 29900 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_325
timestamp 1688980957
transform 1 0 31004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1688980957
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 1688980957
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_441
timestamp 1688980957
transform 1 0 41676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_445
timestamp 1688980957
transform 1 0 42044 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_475
timestamp 1688980957
transform 1 0 44804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_495
timestamp 1688980957
transform 1 0 46644 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_499
timestamp 1688980957
transform 1 0 47012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 1688980957
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_509
timestamp 1688980957
transform 1 0 47932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_521
timestamp 1688980957
transform 1 0 49036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_533
timestamp 1688980957
transform 1 0 50140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_536
timestamp 1688980957
transform 1 0 50416 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_561
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_567
timestamp 1688980957
transform 1 0 53268 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_579
timestamp 1688980957
transform 1 0 54372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_591
timestamp 1688980957
transform 1 0 55476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_603
timestamp 1688980957
transform 1 0 56580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 1688980957
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_49
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_73
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_120
timestamp 1688980957
transform 1 0 12144 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_205
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_217
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_229
timestamp 1688980957
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_241
timestamp 1688980957
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_249
timestamp 1688980957
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_259
timestamp 1688980957
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_262
timestamp 1688980957
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_274
timestamp 1688980957
transform 1 0 26312 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_282
timestamp 1688980957
transform 1 0 27048 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_286
timestamp 1688980957
transform 1 0 27416 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_315
timestamp 1688980957
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_340
timestamp 1688980957
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_352
timestamp 1688980957
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_473
timestamp 1688980957
transform 1 0 44620 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_486
timestamp 1688980957
transform 1 0 45816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_510
timestamp 1688980957
transform 1 0 48024 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_514
timestamp 1688980957
transform 1 0 48392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_518
timestamp 1688980957
transform 1 0 48760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_544
timestamp 1688980957
transform 1 0 51152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_584
timestamp 1688980957
transform 1 0 54832 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1688980957
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1688980957
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_82
timestamp 1688980957
transform 1 0 8648 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_86
timestamp 1688980957
transform 1 0 9016 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_98
timestamp 1688980957
transform 1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_117
timestamp 1688980957
transform 1 0 11868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_121
timestamp 1688980957
transform 1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_129
timestamp 1688980957
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_140
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_208
timestamp 1688980957
transform 1 0 20240 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_303
timestamp 1688980957
transform 1 0 28980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_345
timestamp 1688980957
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_357
timestamp 1688980957
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_369
timestamp 1688980957
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_381
timestamp 1688980957
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 1688980957
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_467
timestamp 1688980957
transform 1 0 44068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_502
timestamp 1688980957
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_521
timestamp 1688980957
transform 1 0 49036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_554
timestamp 1688980957
transform 1 0 52072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_558
timestamp 1688980957
transform 1 0 52440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_586
timestamp 1688980957
transform 1 0 55016 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_590
timestamp 1688980957
transform 1 0 55384 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_602
timestamp 1688980957
transform 1 0 56488 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_614
timestamp 1688980957
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_617
timestamp 1688980957
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_171
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_175
timestamp 1688980957
transform 1 0 17204 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_192
timestamp 1688980957
transform 1 0 18768 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_205
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_217
timestamp 1688980957
transform 1 0 21068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_229
timestamp 1688980957
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_241
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_249
timestamp 1688980957
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_336
timestamp 1688980957
transform 1 0 32016 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_340
timestamp 1688980957
transform 1 0 32384 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_352
timestamp 1688980957
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_473
timestamp 1688980957
transform 1 0 44620 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_526
timestamp 1688980957
transform 1 0 49496 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_549
timestamp 1688980957
transform 1 0 51612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_553
timestamp 1688980957
transform 1 0 51980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 1688980957
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1688980957
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1688980957
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_187
timestamp 1688980957
transform 1 0 18308 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_198
timestamp 1688980957
transform 1 0 19320 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_210
timestamp 1688980957
transform 1 0 20424 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_222
timestamp 1688980957
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_289
timestamp 1688980957
transform 1 0 27692 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_298
timestamp 1688980957
transform 1 0 28520 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_307
timestamp 1688980957
transform 1 0 29348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_315
timestamp 1688980957
transform 1 0 30084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_324
timestamp 1688980957
transform 1 0 30912 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_328
timestamp 1688980957
transform 1 0 31280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_332
timestamp 1688980957
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_473
timestamp 1688980957
transform 1 0 44620 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_513
timestamp 1688980957
transform 1 0 48300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_525
timestamp 1688980957
transform 1 0 49404 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_533
timestamp 1688980957
transform 1 0 50140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_558
timestamp 1688980957
transform 1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_573
timestamp 1688980957
transform 1 0 53820 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_584
timestamp 1688980957
transform 1 0 54832 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_596
timestamp 1688980957
transform 1 0 55936 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_608
timestamp 1688980957
transform 1 0 57040 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 1688980957
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1688980957
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 1688980957
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_293
timestamp 1688980957
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_337
timestamp 1688980957
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_349
timestamp 1688980957
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_393
timestamp 1688980957
transform 1 0 37260 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_405
timestamp 1688980957
transform 1 0 38364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_417
timestamp 1688980957
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_449
timestamp 1688980957
transform 1 0 42412 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_461
timestamp 1688980957
transform 1 0 43516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_473
timestamp 1688980957
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1688980957
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_501
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_505
timestamp 1688980957
transform 1 0 47564 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_517
timestamp 1688980957
transform 1 0 48668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_529
timestamp 1688980957
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1688980957
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_545
timestamp 1688980957
transform 1 0 51244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_557
timestamp 1688980957
transform 1 0 52348 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_561
timestamp 1688980957
transform 1 0 52716 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_573
timestamp 1688980957
transform 1 0 53820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_585
timestamp 1688980957
transform 1 0 54924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1688980957
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_613
timestamp 1688980957
transform 1 0 57500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_617
timestamp 1688980957
transform 1 0 57868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 6072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 43148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold6 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 40940 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 44068 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 44252 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 41308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 41032 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold13
timestamp 1688980957
transform -1 0 39100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 37996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 26404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold18
timestamp 1688980957
transform -1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 25116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 21344 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 39744 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 39284 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold25
timestamp 1688980957
transform -1 0 36156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 33764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 20608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 31740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 30176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 35972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 35972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 44712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 44620 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 29808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold36
timestamp 1688980957
transform -1 0 28980 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 24564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 23644 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 33028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 34500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 45724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold45
timestamp 1688980957
transform 1 0 46276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 46552 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold48
timestamp 1688980957
transform -1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 15272 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 48484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 49956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 26312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 45816 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 45816 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 17664 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 17480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 15456 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 54188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold65
timestamp 1688980957
transform -1 0 53544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 51612 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 49312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 50140 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold70
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 45540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold73
timestamp 1688980957
transform -1 0 44896 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 29808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 49496 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 49772 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 7912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 9936 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 52624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 52624 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold88
timestamp 1688980957
transform -1 0 25208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 27324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 58604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold91
timestamp 1688980957
transform -1 0 57776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 55384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 13984 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 13524 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 13984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 43700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 43056 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 55292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 54280 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 43516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 41860 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold104
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 21620 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 53452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold107
timestamp 1688980957
transform -1 0 51980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 51152 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 50968 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 50600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 53544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 56028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 55476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold114
timestamp 1688980957
transform -1 0 57040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 55844 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 55108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 56028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 44068 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 43976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 54280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 53452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 55016 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 53452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 52348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 47380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 48116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 34592 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold129
timestamp 1688980957
transform -1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 30820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 17204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 16192 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold134
timestamp 1688980957
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 10764 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold137
timestamp 1688980957
transform -1 0 16560 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 14720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 48116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 49864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform -1 0 7176 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 49036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 49036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform -1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 43148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 54832 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 58604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 58420 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 42044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold156
timestamp 1688980957
transform -1 0 38732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform -1 0 36892 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform 1 0 55108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform -1 0 54924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform 1 0 40848 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 40572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 9844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform -1 0 14996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform -1 0 38272 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 38456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 27140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 58604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform 1 0 55660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 17112 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 16284 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform -1 0 8648 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 6256 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 55476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 55476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 29348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 32108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 29440 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 13524 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform -1 0 13616 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 58604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 58328 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 58604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 58052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform 1 0 12788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 12696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 34316 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform 1 0 33028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 35972 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 35880 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold197
timestamp 1688980957
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold200 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform -1 0 13708 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 41308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 58604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 16560 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform -1 0 11408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 20792 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 19780 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 58604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 57316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 54740 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 56028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 54464 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 54280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform 1 0 14260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 13984 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 16560 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 16284 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 44804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform 1 0 11408 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 11132 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 49036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 49404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 15548 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 47472 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 46736 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 23552 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 22816 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform 1 0 11592 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 11408 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 51428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 53176 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 49312 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 48576 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform 1 0 50508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 50048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform 1 0 42964 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 42320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform -1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 18952 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 16560 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform -1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold259
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform -1 0 53176 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 52624 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform -1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform 1 0 19136 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform -1 0 48576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform -1 0 51888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform -1 0 52624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform 1 0 45540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform -1 0 44804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 4140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform -1 0 20148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold276
timestamp 1688980957
transform -1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform -1 0 9568 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform 1 0 46460 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 46092 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 26772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform -1 0 26036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 7912 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 7176 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 18032 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform 1 0 18308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform -1 0 18308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform -1 0 20516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform -1 0 6256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform 1 0 36340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform 1 0 37168 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform 1 0 41216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform -1 0 41216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 21804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform -1 0 21068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform 1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 19044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform 1 0 6440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform -1 0 6072 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform -1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 43884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform -1 0 43976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform -1 0 24104 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 3680 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 48300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold313
timestamp 1688980957
transform 1 0 46920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform -1 0 47196 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 45724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform -1 0 44804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform -1 0 40572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform -1 0 42044 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform -1 0 23920 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform 1 0 43240 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 42320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold326
timestamp 1688980957
transform -1 0 58604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 58604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform 1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform -1 0 35972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform -1 0 23092 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold335
timestamp 1688980957
transform -1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform -1 0 10948 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform -1 0 39284 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform -1 0 40020 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform -1 0 8464 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform -1 0 44528 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform -1 0 43792 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 24656 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform -1 0 24012 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform 1 0 54188 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform -1 0 54096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform -1 0 34684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform -1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 41768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform -1 0 41308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform -1 0 28520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform -1 0 28244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform -1 0 5244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform -1 0 7912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 1688980957
transform 1 0 48944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform -1 0 49496 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform -1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform 1 0 35236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold362
timestamp 1688980957
transform -1 0 35236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform -1 0 24012 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform -1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform 1 0 4048 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform -1 0 34500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform -1 0 36616 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform -1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform -1 0 14628 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 1688980957
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 1688980957
transform -1 0 16928 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform 1 0 33028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 1688980957
transform -1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform 1 0 37996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform -1 0 37996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform 1 0 30544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold383
timestamp 1688980957
transform -1 0 32016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform -1 0 31556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform -1 0 30820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 1688980957
transform -1 0 58604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform -1 0 58052 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform 1 0 55108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform -1 0 55108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform 1 0 2116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 1688980957
transform 1 0 2208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 1688980957
transform 1 0 33120 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold393
timestamp 1688980957
transform -1 0 33028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold394
timestamp 1688980957
transform -1 0 36248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold395
timestamp 1688980957
transform -1 0 36892 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 1688980957
transform -1 0 4968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 1688980957
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 1688980957
transform 1 0 50508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold399
timestamp 1688980957
transform -1 0 52256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 1688980957
transform -1 0 51704 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold401
timestamp 1688980957
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold402
timestamp 1688980957
transform -1 0 49956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 1688980957
transform -1 0 49312 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold404
timestamp 1688980957
transform -1 0 6992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 1688980957
transform -1 0 7728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold406
timestamp 1688980957
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold407
timestamp 1688980957
transform -1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 1688980957
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold409
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 1688980957
transform 1 0 38916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold411
timestamp 1688980957
transform -1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 1688980957
transform -1 0 36156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 1688980957
transform 1 0 37444 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 1688980957
transform -1 0 37444 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 1688980957
transform -1 0 36708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 1688980957
transform -1 0 35972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold417
timestamp 1688980957
transform -1 0 28060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 1688980957
transform -1 0 29532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 1688980957
transform -1 0 52348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 1688980957
transform -1 0 53452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 1688980957
transform -1 0 32016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 1688980957
transform -1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 1688980957
transform 1 0 7544 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 1688980957
transform -1 0 6992 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 1688980957
transform -1 0 31740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 1688980957
transform -1 0 31648 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 1688980957
transform -1 0 33948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 1688980957
transform -1 0 35420 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 1688980957
transform -1 0 39468 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold432
timestamp 1688980957
transform -1 0 38732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 1688980957
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 1688980957
transform -1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 1688980957
transform 1 0 40388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 1688980957
transform -1 0 40940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 1688980957
transform 1 0 37720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 1688980957
transform -1 0 37720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 1688980957
transform -1 0 48300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 1688980957
transform 1 0 46644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 1688980957
transform 1 0 26956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 1688980957
transform -1 0 26312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 1688980957
transform 1 0 37720 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 1688980957
transform -1 0 37720 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 1688980957
transform 1 0 28796 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 1688980957
transform 1 0 28704 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 1688980957
transform -1 0 58604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 1688980957
transform -1 0 58052 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 1688980957
transform -1 0 3588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 1688980957
transform 1 0 38456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 1688980957
transform -1 0 38456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 1688980957
transform -1 0 51980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 1688980957
transform -1 0 51152 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 1688980957
transform 1 0 45172 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 1688980957
transform -1 0 46644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold457
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 1688980957
transform 1 0 25024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 1688980957
transform 1 0 55292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 1688980957
transform -1 0 54556 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 1688980957
transform -1 0 44804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 1688980957
transform -1 0 44068 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 1688980957
transform -1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 1688980957
transform -1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 1688980957
transform -1 0 49404 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 1688980957
transform -1 0 49496 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 1688980957
transform 1 0 30728 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 1688980957
transform -1 0 30728 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 1688980957
transform -1 0 28428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold470
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 1688980957
transform -1 0 25300 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 1688980957
transform 1 0 54372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 1688980957
transform -1 0 54832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 1688980957
transform 1 0 18584 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 1688980957
transform -1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 1688980957
transform -1 0 23000 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 1688980957
transform 1 0 16928 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 1688980957
transform -1 0 18400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 1688980957
transform -1 0 20884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 1688980957
transform -1 0 23092 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 1688980957
transform 1 0 50968 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 1688980957
transform -1 0 50968 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 1688980957
transform -1 0 46644 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 1688980957
transform 1 0 45172 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 1688980957
transform 1 0 24104 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 1688980957
transform -1 0 24104 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 1688980957
transform -1 0 58604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 1688980957
transform -1 0 57316 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 1688980957
transform 1 0 27048 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 1688980957
transform -1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 1688980957
transform -1 0 28980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold493
timestamp 1688980957
transform -1 0 28060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 1688980957
transform -1 0 52716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 1688980957
transform -1 0 53452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold496
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold497
timestamp 1688980957
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold498
timestamp 1688980957
transform -1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 1688980957
transform 1 0 55108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 1688980957
transform -1 0 56212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold501
timestamp 1688980957
transform -1 0 54832 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold502
timestamp 1688980957
transform -1 0 54372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold503
timestamp 1688980957
transform 1 0 43976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 1688980957
transform -1 0 45816 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 1688980957
transform 1 0 42596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold506
timestamp 1688980957
transform -1 0 42412 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold507
timestamp 1688980957
transform 1 0 51612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold508
timestamp 1688980957
transform -1 0 52440 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 1688980957
transform -1 0 26312 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 1688980957
transform -1 0 27692 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold511
timestamp 1688980957
transform -1 0 25208 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold512
timestamp 1688980957
transform -1 0 25116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold513
timestamp 1688980957
transform 1 0 25300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 1688980957
transform -1 0 25300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold516
timestamp 1688980957
transform -1 0 28520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold517
timestamp 1688980957
transform 1 0 48392 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold518
timestamp 1688980957
transform -1 0 48208 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 1688980957
transform -1 0 47104 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold521
timestamp 1688980957
transform 1 0 29256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 1688980957
transform -1 0 28980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 1688980957
transform 1 0 19320 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 1688980957
transform 1 0 18952 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 1688980957
transform -1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 1688980957
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold527
timestamp 1688980957
transform -1 0 32016 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold528
timestamp 1688980957
transform -1 0 30912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold529
timestamp 1688980957
transform 1 0 31464 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 1688980957
transform -1 0 31740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 1688980957
transform 1 0 43056 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 1688980957
transform -1 0 42228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 1688980957
transform -1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 1688980957
transform 1 0 29716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 1688980957
transform -1 0 23736 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 1688980957
transform -1 0 23920 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 1688980957
transform -1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 1688980957
transform 1 0 46644 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 1688980957
transform -1 0 46644 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 1688980957
transform -1 0 22816 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 1688980957
transform -1 0 32384 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 1688980957
transform -1 0 32844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 1688980957
transform -1 0 42228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 1688980957
transform -1 0 40572 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 1688980957
transform -1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold548
timestamp 1688980957
transform -1 0 41308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 1688980957
transform -1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold550
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold551
timestamp 1688980957
transform 1 0 16928 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 1688980957
transform -1 0 13340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 1688980957
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold554
timestamp 1688980957
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold555
timestamp 1688980957
transform -1 0 44620 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 1688980957
transform -1 0 44068 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 1688980957
transform -1 0 45172 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold558 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold561
timestamp 1688980957
transform -1 0 17112 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 1688980957
transform -1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold563
timestamp 1688980957
transform -1 0 11408 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold565
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold566
timestamp 1688980957
transform -1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold567
timestamp 1688980957
transform -1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold568
timestamp 1688980957
transform -1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold569 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold570
timestamp 1688980957
transform -1 0 16468 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold571
timestamp 1688980957
transform 1 0 38640 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold572
timestamp 1688980957
transform -1 0 39560 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold573
timestamp 1688980957
transform -1 0 50508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold574
timestamp 1688980957
transform -1 0 49956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold575
timestamp 1688980957
transform 1 0 34500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold576
timestamp 1688980957
transform -1 0 35512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold577
timestamp 1688980957
transform -1 0 58604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold578
timestamp 1688980957
transform -1 0 58604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold579
timestamp 1688980957
transform -1 0 58604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold580
timestamp 1688980957
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold581
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold582
timestamp 1688980957
transform -1 0 40664 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold583
timestamp 1688980957
transform -1 0 51244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 1688980957
transform -1 0 50876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold585
timestamp 1688980957
transform 1 0 42320 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold586
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold587
timestamp 1688980957
transform -1 0 24288 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold588
timestamp 1688980957
transform -1 0 22540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold589
timestamp 1688980957
transform -1 0 47288 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold590
timestamp 1688980957
transform -1 0 48300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold591
timestamp 1688980957
transform -1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold592
timestamp 1688980957
transform -1 0 46736 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold593
timestamp 1688980957
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold594
timestamp 1688980957
transform 1 0 29716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold595
timestamp 1688980957
transform -1 0 39100 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold596
timestamp 1688980957
transform -1 0 37996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold597
timestamp 1688980957
transform -1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold598
timestamp 1688980957
transform -1 0 27692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold599
timestamp 1688980957
transform -1 0 54280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold600
timestamp 1688980957
transform 1 0 53636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold601
timestamp 1688980957
transform -1 0 57040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold602
timestamp 1688980957
transform -1 0 56304 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold603
timestamp 1688980957
transform 1 0 43424 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold604
timestamp 1688980957
transform -1 0 44804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold605
timestamp 1688980957
transform -1 0 52440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold606
timestamp 1688980957
transform 1 0 51612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold607
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold608
timestamp 1688980957
transform 1 0 20332 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold609
timestamp 1688980957
transform -1 0 25576 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold610
timestamp 1688980957
transform -1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold611
timestamp 1688980957
transform -1 0 19596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold612
timestamp 1688980957
transform -1 0 19412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold613
timestamp 1688980957
transform -1 0 24104 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold614
timestamp 1688980957
transform -1 0 23920 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold615
timestamp 1688980957
transform -1 0 29256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold616
timestamp 1688980957
transform -1 0 29532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold617
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold618
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold619
timestamp 1688980957
transform 1 0 33580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold620
timestamp 1688980957
transform -1 0 32936 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold621
timestamp 1688980957
transform 1 0 2208 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold622
timestamp 1688980957
transform -1 0 3680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold623
timestamp 1688980957
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold624
timestamp 1688980957
transform -1 0 30268 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold625
timestamp 1688980957
transform -1 0 28980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold626
timestamp 1688980957
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold627
timestamp 1688980957
transform -1 0 18952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold628
timestamp 1688980957
transform -1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold629
timestamp 1688980957
transform 1 0 37812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold630
timestamp 1688980957
transform -1 0 39008 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold631
timestamp 1688980957
transform -1 0 38916 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold632
timestamp 1688980957
transform 1 0 4140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold633
timestamp 1688980957
transform -1 0 3680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold634
timestamp 1688980957
transform -1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold635
timestamp 1688980957
transform -1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold636
timestamp 1688980957
transform 1 0 33764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold637
timestamp 1688980957
transform -1 0 34592 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold638
timestamp 1688980957
transform -1 0 34592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold639
timestamp 1688980957
transform 1 0 47012 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold640
timestamp 1688980957
transform -1 0 47840 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold641
timestamp 1688980957
transform -1 0 46276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold642
timestamp 1688980957
transform -1 0 53360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold643
timestamp 1688980957
transform -1 0 54096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold644
timestamp 1688980957
transform -1 0 53360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold645
timestamp 1688980957
transform -1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold646
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold647
timestamp 1688980957
transform -1 0 42320 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold648
timestamp 1688980957
transform 1 0 22080 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold649
timestamp 1688980957
transform -1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold650
timestamp 1688980957
transform -1 0 23000 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold651
timestamp 1688980957
transform -1 0 58604 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold652
timestamp 1688980957
transform -1 0 57684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold653
timestamp 1688980957
transform -1 0 57776 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold654
timestamp 1688980957
transform -1 0 58604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold655
timestamp 1688980957
transform -1 0 56304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold656
timestamp 1688980957
transform 1 0 55476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold657
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold658
timestamp 1688980957
transform -1 0 11224 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold659
timestamp 1688980957
transform -1 0 9844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  hold660
timestamp 1688980957
transform 1 0 15088 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold661
timestamp 1688980957
transform -1 0 21252 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold662
timestamp 1688980957
transform -1 0 20516 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold663
timestamp 1688980957
transform -1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold664
timestamp 1688980957
transform -1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold665
timestamp 1688980957
transform -1 0 8280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold666
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold667
timestamp 1688980957
transform 1 0 50876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold668
timestamp 1688980957
transform -1 0 52348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold669
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold670
timestamp 1688980957
transform -1 0 15824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold671
timestamp 1688980957
transform -1 0 31372 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold672
timestamp 1688980957
transform -1 0 34500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold673
timestamp 1688980957
transform -1 0 43792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold674
timestamp 1688980957
transform -1 0 47472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold675
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold676
timestamp 1688980957
transform 1 0 40204 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold677
timestamp 1688980957
transform -1 0 41400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold678
timestamp 1688980957
transform -1 0 39468 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold679
timestamp 1688980957
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold680
timestamp 1688980957
transform -1 0 11224 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold681
timestamp 1688980957
transform -1 0 11040 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold682
timestamp 1688980957
transform -1 0 34316 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold683
timestamp 1688980957
transform -1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold684
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold685
timestamp 1688980957
transform 1 0 45264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold686
timestamp 1688980957
transform 1 0 46000 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold687
timestamp 1688980957
transform -1 0 52440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold688
timestamp 1688980957
transform 1 0 52900 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold689
timestamp 1688980957
transform -1 0 52440 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold690
timestamp 1688980957
transform -1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold691
timestamp 1688980957
transform -1 0 18768 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold692
timestamp 1688980957
transform 1 0 29716 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold693
timestamp 1688980957
transform 1 0 30360 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold694
timestamp 1688980957
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold695
timestamp 1688980957
transform -1 0 58144 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold696
timestamp 1688980957
transform -1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold697
timestamp 1688980957
transform -1 0 13524 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold698
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold699
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold700
timestamp 1688980957
transform 1 0 49128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold701
timestamp 1688980957
transform -1 0 49128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold702
timestamp 1688980957
transform -1 0 3680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold703
timestamp 1688980957
transform -1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold704
timestamp 1688980957
transform -1 0 3312 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold705
timestamp 1688980957
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold706
timestamp 1688980957
transform -1 0 3496 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold707
timestamp 1688980957
transform -1 0 4600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold708
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold709
timestamp 1688980957
transform -1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold710
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold711
timestamp 1688980957
transform -1 0 9568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold712
timestamp 1688980957
transform -1 0 8372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold713
timestamp 1688980957
transform -1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold714
timestamp 1688980957
transform -1 0 14720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold715
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold716
timestamp 1688980957
transform 1 0 28152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold717
timestamp 1688980957
transform -1 0 52072 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold718
timestamp 1688980957
transform -1 0 10856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold719
timestamp 1688980957
transform -1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold720
timestamp 1688980957
transform -1 0 48300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold721
timestamp 1688980957
transform 1 0 16744 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold722
timestamp 1688980957
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold723
timestamp 1688980957
transform 1 0 11040 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold724
timestamp 1688980957
transform 1 0 49680 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold725
timestamp 1688980957
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 35972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 36616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 40112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 43608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 47472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 51980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 55200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 54556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 55568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform -1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1688980957
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform -1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform -1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform -1 0 29348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform -1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 36064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform -1 0 37076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 39468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform -1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform -1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 46920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 46920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 52164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 52256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 55384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 57224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform -1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform -1 0 57684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 58328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 11592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 14168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform -1 0 20976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform -1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1688980957
transform 1 0 1472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output69 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform 1 0 24196 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform 1 0 30544 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 33948 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform -1 0 36156 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform 1 0 40756 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform -1 0 45540 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform -1 0 47196 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform 1 0 47564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform 1 0 49036 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform -1 0 52164 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform 1 0 54004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform -1 0 57132 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform -1 0 57776 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform 1 0 57132 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform -1 0 13984 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire112
timestamp 1688980957
transform -1 0 9384 0 -1 3264
box -38 -48 406 592
<< labels >>
flabel metal4 s 8166 2128 8486 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 22610 2128 22930 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 37054 2128 37374 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 51498 2128 51818 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 15388 2128 15708 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 29832 2128 30152 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 44276 2128 44596 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 58720 2128 59040 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal tristate
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal tristate
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
