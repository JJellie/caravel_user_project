// This is the unpowered netlist.
module wishbone_nn (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \fifo_in.FIFO[0][0] ;
 wire \fifo_in.FIFO[0][10] ;
 wire \fifo_in.FIFO[0][11] ;
 wire \fifo_in.FIFO[0][12] ;
 wire \fifo_in.FIFO[0][13] ;
 wire \fifo_in.FIFO[0][14] ;
 wire \fifo_in.FIFO[0][15] ;
 wire \fifo_in.FIFO[0][16] ;
 wire \fifo_in.FIFO[0][17] ;
 wire \fifo_in.FIFO[0][18] ;
 wire \fifo_in.FIFO[0][19] ;
 wire \fifo_in.FIFO[0][1] ;
 wire \fifo_in.FIFO[0][20] ;
 wire \fifo_in.FIFO[0][21] ;
 wire \fifo_in.FIFO[0][22] ;
 wire \fifo_in.FIFO[0][23] ;
 wire \fifo_in.FIFO[0][24] ;
 wire \fifo_in.FIFO[0][25] ;
 wire \fifo_in.FIFO[0][26] ;
 wire \fifo_in.FIFO[0][27] ;
 wire \fifo_in.FIFO[0][28] ;
 wire \fifo_in.FIFO[0][29] ;
 wire \fifo_in.FIFO[0][2] ;
 wire \fifo_in.FIFO[0][30] ;
 wire \fifo_in.FIFO[0][31] ;
 wire \fifo_in.FIFO[0][3] ;
 wire \fifo_in.FIFO[0][4] ;
 wire \fifo_in.FIFO[0][5] ;
 wire \fifo_in.FIFO[0][6] ;
 wire \fifo_in.FIFO[0][7] ;
 wire \fifo_in.FIFO[0][8] ;
 wire \fifo_in.FIFO[0][9] ;
 wire \fifo_in.FIFO[1][0] ;
 wire \fifo_in.FIFO[1][10] ;
 wire \fifo_in.FIFO[1][11] ;
 wire \fifo_in.FIFO[1][12] ;
 wire \fifo_in.FIFO[1][13] ;
 wire \fifo_in.FIFO[1][14] ;
 wire \fifo_in.FIFO[1][15] ;
 wire \fifo_in.FIFO[1][16] ;
 wire \fifo_in.FIFO[1][17] ;
 wire \fifo_in.FIFO[1][18] ;
 wire \fifo_in.FIFO[1][19] ;
 wire \fifo_in.FIFO[1][1] ;
 wire \fifo_in.FIFO[1][20] ;
 wire \fifo_in.FIFO[1][21] ;
 wire \fifo_in.FIFO[1][22] ;
 wire \fifo_in.FIFO[1][23] ;
 wire \fifo_in.FIFO[1][24] ;
 wire \fifo_in.FIFO[1][25] ;
 wire \fifo_in.FIFO[1][26] ;
 wire \fifo_in.FIFO[1][27] ;
 wire \fifo_in.FIFO[1][28] ;
 wire \fifo_in.FIFO[1][29] ;
 wire \fifo_in.FIFO[1][2] ;
 wire \fifo_in.FIFO[1][30] ;
 wire \fifo_in.FIFO[1][31] ;
 wire \fifo_in.FIFO[1][3] ;
 wire \fifo_in.FIFO[1][4] ;
 wire \fifo_in.FIFO[1][5] ;
 wire \fifo_in.FIFO[1][6] ;
 wire \fifo_in.FIFO[1][7] ;
 wire \fifo_in.FIFO[1][8] ;
 wire \fifo_in.FIFO[1][9] ;
 wire \fifo_in.FIFO[2][0] ;
 wire \fifo_in.FIFO[2][10] ;
 wire \fifo_in.FIFO[2][11] ;
 wire \fifo_in.FIFO[2][12] ;
 wire \fifo_in.FIFO[2][13] ;
 wire \fifo_in.FIFO[2][14] ;
 wire \fifo_in.FIFO[2][15] ;
 wire \fifo_in.FIFO[2][16] ;
 wire \fifo_in.FIFO[2][17] ;
 wire \fifo_in.FIFO[2][18] ;
 wire \fifo_in.FIFO[2][19] ;
 wire \fifo_in.FIFO[2][1] ;
 wire \fifo_in.FIFO[2][20] ;
 wire \fifo_in.FIFO[2][21] ;
 wire \fifo_in.FIFO[2][22] ;
 wire \fifo_in.FIFO[2][23] ;
 wire \fifo_in.FIFO[2][24] ;
 wire \fifo_in.FIFO[2][25] ;
 wire \fifo_in.FIFO[2][26] ;
 wire \fifo_in.FIFO[2][27] ;
 wire \fifo_in.FIFO[2][28] ;
 wire \fifo_in.FIFO[2][29] ;
 wire \fifo_in.FIFO[2][2] ;
 wire \fifo_in.FIFO[2][30] ;
 wire \fifo_in.FIFO[2][31] ;
 wire \fifo_in.FIFO[2][3] ;
 wire \fifo_in.FIFO[2][4] ;
 wire \fifo_in.FIFO[2][5] ;
 wire \fifo_in.FIFO[2][6] ;
 wire \fifo_in.FIFO[2][7] ;
 wire \fifo_in.FIFO[2][8] ;
 wire \fifo_in.FIFO[2][9] ;
 wire \fifo_in.FIFO[3][0] ;
 wire \fifo_in.FIFO[3][10] ;
 wire \fifo_in.FIFO[3][11] ;
 wire \fifo_in.FIFO[3][12] ;
 wire \fifo_in.FIFO[3][13] ;
 wire \fifo_in.FIFO[3][14] ;
 wire \fifo_in.FIFO[3][15] ;
 wire \fifo_in.FIFO[3][16] ;
 wire \fifo_in.FIFO[3][17] ;
 wire \fifo_in.FIFO[3][18] ;
 wire \fifo_in.FIFO[3][19] ;
 wire \fifo_in.FIFO[3][1] ;
 wire \fifo_in.FIFO[3][20] ;
 wire \fifo_in.FIFO[3][21] ;
 wire \fifo_in.FIFO[3][22] ;
 wire \fifo_in.FIFO[3][23] ;
 wire \fifo_in.FIFO[3][24] ;
 wire \fifo_in.FIFO[3][25] ;
 wire \fifo_in.FIFO[3][26] ;
 wire \fifo_in.FIFO[3][27] ;
 wire \fifo_in.FIFO[3][28] ;
 wire \fifo_in.FIFO[3][29] ;
 wire \fifo_in.FIFO[3][2] ;
 wire \fifo_in.FIFO[3][30] ;
 wire \fifo_in.FIFO[3][31] ;
 wire \fifo_in.FIFO[3][3] ;
 wire \fifo_in.FIFO[3][4] ;
 wire \fifo_in.FIFO[3][5] ;
 wire \fifo_in.FIFO[3][6] ;
 wire \fifo_in.FIFO[3][7] ;
 wire \fifo_in.FIFO[3][8] ;
 wire \fifo_in.FIFO[3][9] ;
 wire \fifo_in.FIFO[4][0] ;
 wire \fifo_in.FIFO[4][10] ;
 wire \fifo_in.FIFO[4][11] ;
 wire \fifo_in.FIFO[4][12] ;
 wire \fifo_in.FIFO[4][13] ;
 wire \fifo_in.FIFO[4][14] ;
 wire \fifo_in.FIFO[4][15] ;
 wire \fifo_in.FIFO[4][16] ;
 wire \fifo_in.FIFO[4][17] ;
 wire \fifo_in.FIFO[4][18] ;
 wire \fifo_in.FIFO[4][19] ;
 wire \fifo_in.FIFO[4][1] ;
 wire \fifo_in.FIFO[4][20] ;
 wire \fifo_in.FIFO[4][21] ;
 wire \fifo_in.FIFO[4][22] ;
 wire \fifo_in.FIFO[4][23] ;
 wire \fifo_in.FIFO[4][24] ;
 wire \fifo_in.FIFO[4][25] ;
 wire \fifo_in.FIFO[4][26] ;
 wire \fifo_in.FIFO[4][27] ;
 wire \fifo_in.FIFO[4][28] ;
 wire \fifo_in.FIFO[4][29] ;
 wire \fifo_in.FIFO[4][2] ;
 wire \fifo_in.FIFO[4][30] ;
 wire \fifo_in.FIFO[4][31] ;
 wire \fifo_in.FIFO[4][3] ;
 wire \fifo_in.FIFO[4][4] ;
 wire \fifo_in.FIFO[4][5] ;
 wire \fifo_in.FIFO[4][6] ;
 wire \fifo_in.FIFO[4][7] ;
 wire \fifo_in.FIFO[4][8] ;
 wire \fifo_in.FIFO[4][9] ;
 wire \fifo_in.FIFO[5][0] ;
 wire \fifo_in.FIFO[5][10] ;
 wire \fifo_in.FIFO[5][11] ;
 wire \fifo_in.FIFO[5][12] ;
 wire \fifo_in.FIFO[5][13] ;
 wire \fifo_in.FIFO[5][14] ;
 wire \fifo_in.FIFO[5][15] ;
 wire \fifo_in.FIFO[5][16] ;
 wire \fifo_in.FIFO[5][17] ;
 wire \fifo_in.FIFO[5][18] ;
 wire \fifo_in.FIFO[5][19] ;
 wire \fifo_in.FIFO[5][1] ;
 wire \fifo_in.FIFO[5][20] ;
 wire \fifo_in.FIFO[5][21] ;
 wire \fifo_in.FIFO[5][22] ;
 wire \fifo_in.FIFO[5][23] ;
 wire \fifo_in.FIFO[5][24] ;
 wire \fifo_in.FIFO[5][25] ;
 wire \fifo_in.FIFO[5][26] ;
 wire \fifo_in.FIFO[5][27] ;
 wire \fifo_in.FIFO[5][28] ;
 wire \fifo_in.FIFO[5][29] ;
 wire \fifo_in.FIFO[5][2] ;
 wire \fifo_in.FIFO[5][30] ;
 wire \fifo_in.FIFO[5][31] ;
 wire \fifo_in.FIFO[5][3] ;
 wire \fifo_in.FIFO[5][4] ;
 wire \fifo_in.FIFO[5][5] ;
 wire \fifo_in.FIFO[5][6] ;
 wire \fifo_in.FIFO[5][7] ;
 wire \fifo_in.FIFO[5][8] ;
 wire \fifo_in.FIFO[5][9] ;
 wire \fifo_in.FIFO[6][0] ;
 wire \fifo_in.FIFO[6][10] ;
 wire \fifo_in.FIFO[6][11] ;
 wire \fifo_in.FIFO[6][12] ;
 wire \fifo_in.FIFO[6][13] ;
 wire \fifo_in.FIFO[6][14] ;
 wire \fifo_in.FIFO[6][15] ;
 wire \fifo_in.FIFO[6][16] ;
 wire \fifo_in.FIFO[6][17] ;
 wire \fifo_in.FIFO[6][18] ;
 wire \fifo_in.FIFO[6][19] ;
 wire \fifo_in.FIFO[6][1] ;
 wire \fifo_in.FIFO[6][20] ;
 wire \fifo_in.FIFO[6][21] ;
 wire \fifo_in.FIFO[6][22] ;
 wire \fifo_in.FIFO[6][23] ;
 wire \fifo_in.FIFO[6][24] ;
 wire \fifo_in.FIFO[6][25] ;
 wire \fifo_in.FIFO[6][26] ;
 wire \fifo_in.FIFO[6][27] ;
 wire \fifo_in.FIFO[6][28] ;
 wire \fifo_in.FIFO[6][29] ;
 wire \fifo_in.FIFO[6][2] ;
 wire \fifo_in.FIFO[6][30] ;
 wire \fifo_in.FIFO[6][31] ;
 wire \fifo_in.FIFO[6][3] ;
 wire \fifo_in.FIFO[6][4] ;
 wire \fifo_in.FIFO[6][5] ;
 wire \fifo_in.FIFO[6][6] ;
 wire \fifo_in.FIFO[6][7] ;
 wire \fifo_in.FIFO[6][8] ;
 wire \fifo_in.FIFO[6][9] ;
 wire \fifo_in.FIFO[7][0] ;
 wire \fifo_in.FIFO[7][10] ;
 wire \fifo_in.FIFO[7][11] ;
 wire \fifo_in.FIFO[7][12] ;
 wire \fifo_in.FIFO[7][13] ;
 wire \fifo_in.FIFO[7][14] ;
 wire \fifo_in.FIFO[7][15] ;
 wire \fifo_in.FIFO[7][16] ;
 wire \fifo_in.FIFO[7][17] ;
 wire \fifo_in.FIFO[7][18] ;
 wire \fifo_in.FIFO[7][19] ;
 wire \fifo_in.FIFO[7][1] ;
 wire \fifo_in.FIFO[7][20] ;
 wire \fifo_in.FIFO[7][21] ;
 wire \fifo_in.FIFO[7][22] ;
 wire \fifo_in.FIFO[7][23] ;
 wire \fifo_in.FIFO[7][24] ;
 wire \fifo_in.FIFO[7][25] ;
 wire \fifo_in.FIFO[7][26] ;
 wire \fifo_in.FIFO[7][27] ;
 wire \fifo_in.FIFO[7][28] ;
 wire \fifo_in.FIFO[7][29] ;
 wire \fifo_in.FIFO[7][2] ;
 wire \fifo_in.FIFO[7][30] ;
 wire \fifo_in.FIFO[7][31] ;
 wire \fifo_in.FIFO[7][3] ;
 wire \fifo_in.FIFO[7][4] ;
 wire \fifo_in.FIFO[7][5] ;
 wire \fifo_in.FIFO[7][6] ;
 wire \fifo_in.FIFO[7][7] ;
 wire \fifo_in.FIFO[7][8] ;
 wire \fifo_in.FIFO[7][9] ;
 wire \fifo_in.count[0] ;
 wire \fifo_in.count[1] ;
 wire \fifo_in.count[2] ;
 wire \fifo_in.data_o[0] ;
 wire \fifo_in.data_o[10] ;
 wire \fifo_in.data_o[11] ;
 wire \fifo_in.data_o[12] ;
 wire \fifo_in.data_o[13] ;
 wire \fifo_in.data_o[14] ;
 wire \fifo_in.data_o[15] ;
 wire \fifo_in.data_o[16] ;
 wire \fifo_in.data_o[17] ;
 wire \fifo_in.data_o[18] ;
 wire \fifo_in.data_o[19] ;
 wire \fifo_in.data_o[1] ;
 wire \fifo_in.data_o[20] ;
 wire \fifo_in.data_o[21] ;
 wire \fifo_in.data_o[22] ;
 wire \fifo_in.data_o[23] ;
 wire \fifo_in.data_o[24] ;
 wire \fifo_in.data_o[25] ;
 wire \fifo_in.data_o[26] ;
 wire \fifo_in.data_o[27] ;
 wire \fifo_in.data_o[28] ;
 wire \fifo_in.data_o[29] ;
 wire \fifo_in.data_o[2] ;
 wire \fifo_in.data_o[30] ;
 wire \fifo_in.data_o[31] ;
 wire \fifo_in.data_o[3] ;
 wire \fifo_in.data_o[4] ;
 wire \fifo_in.data_o[5] ;
 wire \fifo_in.data_o[6] ;
 wire \fifo_in.data_o[7] ;
 wire \fifo_in.data_o[8] ;
 wire \fifo_in.data_o[9] ;
 wire \fifo_in.read_addr[0] ;
 wire \fifo_in.read_addr[1] ;
 wire \fifo_in.read_addr[2] ;
 wire \fifo_in.write_addr[0] ;
 wire \fifo_in.write_addr[1] ;
 wire \fifo_in.write_addr[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__0518__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__S (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__D (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0551__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0552__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0553__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0559__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0563__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0578__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__S (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__S (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0616__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0624__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__S (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__S (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__S (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__S (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__S (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__S (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A_N (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__D (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A2 (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__A2 (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0930__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__S (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0951__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0958__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__S (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1282__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1295__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1298__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_98 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _0517_ (.A(net70),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(net123),
    .Y(_0399_));
 sky130_fd_sc_hd__and4bb_1 _0519_ (.A_N(\fifo_in.write_addr[0] ),
    .B_N(net137),
    .C(net34),
    .D(net68),
    .X(_0400_));
 sky130_fd_sc_hd__nor3b_4 _0520_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C_N(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__mux2_1 _0521_ (.A0(net824),
    .A1(net452),
    .S(_0401_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0522_ (.A0(net839),
    .A1(net541),
    .S(net121),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0523_ (.A0(net558),
    .A1(net538),
    .S(net121),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0524_ (.A0(net383),
    .A1(net246),
    .S(net121),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0525_ (.A0(net259),
    .A1(net204),
    .S(net121),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0526_ (.A0(net292),
    .A1(net253),
    .S(net121),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0527_ (.A0(net790),
    .A1(net230),
    .S(net121),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0528_ (.A0(net525),
    .A1(net465),
    .S(net121),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _0529_ (.A(\fifo_in.write_addr[0] ),
    .B(net68),
    .C(net34),
    .X(_0402_));
 sky130_fd_sc_hd__nand3_2 _0530_ (.A(\fifo_in.write_addr[0] ),
    .B(net68),
    .C(net34),
    .Y(_0403_));
 sky130_fd_sc_hd__a21o_1 _0531_ (.A1(net68),
    .A2(net34),
    .B1(\fifo_in.write_addr[0] ),
    .X(_0404_));
 sky130_fd_sc_hd__and3b_1 _0532_ (.A_N(net137),
    .B(net844),
    .C(_0404_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _0533_ (.A(net841),
    .B(_0402_),
    .X(_0405_));
 sky130_fd_sc_hd__nor2_1 _0534_ (.A(net137),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__o21a_1 _0535_ (.A1(net841),
    .A2(_0402_),
    .B1(_0406_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _0536_ (.A(net846),
    .B(_0405_),
    .Y(_0407_));
 sky130_fd_sc_hd__or2_1 _0537_ (.A(net846),
    .B(_0405_),
    .X(_0408_));
 sky130_fd_sc_hd__and3b_1 _0538_ (.A_N(net137),
    .B(net847),
    .C(_0408_),
    .X(_0010_));
 sky130_fd_sc_hd__or3_1 _0539_ (.A(net773),
    .B(net760),
    .C(net771),
    .X(_0409_));
 sky130_fd_sc_hd__and3b_1 _0540_ (.A_N(net68),
    .B(net34),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__and4b_1 _0541_ (.A_N(net68),
    .B(net34),
    .C(_0409_),
    .D(net130),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _0542_ (.A(net137),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__o21a_1 _0543_ (.A1(net130),
    .A2(_0410_),
    .B1(_0412_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0544_ (.A(net125),
    .B(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _0545_ (.A(net125),
    .B(_0411_),
    .Y(_0414_));
 sky130_fd_sc_hd__and3b_1 _0546_ (.A_N(net137),
    .B(_0413_),
    .C(_0414_),
    .X(_0012_));
 sky130_fd_sc_hd__a21oi_1 _0547_ (.A1(_0399_),
    .A2(_0414_),
    .B1(net137),
    .Y(_0415_));
 sky130_fd_sc_hd__o21a_1 _0548_ (.A1(_0399_),
    .A2(_0414_),
    .B1(_0415_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_4 _0549_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0400_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _0550_ (.A0(net449),
    .A1(net273),
    .S(net120),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(net220),
    .A1(net209),
    .S(net120),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0552_ (.A0(net588),
    .A1(net474),
    .S(net120),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0553_ (.A0(net492),
    .A1(net415),
    .S(net120),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0554_ (.A0(net371),
    .A1(net339),
    .S(net120),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0555_ (.A0(net361),
    .A1(net336),
    .S(net120),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(net498),
    .A1(net276),
    .S(net120),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0557_ (.A0(net311),
    .A1(net187),
    .S(net120),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net278),
    .A1(net243),
    .S(net120),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0559_ (.A0(net412),
    .A1(net398),
    .S(net120),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(net355),
    .A1(net157),
    .S(net120),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0561_ (.A0(net482),
    .A1(net227),
    .S(net120),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0562_ (.A0(net625),
    .A1(net609),
    .S(net120),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(net654),
    .A1(net636),
    .S(net120),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0564_ (.A0(net596),
    .A1(net175),
    .S(net120),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0565_ (.A0(net523),
    .A1(net164),
    .S(net119),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(net319),
    .A1(net268),
    .S(net119),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0567_ (.A0(net531),
    .A1(net501),
    .S(net119),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0568_ (.A0(net576),
    .A1(net548),
    .S(net119),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0569_ (.A0(net469),
    .A1(net152),
    .S(net119),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(net467),
    .A1(net295),
    .S(net119),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0571_ (.A0(net299),
    .A1(net145),
    .S(net119),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(net408),
    .A1(net184),
    .S(net119),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0573_ (.A0(net389),
    .A1(net212),
    .S(net119),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(net644),
    .A1(net452),
    .S(net119),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0575_ (.A0(net594),
    .A1(net541),
    .S(net119),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0576_ (.A0(net621),
    .A1(net538),
    .S(net119),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0577_ (.A0(net404),
    .A1(net246),
    .S(net119),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(net248),
    .A1(net204),
    .S(net119),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(net317),
    .A1(net253),
    .S(net119),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0580_ (.A0(net359),
    .A1(net230),
    .S(net119),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0581_ (.A0(net598),
    .A1(net465),
    .S(_0416_),
    .X(_0045_));
 sky130_fd_sc_hd__or4b_4 _0582_ (.A(\fifo_in.write_addr[1] ),
    .B(net137),
    .C(_0403_),
    .D_N(\fifo_in.write_addr[2] ),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _0583_ (.A0(net273),
    .A1(net410),
    .S(net118),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net209),
    .A1(net323),
    .S(net118),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(net474),
    .A1(net535),
    .S(net118),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net415),
    .A1(net421),
    .S(net118),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(net339),
    .A1(net365),
    .S(net118),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0588_ (.A0(net336),
    .A1(net613),
    .S(net118),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(net276),
    .A1(net513),
    .S(net118),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net187),
    .A1(net270),
    .S(net118),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net243),
    .A1(net429),
    .S(net118),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(net398),
    .A1(net619),
    .S(net118),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net157),
    .A1(net503),
    .S(net118),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net227),
    .A1(net802),
    .S(net118),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(net609),
    .A1(net648),
    .S(net118),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net636),
    .A1(net666),
    .S(net117),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net175),
    .A1(net602),
    .S(net118),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net164),
    .A1(net486),
    .S(net117),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net268),
    .A1(net810),
    .S(net117),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net501),
    .A1(net533),
    .S(net117),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(net548),
    .A1(net684),
    .S(net117),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net152),
    .A1(net433),
    .S(net117),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0603_ (.A0(net295),
    .A1(net456),
    .S(net117),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(net145),
    .A1(net257),
    .S(net117),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(net184),
    .A1(net385),
    .S(net117),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0606_ (.A0(net212),
    .A1(net369),
    .S(net117),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(net452),
    .A1(net600),
    .S(net117),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0608_ (.A0(net541),
    .A1(net578),
    .S(net117),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0609_ (.A0(net538),
    .A1(net640),
    .S(net117),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(net246),
    .A1(net400),
    .S(net117),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0611_ (.A0(net204),
    .A1(net781),
    .S(net117),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0612_ (.A0(net253),
    .A1(net309),
    .S(net117),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0613_ (.A0(net230),
    .A1(net325),
    .S(_0417_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(net465),
    .A1(net586),
    .S(net118),
    .X(_0077_));
 sky130_fd_sc_hd__and3b_4 _0615_ (.A_N(\fifo_in.write_addr[1] ),
    .B(_0400_),
    .C(\fifo_in.write_addr[2] ),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _0616_ (.A0(net431),
    .A1(net273),
    .S(net116),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(net232),
    .A1(net209),
    .S(net116),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(net543),
    .A1(net474),
    .S(net116),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(net462),
    .A1(net415),
    .S(net116),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(net375),
    .A1(net339),
    .S(net116),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(net393),
    .A1(net336),
    .S(net116),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(net443),
    .A1(net276),
    .S(net116),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(net439),
    .A1(net187),
    .S(net116),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(net852),
    .A1(net243),
    .S(net116),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0625_ (.A0(net680),
    .A1(net398),
    .S(net116),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(net379),
    .A1(net157),
    .S(net116),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(net307),
    .A1(net227),
    .S(net116),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(net629),
    .A1(net609),
    .S(net116),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(net682),
    .A1(net636),
    .S(net116),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(net556),
    .A1(net175),
    .S(net116),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0631_ (.A0(net568),
    .A1(net164),
    .S(net115),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(net331),
    .A1(net268),
    .S(net115),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(net550),
    .A1(net501),
    .S(net115),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(net686),
    .A1(net548),
    .S(net115),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(net476),
    .A1(net152),
    .S(net115),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net488),
    .A1(net295),
    .S(net115),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0637_ (.A0(net288),
    .A1(net145),
    .S(net115),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(net280),
    .A1(net184),
    .S(net115),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(net377),
    .A1(net212),
    .S(net115),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0640_ (.A0(net642),
    .A1(net452),
    .S(net115),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0641_ (.A0(net604),
    .A1(net541),
    .S(net115),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(net611),
    .A1(net538),
    .S(net115),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(net406),
    .A1(net246),
    .S(net115),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0644_ (.A0(net250),
    .A1(net204),
    .S(net115),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0645_ (.A0(net343),
    .A1(net253),
    .S(net115),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net351),
    .A1(net230),
    .S(net115),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(net627),
    .A1(net465),
    .S(_0418_),
    .X(_0109_));
 sky130_fd_sc_hd__nand2b_4 _0648_ (.A_N(net137),
    .B(_0410_),
    .Y(_0419_));
 sky130_fd_sc_hd__mux4_1 _0649_ (.A0(net431),
    .A1(net410),
    .A2(net449),
    .A3(net505),
    .S0(net130),
    .S1(net125),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_1 _0650_ (.A0(net301),
    .A1(\fifo_in.FIFO[1][0] ),
    .A2(net282),
    .A3(net315),
    .S0(net130),
    .S1(net125),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _0651_ (.A0(_0421_),
    .A1(_0420_),
    .S(net123),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(_0422_),
    .A1(net804),
    .S(net105),
    .X(_0110_));
 sky130_fd_sc_hd__mux4_1 _0653_ (.A0(net232),
    .A1(net323),
    .A2(net220),
    .A3(net363),
    .S0(net130),
    .S1(net125),
    .X(_0423_));
 sky130_fd_sc_hd__mux4_1 _0654_ (.A0(net224),
    .A1(net234),
    .A2(net218),
    .A3(net796),
    .S0(net130),
    .S1(net125),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(_0424_),
    .A1(_0423_),
    .S(net123),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(net797),
    .A1(net704),
    .S(net105),
    .X(_0111_));
 sky130_fd_sc_hd__mux4_1 _0657_ (.A0(net543),
    .A1(net535),
    .A2(net588),
    .A3(net529),
    .S0(net130),
    .S1(net125),
    .X(_0426_));
 sky130_fd_sc_hd__mux4_1 _0658_ (.A0(net517),
    .A1(net819),
    .A2(net564),
    .A3(net494),
    .S0(net130),
    .S1(net125),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(_0427_),
    .A1(_0426_),
    .S(net123),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net820),
    .A1(net706),
    .S(net105),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_1 _0661_ (.A0(net462),
    .A1(net421),
    .A2(net492),
    .A3(net545),
    .S0(net130),
    .S1(net125),
    .X(_0429_));
 sky130_fd_sc_hd__mux4_1 _0662_ (.A0(net478),
    .A1(net837),
    .A2(net507),
    .A3(net441),
    .S0(net131),
    .S1(net125),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _0663_ (.A0(_0430_),
    .A1(_0429_),
    .S(net123),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(net838),
    .A1(net702),
    .S(net105),
    .X(_0113_));
 sky130_fd_sc_hd__mux4_1 _0665_ (.A0(net375),
    .A1(net365),
    .A2(net371),
    .A3(net381),
    .S0(net130),
    .S1(net125),
    .X(_0432_));
 sky130_fd_sc_hd__mux4_1 _0666_ (.A0(net511),
    .A1(\fifo_in.FIFO[1][4] ),
    .A2(net353),
    .A3(net347),
    .S0(net130),
    .S1(net125),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(_0433_),
    .A1(_0432_),
    .S(net123),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _0668_ (.A0(_0434_),
    .A1(net835),
    .S(net105),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _0669_ (.A0(net393),
    .A1(net613),
    .A2(net361),
    .A3(net395),
    .S0(net131),
    .S1(net126),
    .X(_0435_));
 sky130_fd_sc_hd__mux4_1 _0670_ (.A0(net617),
    .A1(net345),
    .A2(net367),
    .A3(net829),
    .S0(net134),
    .S1(net126),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(net830),
    .A1(_0435_),
    .S(net123),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(_0437_),
    .A1(net700),
    .S(net105),
    .X(_0115_));
 sky130_fd_sc_hd__mux4_1 _0673_ (.A0(net443),
    .A1(net513),
    .A2(net498),
    .A3(net427),
    .S0(net130),
    .S1(net125),
    .X(_0438_));
 sky130_fd_sc_hd__mux4_1 _0674_ (.A0(net313),
    .A1(net808),
    .A2(net329),
    .A3(net286),
    .S0(net130),
    .S1(net125),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _0675_ (.A0(_0439_),
    .A1(_0438_),
    .S(net123),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _0676_ (.A0(net809),
    .A1(net708),
    .S(net105),
    .X(_0116_));
 sky130_fd_sc_hd__mux4_1 _0677_ (.A0(net439),
    .A1(net270),
    .A2(net311),
    .A3(net303),
    .S0(net130),
    .S1(net126),
    .X(_0441_));
 sky130_fd_sc_hd__mux4_1 _0678_ (.A0(net197),
    .A1(net199),
    .A2(net201),
    .A3(net765),
    .S0(net131),
    .S1(net126),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(_0442_),
    .A1(_0441_),
    .S(net123),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _0680_ (.A0(net766),
    .A1(net750),
    .S(net105),
    .X(_0117_));
 sky130_fd_sc_hd__mux4_1 _0681_ (.A0(\fifo_in.FIFO[4][8] ),
    .A1(net429),
    .A2(net278),
    .A3(net423),
    .S0(net131),
    .S1(net126),
    .X(_0444_));
 sky130_fd_sc_hd__mux4_1 _0682_ (.A0(net437),
    .A1(net402),
    .A2(net425),
    .A3(net391),
    .S0(net131),
    .S1(net126),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _0683_ (.A0(_0445_),
    .A1(_0444_),
    .S(net799),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(net800),
    .A1(net746),
    .S(net105),
    .X(_0118_));
 sky130_fd_sc_hd__mux4_1 _0685_ (.A0(net680),
    .A1(net619),
    .A2(net412),
    .A3(net823),
    .S0(net131),
    .S1(net126),
    .X(_0447_));
 sky130_fd_sc_hd__mux4_1 _0686_ (.A0(net674),
    .A1(net615),
    .A2(net662),
    .A3(net562),
    .S0(net131),
    .S1(net126),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(_0448_),
    .A1(_0447_),
    .S(net123),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(_0449_),
    .A1(net726),
    .S(net105),
    .X(_0119_));
 sky130_fd_sc_hd__mux4_1 _0689_ (.A0(net379),
    .A1(net503),
    .A2(net355),
    .A3(net349),
    .S0(net131),
    .S1(net126),
    .X(_0450_));
 sky130_fd_sc_hd__mux4_1 _0690_ (.A0(net787),
    .A1(net177),
    .A2(net166),
    .A3(net159),
    .S0(net131),
    .S1(net126),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(_0451_),
    .A1(_0450_),
    .S(net123),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(net788),
    .A1(net752),
    .S(net105),
    .X(_0120_));
 sky130_fd_sc_hd__mux4_1 _0693_ (.A0(net307),
    .A1(net802),
    .A2(net482),
    .A3(net471),
    .S0(net131),
    .S1(net126),
    .X(_0453_));
 sky130_fd_sc_hd__mux4_1 _0694_ (.A0(net490),
    .A1(net419),
    .A2(net458),
    .A3(net447),
    .S0(net131),
    .S1(net126),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(_0454_),
    .A1(_0453_),
    .S(net123),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(net803),
    .A1(net748),
    .S(net105),
    .X(_0121_));
 sky130_fd_sc_hd__mux4_1 _0697_ (.A0(net629),
    .A1(net648),
    .A2(net625),
    .A3(net650),
    .S0(net131),
    .S1(net126),
    .X(_0456_));
 sky130_fd_sc_hd__mux4_1 _0698_ (.A0(net631),
    .A1(net664),
    .A2(net652),
    .A3(net818),
    .S0(net131),
    .S1(net126),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(_0457_),
    .A1(_0456_),
    .S(net123),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(_0458_),
    .A1(net736),
    .S(net105),
    .X(_0122_));
 sky130_fd_sc_hd__mux4_1 _0701_ (.A0(net682),
    .A1(net666),
    .A2(net654),
    .A3(net676),
    .S0(net133),
    .S1(net128),
    .X(_0459_));
 sky130_fd_sc_hd__mux4_1 _0702_ (.A0(net672),
    .A1(net668),
    .A2(net660),
    .A3(net831),
    .S0(net133),
    .S1(net128),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(_0460_),
    .A1(_0459_),
    .S(net799),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(net832),
    .A1(net754),
    .S(net105),
    .X(_0123_));
 sky130_fd_sc_hd__mux4_1 _0705_ (.A0(net556),
    .A1(net602),
    .A2(net596),
    .A3(net580),
    .S0(net131),
    .S1(net126),
    .X(_0462_));
 sky130_fd_sc_hd__mux4_1 _0706_ (.A0(net214),
    .A1(net195),
    .A2(net191),
    .A3(net762),
    .S0(net131),
    .S1(net126),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(_0463_),
    .A1(_0462_),
    .S(net123),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(net763),
    .A1(net732),
    .S(net105),
    .X(_0124_));
 sky130_fd_sc_hd__mux4_1 _0709_ (.A0(net568),
    .A1(net486),
    .A2(net523),
    .A3(net521),
    .S0(net133),
    .S1(net128),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_1 _0710_ (.A0(net181),
    .A1(net775),
    .A2(net179),
    .A3(net168),
    .S0(net133),
    .S1(net128),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(_0466_),
    .A1(_0465_),
    .S(net124),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _0712_ (.A0(net776),
    .A1(net758),
    .S(net104),
    .X(_0125_));
 sky130_fd_sc_hd__mux4_1 _0713_ (.A0(net331),
    .A1(net810),
    .A2(net319),
    .A3(net321),
    .S0(net133),
    .S1(net128),
    .X(_0468_));
 sky130_fd_sc_hd__mux4_1 _0714_ (.A0(net515),
    .A1(net566),
    .A2(net584),
    .A3(net606),
    .S0(net133),
    .S1(net128),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(_0469_),
    .A1(_0468_),
    .S(net124),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(net811),
    .A1(net756),
    .S(net104),
    .X(_0126_));
 sky130_fd_sc_hd__mux4_1 _0717_ (.A0(net550),
    .A1(net533),
    .A2(net531),
    .A3(net572),
    .S0(net133),
    .S1(net128),
    .X(_0471_));
 sky130_fd_sc_hd__mux4_1 _0718_ (.A0(net554),
    .A1(net509),
    .A2(net560),
    .A3(net821),
    .S0(net133),
    .S1(net128),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(_0472_),
    .A1(_0471_),
    .S(net124),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(net822),
    .A1(net714),
    .S(net104),
    .X(_0127_));
 sky130_fd_sc_hd__mux4_1 _0721_ (.A0(net686),
    .A1(net684),
    .A2(net576),
    .A3(net570),
    .S0(net133),
    .S1(net128),
    .X(_0474_));
 sky130_fd_sc_hd__mux4_1 _0722_ (.A0(net574),
    .A1(net816),
    .A2(net582),
    .A3(net590),
    .S0(net133),
    .S1(net128),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(_0475_),
    .A1(_0474_),
    .S(net124),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(net817),
    .A1(net734),
    .S(net104),
    .X(_0128_));
 sky130_fd_sc_hd__mux4_1 _0725_ (.A0(net476),
    .A1(net433),
    .A2(net469),
    .A3(net552),
    .S0(net133),
    .S1(net128),
    .X(_0477_));
 sky130_fd_sc_hd__mux4_1 _0726_ (.A0(net161),
    .A1(net768),
    .A2(net170),
    .A3(net154),
    .S0(net133),
    .S1(net128),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(_0478_),
    .A1(_0477_),
    .S(net124),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net769),
    .A1(net710),
    .S(net104),
    .X(_0129_));
 sky130_fd_sc_hd__mux4_1 _0729_ (.A0(net488),
    .A1(net456),
    .A2(net467),
    .A3(net519),
    .S0(net133),
    .S1(net128),
    .X(_0480_));
 sky130_fd_sc_hd__mux4_1 _0730_ (.A0(net341),
    .A1(net305),
    .A2(net333),
    .A3(net814),
    .S0(net133),
    .S1(net128),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(_0481_),
    .A1(_0480_),
    .S(net124),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net815),
    .A1(net720),
    .S(net104),
    .X(_0130_));
 sky130_fd_sc_hd__mux4_1 _0733_ (.A0(net288),
    .A1(net257),
    .A2(net299),
    .A3(net435),
    .S0(net133),
    .S1(net128),
    .X(_0483_));
 sky130_fd_sc_hd__mux4_1 _0734_ (.A0(net172),
    .A1(net147),
    .A2(net149),
    .A3(net784),
    .S0(net133),
    .S1(net128),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(_0484_),
    .A1(_0483_),
    .S(net124),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net785),
    .A1(net724),
    .S(net104),
    .X(_0131_));
 sky130_fd_sc_hd__mux4_1 _0737_ (.A0(net280),
    .A1(net385),
    .A2(net408),
    .A3(net417),
    .S0(net132),
    .S1(net127),
    .X(_0486_));
 sky130_fd_sc_hd__mux4_1 _0738_ (.A0(net216),
    .A1(net189),
    .A2(net193),
    .A3(net778),
    .S0(net132),
    .S1(net127),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(_0487_),
    .A1(_0486_),
    .S(net124),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net779),
    .A1(net742),
    .S(net104),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_1 _0741_ (.A0(net377),
    .A1(net369),
    .A2(net389),
    .A3(net445),
    .S0(net134),
    .S1(net129),
    .X(_0489_));
 sky130_fd_sc_hd__mux4_1 _0742_ (.A0(net265),
    .A1(net812),
    .A2(net240),
    .A3(net236),
    .S0(net132),
    .S1(net127),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(_0490_),
    .A1(_0489_),
    .S(net124),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(net813),
    .A1(net730),
    .S(net104),
    .X(_0133_));
 sky130_fd_sc_hd__mux4_1 _0745_ (.A0(net642),
    .A1(net600),
    .A2(net644),
    .A3(net670),
    .S0(net132),
    .S1(net127),
    .X(_0492_));
 sky130_fd_sc_hd__mux4_1 _0746_ (.A0(net824),
    .A1(net454),
    .A2(net460),
    .A3(net480),
    .S0(net132),
    .S1(net127),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(_0493_),
    .A1(_0492_),
    .S(net124),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(net825),
    .A1(net728),
    .S(net104),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _0749_ (.A0(net604),
    .A1(net578),
    .A2(net594),
    .A3(net623),
    .S0(net132),
    .S1(net127),
    .X(_0495_));
 sky130_fd_sc_hd__mux4_1 _0750_ (.A0(net839),
    .A1(net656),
    .A2(net678),
    .A3(net658),
    .S0(net132),
    .S1(net127),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(_0496_),
    .A1(_0495_),
    .S(net124),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(net840),
    .A1(net712),
    .S(net104),
    .X(_0135_));
 sky130_fd_sc_hd__mux4_1 _0753_ (.A0(net611),
    .A1(net640),
    .A2(net621),
    .A3(net646),
    .S0(net134),
    .S1(net129),
    .X(_0498_));
 sky130_fd_sc_hd__mux4_1 _0754_ (.A0(net558),
    .A1(net633),
    .A2(net826),
    .A3(net592),
    .S0(net134),
    .S1(net129),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(net827),
    .A1(_0498_),
    .S(net124),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(net828),
    .A1(net722),
    .S(net104),
    .X(_0136_));
 sky130_fd_sc_hd__mux4_1 _0757_ (.A0(net406),
    .A1(net400),
    .A2(net404),
    .A3(net496),
    .S0(net134),
    .S1(net129),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _0758_ (.A0(net383),
    .A1(net806),
    .A2(net284),
    .A3(net373),
    .S0(net132),
    .S1(net127),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _0759_ (.A0(_0502_),
    .A1(_0501_),
    .S(net124),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(net807),
    .A1(net744),
    .S(net104),
    .X(_0137_));
 sky130_fd_sc_hd__mux4_1 _0761_ (.A0(net250),
    .A1(net781),
    .A2(net248),
    .A3(net387),
    .S0(net132),
    .S1(net127),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _0762_ (.A0(net259),
    .A1(net222),
    .A2(net263),
    .A3(net206),
    .S0(net132),
    .S1(net127),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _0763_ (.A0(_0505_),
    .A1(_0504_),
    .S(net124),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(net782),
    .A1(net738),
    .S(net104),
    .X(_0138_));
 sky130_fd_sc_hd__mux4_1 _0765_ (.A0(net343),
    .A1(net309),
    .A2(net317),
    .A3(net297),
    .S0(net132),
    .S1(net127),
    .X(_0507_));
 sky130_fd_sc_hd__mux4_1 _0766_ (.A0(net292),
    .A1(net793),
    .A2(net290),
    .A3(net255),
    .S0(net132),
    .S1(net127),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(_0508_),
    .A1(_0507_),
    .S(net124),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(net794),
    .A1(net740),
    .S(net104),
    .X(_0139_));
 sky130_fd_sc_hd__mux4_1 _0769_ (.A0(net351),
    .A1(net325),
    .A2(net359),
    .A3(net357),
    .S0(net132),
    .S1(net127),
    .X(_0510_));
 sky130_fd_sc_hd__mux4_1 _0770_ (.A0(net790),
    .A1(net327),
    .A2(net238),
    .A3(net261),
    .S0(net132),
    .S1(net127),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(_0511_),
    .A1(_0510_),
    .S(net124),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(net791),
    .A1(net716),
    .S(net104),
    .X(_0140_));
 sky130_fd_sc_hd__mux4_1 _0773_ (.A0(net627),
    .A1(net586),
    .A2(net598),
    .A3(net638),
    .S0(net132),
    .S1(net127),
    .X(_0513_));
 sky130_fd_sc_hd__mux4_1 _0774_ (.A0(net525),
    .A1(net833),
    .A2(net527),
    .A3(net484),
    .S0(net132),
    .S1(net127),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(_0514_),
    .A1(_0513_),
    .S(net799),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(net834),
    .A1(net718),
    .S(_0419_),
    .X(_0141_));
 sky130_fd_sc_hd__or4b_4 _0777_ (.A(\fifo_in.write_addr[2] ),
    .B(net137),
    .C(_0403_),
    .D_N(\fifo_in.write_addr[1] ),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(net273),
    .A1(net315),
    .S(net114),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(net209),
    .A1(net796),
    .S(net114),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(net474),
    .A1(net494),
    .S(net114),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(net415),
    .A1(net441),
    .S(net114),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(net339),
    .A1(net347),
    .S(net114),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(net336),
    .A1(net829),
    .S(net114),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(net276),
    .A1(net286),
    .S(net114),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(net187),
    .A1(net765),
    .S(net114),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(net243),
    .A1(net391),
    .S(net114),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(net398),
    .A1(net562),
    .S(net114),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(net157),
    .A1(net159),
    .S(net114),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net227),
    .A1(net447),
    .S(net114),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(net609),
    .A1(net818),
    .S(net114),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(net636),
    .A1(net831),
    .S(net114),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net175),
    .A1(net762),
    .S(net114),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(net164),
    .A1(net168),
    .S(net113),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(net268),
    .A1(net606),
    .S(net113),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(net501),
    .A1(net821),
    .S(net113),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(net548),
    .A1(net590),
    .S(net113),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(net152),
    .A1(net154),
    .S(net113),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0798_ (.A0(net295),
    .A1(net814),
    .S(net113),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0799_ (.A0(net145),
    .A1(net784),
    .S(net113),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(net184),
    .A1(net778),
    .S(net113),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(net212),
    .A1(net236),
    .S(net113),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _0802_ (.A0(net452),
    .A1(net480),
    .S(net113),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(net541),
    .A1(net658),
    .S(net113),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(net538),
    .A1(net592),
    .S(net113),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(net246),
    .A1(net373),
    .S(net113),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(net204),
    .A1(net206),
    .S(net113),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _0807_ (.A0(net253),
    .A1(net255),
    .S(net113),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(net230),
    .A1(net261),
    .S(net113),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(net465),
    .A1(net484),
    .S(_0516_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2b_1 _0810_ (.A_N(\fifo_in.write_addr[0] ),
    .B(net130),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2b_1 _0811_ (.A_N(net130),
    .B(\fifo_in.write_addr[0] ),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_2 _0812_ (.A(_0330_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__and2b_1 _0813_ (.A_N(net125),
    .B(\fifo_in.write_addr[1] ),
    .X(_0333_));
 sky130_fd_sc_hd__xnor2_2 _0814_ (.A(net125),
    .B(\fifo_in.write_addr[1] ),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2b_1 _0816_ (.A_N(net123),
    .B(\fifo_in.write_addr[2] ),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2b_1 _0817_ (.A_N(\fifo_in.write_addr[2] ),
    .B(net123),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _0818_ (.A(_0336_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__nor4_1 _0819_ (.A(net137),
    .B(_0332_),
    .C(_0335_),
    .D(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__a21o_1 _0820_ (.A1(net760),
    .A2(_0339_),
    .B1(_0332_),
    .X(_0174_));
 sky130_fd_sc_hd__xor2_1 _0821_ (.A(_0330_),
    .B(_0334_),
    .X(_0340_));
 sky130_fd_sc_hd__a21oi_1 _0822_ (.A1(_0330_),
    .A2(_0334_),
    .B1(_0333_),
    .Y(_0341_));
 sky130_fd_sc_hd__or2_1 _0823_ (.A(_0338_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a31o_1 _0824_ (.A1(_0332_),
    .A2(_0336_),
    .A3(_0342_),
    .B1(_0340_),
    .X(_0343_));
 sky130_fd_sc_hd__nand4_1 _0825_ (.A(_0332_),
    .B(_0336_),
    .C(_0340_),
    .D(_0342_),
    .Y(_0344_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(net773),
    .A2(_0339_),
    .B1(_0343_),
    .B2(_0344_),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _0827_ (.A(_0338_),
    .B(_0341_),
    .Y(_0345_));
 sky130_fd_sc_hd__o221a_1 _0828_ (.A1(_0332_),
    .A2(_0335_),
    .B1(_0338_),
    .B2(_0341_),
    .C1(_0336_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _0829_ (.A(_0345_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__a21o_1 _0830_ (.A1(_0342_),
    .A2(_0345_),
    .B1(_0346_),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _0831_ (.A1(net771),
    .A2(_0339_),
    .B1(_0347_),
    .B2(_0348_),
    .X(_0176_));
 sky130_fd_sc_hd__or4_1 _0832_ (.A(net14),
    .B(net17),
    .C(net695),
    .D(net19),
    .X(_0349_));
 sky130_fd_sc_hd__or4_1 _0833_ (.A(net9),
    .B(net12),
    .C(net11),
    .D(net15),
    .X(_0350_));
 sky130_fd_sc_hd__or4b_1 _0834_ (.A(net18),
    .B(net21),
    .C(net20),
    .D_N(net23),
    .X(_0351_));
 sky130_fd_sc_hd__or3b_1 _0835_ (.A(net26),
    .B(net25),
    .C_N(net22),
    .X(_0352_));
 sky130_fd_sc_hd__or4_1 _0836_ (.A(net696),
    .B(_0350_),
    .C(_0351_),
    .D(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__or4_1 _0837_ (.A(net28),
    .B(net31),
    .C(net689),
    .D(net33),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _0838_ (.A(net13),
    .B(net27),
    .C(net24),
    .D(net29),
    .X(_0355_));
 sky130_fd_sc_hd__or4_1 _0839_ (.A(net32),
    .B(net4),
    .C(net3),
    .D(net6),
    .X(_0356_));
 sky130_fd_sc_hd__or4_1 _0840_ (.A(net5),
    .B(net8),
    .C(net7),
    .D(net10),
    .X(_0357_));
 sky130_fd_sc_hd__or4_1 _0841_ (.A(net690),
    .B(_0355_),
    .C(_0356_),
    .D(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__nor2_1 _0842_ (.A(net697),
    .B(net691),
    .Y(_0359_));
 sky130_fd_sc_hd__nand3b_4 _0843_ (.A_N(net68),
    .B(net34),
    .C(net67),
    .Y(_0360_));
 sky130_fd_sc_hd__o21a_1 _0844_ (.A1(net141),
    .A2(\fifo_in.data_o[0] ),
    .B1(net692),
    .X(_0361_));
 sky130_fd_sc_hd__a21oi_1 _0845_ (.A1(_0398_),
    .A2(net135),
    .B1(net137),
    .Y(_0362_));
 sky130_fd_sc_hd__o21a_1 _0846_ (.A1(net135),
    .A2(net142),
    .B1(_0362_),
    .X(_0177_));
 sky130_fd_sc_hd__nor4_1 _0847_ (.A(net141),
    .B(net697),
    .C(net691),
    .D(net135),
    .Y(_0363_));
 sky130_fd_sc_hd__a22oi_1 _0848_ (.A1(net81),
    .A2(net135),
    .B1(net110),
    .B2(net704),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _0849_ (.A(net137),
    .B(net705),
    .Y(_0178_));
 sky130_fd_sc_hd__a22oi_1 _0850_ (.A1(net92),
    .A2(net135),
    .B1(net110),
    .B2(net706),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _0851_ (.A(net137),
    .B(net707),
    .Y(_0179_));
 sky130_fd_sc_hd__a22oi_1 _0852_ (.A1(net95),
    .A2(net135),
    .B1(net110),
    .B2(net702),
    .Y(_0366_));
 sky130_fd_sc_hd__nor2_1 _0853_ (.A(net138),
    .B(net703),
    .Y(_0180_));
 sky130_fd_sc_hd__a22oi_1 _0854_ (.A1(net96),
    .A2(net135),
    .B1(net110),
    .B2(\fifo_in.data_o[4] ),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(net138),
    .B(net699),
    .Y(_0181_));
 sky130_fd_sc_hd__a22oi_1 _0856_ (.A1(net97),
    .A2(net135),
    .B1(net110),
    .B2(net700),
    .Y(_0368_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(net138),
    .B(net701),
    .Y(_0182_));
 sky130_fd_sc_hd__a22oi_1 _0858_ (.A1(net98),
    .A2(net135),
    .B1(net110),
    .B2(net708),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _0859_ (.A(net138),
    .B(net709),
    .Y(_0183_));
 sky130_fd_sc_hd__a22oi_1 _0860_ (.A1(net99),
    .A2(_0360_),
    .B1(net110),
    .B2(net750),
    .Y(_0370_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(net138),
    .B(net751),
    .Y(_0184_));
 sky130_fd_sc_hd__a22oi_1 _0862_ (.A1(net100),
    .A2(net135),
    .B1(net110),
    .B2(net746),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _0863_ (.A(net138),
    .B(net747),
    .Y(_0185_));
 sky130_fd_sc_hd__a22oi_1 _0864_ (.A1(net101),
    .A2(net135),
    .B1(net110),
    .B2(net726),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_1 _0865_ (.A(net138),
    .B(net727),
    .Y(_0186_));
 sky130_fd_sc_hd__a22oi_1 _0866_ (.A1(net71),
    .A2(net135),
    .B1(net110),
    .B2(net752),
    .Y(_0373_));
 sky130_fd_sc_hd__nor2_1 _0867_ (.A(net138),
    .B(net753),
    .Y(_0187_));
 sky130_fd_sc_hd__a22oi_1 _0868_ (.A1(net72),
    .A2(net135),
    .B1(net110),
    .B2(net748),
    .Y(_0374_));
 sky130_fd_sc_hd__nor2_1 _0869_ (.A(net138),
    .B(net749),
    .Y(_0188_));
 sky130_fd_sc_hd__a22oi_1 _0870_ (.A1(net73),
    .A2(net135),
    .B1(net110),
    .B2(net736),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_1 _0871_ (.A(net138),
    .B(net737),
    .Y(_0189_));
 sky130_fd_sc_hd__a22oi_1 _0872_ (.A1(net74),
    .A2(net135),
    .B1(net110),
    .B2(net754),
    .Y(_0376_));
 sky130_fd_sc_hd__nor2_1 _0873_ (.A(net138),
    .B(net755),
    .Y(_0190_));
 sky130_fd_sc_hd__a22oi_1 _0874_ (.A1(net75),
    .A2(net135),
    .B1(net110),
    .B2(net732),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _0875_ (.A(net138),
    .B(net733),
    .Y(_0191_));
 sky130_fd_sc_hd__a22oi_1 _0876_ (.A1(net76),
    .A2(net136),
    .B1(net110),
    .B2(net758),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(net139),
    .B(net759),
    .Y(_0192_));
 sky130_fd_sc_hd__a22oi_1 _0878_ (.A1(net77),
    .A2(net136),
    .B1(net110),
    .B2(net756),
    .Y(_0379_));
 sky130_fd_sc_hd__nor2_1 _0879_ (.A(net139),
    .B(net757),
    .Y(_0193_));
 sky130_fd_sc_hd__a22oi_1 _0880_ (.A1(net78),
    .A2(net136),
    .B1(net111),
    .B2(net714),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _0881_ (.A(net139),
    .B(net715),
    .Y(_0194_));
 sky130_fd_sc_hd__a22oi_1 _0882_ (.A1(net79),
    .A2(net136),
    .B1(net111),
    .B2(net734),
    .Y(_0381_));
 sky130_fd_sc_hd__nor2_1 _0883_ (.A(net139),
    .B(net735),
    .Y(_0195_));
 sky130_fd_sc_hd__a22oi_1 _0884_ (.A1(net80),
    .A2(net136),
    .B1(net111),
    .B2(net710),
    .Y(_0382_));
 sky130_fd_sc_hd__nor2_1 _0885_ (.A(net139),
    .B(net711),
    .Y(_0196_));
 sky130_fd_sc_hd__a22oi_1 _0886_ (.A1(net82),
    .A2(net136),
    .B1(net111),
    .B2(net720),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(net139),
    .B(net721),
    .Y(_0197_));
 sky130_fd_sc_hd__a22oi_1 _0888_ (.A1(net83),
    .A2(net136),
    .B1(net111),
    .B2(net724),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(net139),
    .B(net725),
    .Y(_0198_));
 sky130_fd_sc_hd__a22oi_1 _0890_ (.A1(net84),
    .A2(net136),
    .B1(net111),
    .B2(net742),
    .Y(_0385_));
 sky130_fd_sc_hd__nor2_1 _0891_ (.A(net139),
    .B(net743),
    .Y(_0199_));
 sky130_fd_sc_hd__a22oi_1 _0892_ (.A1(net85),
    .A2(net136),
    .B1(net111),
    .B2(net730),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_1 _0893_ (.A(net139),
    .B(net731),
    .Y(_0200_));
 sky130_fd_sc_hd__a22oi_1 _0894_ (.A1(net86),
    .A2(net136),
    .B1(net111),
    .B2(net728),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(net139),
    .B(net729),
    .Y(_0201_));
 sky130_fd_sc_hd__a22oi_1 _0896_ (.A1(net87),
    .A2(net136),
    .B1(net111),
    .B2(net712),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(net139),
    .B(net713),
    .Y(_0202_));
 sky130_fd_sc_hd__a22oi_1 _0898_ (.A1(net88),
    .A2(net136),
    .B1(net111),
    .B2(net722),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_1 _0899_ (.A(net139),
    .B(net723),
    .Y(_0203_));
 sky130_fd_sc_hd__a22oi_1 _0900_ (.A1(net89),
    .A2(net136),
    .B1(net111),
    .B2(net744),
    .Y(_0390_));
 sky130_fd_sc_hd__nor2_1 _0901_ (.A(net139),
    .B(net745),
    .Y(_0204_));
 sky130_fd_sc_hd__a22oi_1 _0902_ (.A1(net90),
    .A2(net136),
    .B1(net111),
    .B2(net738),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _0903_ (.A(net139),
    .B(net739),
    .Y(_0205_));
 sky130_fd_sc_hd__a22oi_1 _0904_ (.A1(net91),
    .A2(net136),
    .B1(net111),
    .B2(net740),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _0905_ (.A(net139),
    .B(net741),
    .Y(_0206_));
 sky130_fd_sc_hd__a22oi_1 _0906_ (.A1(net93),
    .A2(net136),
    .B1(net111),
    .B2(net716),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_1 _0907_ (.A(net139),
    .B(net717),
    .Y(_0207_));
 sky130_fd_sc_hd__a22oi_1 _0908_ (.A1(net94),
    .A2(_0360_),
    .B1(net111),
    .B2(net718),
    .Y(_0394_));
 sky130_fd_sc_hd__nor2_1 _0909_ (.A(net1),
    .B(net719),
    .Y(_0208_));
 sky130_fd_sc_hd__and4b_1 _0910_ (.A_N(net137),
    .B(net67),
    .C(net692),
    .D(net34),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_4 _0911_ (.A(net137),
    .B(_0407_),
    .Y(_0395_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(net505),
    .A1(net273),
    .S(net103),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0913_ (.A0(net363),
    .A1(net209),
    .S(net103),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(net529),
    .A1(net474),
    .S(net103),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0915_ (.A0(net545),
    .A1(net415),
    .S(net103),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(net381),
    .A1(net339),
    .S(net103),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0917_ (.A0(net395),
    .A1(net336),
    .S(net103),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(net427),
    .A1(net276),
    .S(net103),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0919_ (.A0(net303),
    .A1(net187),
    .S(net103),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(net423),
    .A1(net243),
    .S(net103),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0921_ (.A0(net823),
    .A1(net398),
    .S(net103),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(net349),
    .A1(net157),
    .S(net103),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(net471),
    .A1(net227),
    .S(net103),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(net650),
    .A1(net609),
    .S(net103),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(net676),
    .A1(net636),
    .S(net103),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _0926_ (.A0(net580),
    .A1(net175),
    .S(net103),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(net521),
    .A1(net164),
    .S(net102),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net321),
    .A1(net268),
    .S(net102),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(net572),
    .A1(net501),
    .S(net102),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(net570),
    .A1(net548),
    .S(net102),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(net552),
    .A1(net152),
    .S(net102),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net519),
    .A1(net295),
    .S(net102),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(net435),
    .A1(net145),
    .S(net102),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net417),
    .A1(net184),
    .S(net102),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(net445),
    .A1(net212),
    .S(net102),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(net670),
    .A1(net452),
    .S(net102),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(net623),
    .A1(net541),
    .S(net102),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(net646),
    .A1(net538),
    .S(net102),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(net496),
    .A1(net246),
    .S(net102),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(net387),
    .A1(net204),
    .S(net102),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(net297),
    .A1(net253),
    .S(net102),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(net357),
    .A1(net230),
    .S(net102),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(net638),
    .A1(net465),
    .S(_0395_),
    .X(_0241_));
 sky130_fd_sc_hd__and3b_2 _0944_ (.A_N(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0400_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(net282),
    .A1(net273),
    .S(net108),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(net218),
    .A1(net209),
    .S(net108),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(net564),
    .A1(net474),
    .S(net108),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(net507),
    .A1(net415),
    .S(net108),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(net353),
    .A1(net339),
    .S(net108),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net367),
    .A1(net336),
    .S(net108),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(net329),
    .A1(net276),
    .S(net108),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(net201),
    .A1(net187),
    .S(net108),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(net425),
    .A1(net243),
    .S(net108),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net662),
    .A1(net398),
    .S(net108),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(net166),
    .A1(net157),
    .S(net108),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net458),
    .A1(net227),
    .S(net108),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0957_ (.A0(net652),
    .A1(net609),
    .S(net108),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(net660),
    .A1(net636),
    .S(net108),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(net191),
    .A1(net175),
    .S(net108),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net179),
    .A1(net164),
    .S(net109),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(net584),
    .A1(net268),
    .S(net108),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(net560),
    .A1(net501),
    .S(net109),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(net582),
    .A1(net548),
    .S(net109),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(net170),
    .A1(net152),
    .S(net109),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(net333),
    .A1(net295),
    .S(net109),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(net149),
    .A1(net145),
    .S(net109),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0967_ (.A0(net193),
    .A1(net184),
    .S(net109),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(net240),
    .A1(net212),
    .S(net109),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(net460),
    .A1(net452),
    .S(net109),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(net678),
    .A1(net541),
    .S(net109),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(net826),
    .A1(net538),
    .S(net109),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(net284),
    .A1(net246),
    .S(net109),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(net263),
    .A1(net204),
    .S(net109),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(net290),
    .A1(net253),
    .S(net109),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(net238),
    .A1(net230),
    .S(net109),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(net527),
    .A1(net465),
    .S(net109),
    .X(_0273_));
 sky130_fd_sc_hd__or4_4 _0977_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(net138),
    .D(_0403_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(net273),
    .A1(net854),
    .S(net106),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(net209),
    .A1(net234),
    .S(net106),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(net474),
    .A1(net819),
    .S(net106),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(net415),
    .A1(net837),
    .S(net106),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(net339),
    .A1(net853),
    .S(net106),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _0983_ (.A0(net336),
    .A1(net345),
    .S(net106),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net276),
    .A1(net808),
    .S(net106),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(net187),
    .A1(net199),
    .S(net106),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(net243),
    .A1(net402),
    .S(net106),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(net398),
    .A1(net615),
    .S(net106),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(net157),
    .A1(net177),
    .S(net106),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _0989_ (.A0(net227),
    .A1(net419),
    .S(net106),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(net609),
    .A1(net664),
    .S(net106),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(net636),
    .A1(net668),
    .S(net106),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(net175),
    .A1(net195),
    .S(net107),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(net164),
    .A1(net775),
    .S(net106),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net268),
    .A1(net566),
    .S(net106),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(net501),
    .A1(net509),
    .S(net107),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net548),
    .A1(net816),
    .S(net107),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(net152),
    .A1(net768),
    .S(net107),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(net295),
    .A1(net305),
    .S(net107),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(net145),
    .A1(net147),
    .S(net107),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(net184),
    .A1(net189),
    .S(net107),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(net212),
    .A1(net812),
    .S(net107),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(net452),
    .A1(net454),
    .S(net107),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(net541),
    .A1(net656),
    .S(net107),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(net538),
    .A1(net633),
    .S(net107),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(net246),
    .A1(net806),
    .S(net107),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(net204),
    .A1(net222),
    .S(net107),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(net253),
    .A1(net793),
    .S(net107),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(net230),
    .A1(net327),
    .S(net107),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(net465),
    .A1(net833),
    .S(_0397_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(net301),
    .A1(net273),
    .S(net122),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(net224),
    .A1(net209),
    .S(net122),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(net517),
    .A1(net474),
    .S(net122),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(net478),
    .A1(net415),
    .S(net122),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(net511),
    .A1(net339),
    .S(net122),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(net617),
    .A1(net336),
    .S(net122),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(net313),
    .A1(net276),
    .S(net122),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1017_ (.A0(net197),
    .A1(net187),
    .S(net122),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(net437),
    .A1(net243),
    .S(net122),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(net674),
    .A1(net398),
    .S(net122),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _1020_ (.A0(net787),
    .A1(net157),
    .S(net122),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(net490),
    .A1(net227),
    .S(net122),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(net631),
    .A1(net609),
    .S(net122),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(net672),
    .A1(net636),
    .S(net122),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(net214),
    .A1(net175),
    .S(net122),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1025_ (.A0(net181),
    .A1(net164),
    .S(net121),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1026_ (.A0(net515),
    .A1(net268),
    .S(net121),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(net554),
    .A1(net501),
    .S(net121),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(net574),
    .A1(net548),
    .S(net121),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(net161),
    .A1(net152),
    .S(net121),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(net341),
    .A1(net295),
    .S(net121),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(net172),
    .A1(net145),
    .S(net121),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(net216),
    .A1(net184),
    .S(net121),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1033_ (.A0(net265),
    .A1(net212),
    .S(net121),
    .X(_0329_));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net453),
    .Q(\fifo_in.FIFO[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net542),
    .Q(\fifo_in.FIFO[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net559),
    .Q(\fifo_in.FIFO[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net384),
    .Q(\fifo_in.FIFO[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net260),
    .Q(\fifo_in.FIFO[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net293),
    .Q(\fifo_in.FIFO[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net231),
    .Q(\fifo_in.FIFO[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net526),
    .Q(\fifo_in.FIFO[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net845),
    .Q(\fifo_in.write_addr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1043_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net842),
    .Q(\fifo_in.write_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1044_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net848),
    .Q(\fifo_in.write_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0011_),
    .Q(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0012_),
    .Q(\fifo_in.read_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net850),
    .Q(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net450),
    .Q(\fifo_in.FIFO[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net221),
    .Q(\fifo_in.FIFO[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net589),
    .Q(\fifo_in.FIFO[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net493),
    .Q(\fifo_in.FIFO[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net372),
    .Q(\fifo_in.FIFO[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net362),
    .Q(\fifo_in.FIFO[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net499),
    .Q(\fifo_in.FIFO[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net312),
    .Q(\fifo_in.FIFO[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net279),
    .Q(\fifo_in.FIFO[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net413),
    .Q(\fifo_in.FIFO[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net356),
    .Q(\fifo_in.FIFO[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net483),
    .Q(\fifo_in.FIFO[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net626),
    .Q(\fifo_in.FIFO[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net655),
    .Q(\fifo_in.FIFO[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net597),
    .Q(\fifo_in.FIFO[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net524),
    .Q(\fifo_in.FIFO[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net320),
    .Q(\fifo_in.FIFO[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net532),
    .Q(\fifo_in.FIFO[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net577),
    .Q(\fifo_in.FIFO[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net470),
    .Q(\fifo_in.FIFO[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net468),
    .Q(\fifo_in.FIFO[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net300),
    .Q(\fifo_in.FIFO[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net409),
    .Q(\fifo_in.FIFO[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net390),
    .Q(\fifo_in.FIFO[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net645),
    .Q(\fifo_in.FIFO[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net595),
    .Q(\fifo_in.FIFO[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net622),
    .Q(\fifo_in.FIFO[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net405),
    .Q(\fifo_in.FIFO[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net249),
    .Q(\fifo_in.FIFO[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net318),
    .Q(\fifo_in.FIFO[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net360),
    .Q(\fifo_in.FIFO[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net599),
    .Q(\fifo_in.FIFO[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net411),
    .Q(\fifo_in.FIFO[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net324),
    .Q(\fifo_in.FIFO[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net536),
    .Q(\fifo_in.FIFO[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net422),
    .Q(\fifo_in.FIFO[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net366),
    .Q(\fifo_in.FIFO[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net614),
    .Q(\fifo_in.FIFO[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net514),
    .Q(\fifo_in.FIFO[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net271),
    .Q(\fifo_in.FIFO[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net430),
    .Q(\fifo_in.FIFO[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net620),
    .Q(\fifo_in.FIFO[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net504),
    .Q(\fifo_in.FIFO[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net228),
    .Q(\fifo_in.FIFO[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net649),
    .Q(\fifo_in.FIFO[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net667),
    .Q(\fifo_in.FIFO[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net603),
    .Q(\fifo_in.FIFO[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net487),
    .Q(\fifo_in.FIFO[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net269),
    .Q(\fifo_in.FIFO[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net534),
    .Q(\fifo_in.FIFO[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net685),
    .Q(\fifo_in.FIFO[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net434),
    .Q(\fifo_in.FIFO[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net457),
    .Q(\fifo_in.FIFO[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net258),
    .Q(\fifo_in.FIFO[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net386),
    .Q(\fifo_in.FIFO[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net370),
    .Q(\fifo_in.FIFO[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net601),
    .Q(\fifo_in.FIFO[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net579),
    .Q(\fifo_in.FIFO[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net641),
    .Q(\fifo_in.FIFO[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net401),
    .Q(\fifo_in.FIFO[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net205),
    .Q(\fifo_in.FIFO[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net310),
    .Q(\fifo_in.FIFO[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net326),
    .Q(\fifo_in.FIFO[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net587),
    .Q(\fifo_in.FIFO[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net432),
    .Q(\fifo_in.FIFO[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net233),
    .Q(\fifo_in.FIFO[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net544),
    .Q(\fifo_in.FIFO[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net463),
    .Q(\fifo_in.FIFO[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net376),
    .Q(\fifo_in.FIFO[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net394),
    .Q(\fifo_in.FIFO[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net444),
    .Q(\fifo_in.FIFO[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net440),
    .Q(\fifo_in.FIFO[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net244),
    .Q(\fifo_in.FIFO[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net681),
    .Q(\fifo_in.FIFO[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net380),
    .Q(\fifo_in.FIFO[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net308),
    .Q(\fifo_in.FIFO[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net630),
    .Q(\fifo_in.FIFO[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net683),
    .Q(\fifo_in.FIFO[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net557),
    .Q(\fifo_in.FIFO[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net569),
    .Q(\fifo_in.FIFO[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net332),
    .Q(\fifo_in.FIFO[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net551),
    .Q(\fifo_in.FIFO[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net687),
    .Q(\fifo_in.FIFO[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net477),
    .Q(\fifo_in.FIFO[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net489),
    .Q(\fifo_in.FIFO[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net289),
    .Q(\fifo_in.FIFO[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net281),
    .Q(\fifo_in.FIFO[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net378),
    .Q(\fifo_in.FIFO[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net643),
    .Q(\fifo_in.FIFO[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net605),
    .Q(\fifo_in.FIFO[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net612),
    .Q(\fifo_in.FIFO[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net407),
    .Q(\fifo_in.FIFO[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net251),
    .Q(\fifo_in.FIFO[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net344),
    .Q(\fifo_in.FIFO[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net352),
    .Q(\fifo_in.FIFO[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net628),
    .Q(\fifo_in.FIFO[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net805),
    .Q(\fifo_in.data_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net798),
    .Q(\fifo_in.data_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0112_),
    .Q(\fifo_in.data_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0113_),
    .Q(\fifo_in.data_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net836),
    .Q(\fifo_in.data_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0115_),
    .Q(\fifo_in.data_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0116_),
    .Q(\fifo_in.data_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net767),
    .Q(\fifo_in.data_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net801),
    .Q(\fifo_in.data_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0119_),
    .Q(\fifo_in.data_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net789),
    .Q(\fifo_in.data_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0121_),
    .Q(\fifo_in.data_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0122_),
    .Q(\fifo_in.data_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0123_),
    .Q(\fifo_in.data_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net764),
    .Q(\fifo_in.data_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net777),
    .Q(\fifo_in.data_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0126_),
    .Q(\fifo_in.data_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0127_),
    .Q(\fifo_in.data_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0128_),
    .Q(\fifo_in.data_o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net770),
    .Q(\fifo_in.data_o[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0130_),
    .Q(\fifo_in.data_o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net786),
    .Q(\fifo_in.data_o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net780),
    .Q(\fifo_in.data_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0133_),
    .Q(\fifo_in.data_o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0134_),
    .Q(\fifo_in.data_o[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0135_),
    .Q(\fifo_in.data_o[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0136_),
    .Q(\fifo_in.data_o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0137_),
    .Q(\fifo_in.data_o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net783),
    .Q(\fifo_in.data_o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net795),
    .Q(\fifo_in.data_o[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net792),
    .Q(\fifo_in.data_o[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0141_),
    .Q(\fifo_in.data_o[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net316),
    .Q(\fifo_in.FIFO[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net210),
    .Q(\fifo_in.FIFO[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net495),
    .Q(\fifo_in.FIFO[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net442),
    .Q(\fifo_in.FIFO[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net348),
    .Q(\fifo_in.FIFO[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net337),
    .Q(\fifo_in.FIFO[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net287),
    .Q(\fifo_in.FIFO[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net188),
    .Q(\fifo_in.FIFO[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net392),
    .Q(\fifo_in.FIFO[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net563),
    .Q(\fifo_in.FIFO[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net160),
    .Q(\fifo_in.FIFO[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net448),
    .Q(\fifo_in.FIFO[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net610),
    .Q(\fifo_in.FIFO[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net637),
    .Q(\fifo_in.FIFO[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net176),
    .Q(\fifo_in.FIFO[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net169),
    .Q(\fifo_in.FIFO[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net607),
    .Q(\fifo_in.FIFO[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net502),
    .Q(\fifo_in.FIFO[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net591),
    .Q(\fifo_in.FIFO[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net155),
    .Q(\fifo_in.FIFO[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net296),
    .Q(\fifo_in.FIFO[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net146),
    .Q(\fifo_in.FIFO[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net185),
    .Q(\fifo_in.FIFO[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net237),
    .Q(\fifo_in.FIFO[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net481),
    .Q(\fifo_in.FIFO[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net659),
    .Q(\fifo_in.FIFO[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net593),
    .Q(\fifo_in.FIFO[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net374),
    .Q(\fifo_in.FIFO[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net207),
    .Q(\fifo_in.FIFO[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net256),
    .Q(\fifo_in.FIFO[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net262),
    .Q(\fifo_in.FIFO[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net485),
    .Q(\fifo_in.FIFO[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net761),
    .Q(\fifo_in.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net774),
    .Q(\fifo_in.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net772),
    .Q(\fifo_in.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net143),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0178_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0179_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0180_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0181_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0182_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0183_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0184_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0185_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0186_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0187_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0188_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0189_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0190_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0191_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0192_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0193_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0194_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0195_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0196_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0197_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0198_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0199_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0200_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0201_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0202_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0203_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0204_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0205_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0206_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0207_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0208_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net693),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net506),
    .Q(\fifo_in.FIFO[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net364),
    .Q(\fifo_in.FIFO[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net530),
    .Q(\fifo_in.FIFO[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net546),
    .Q(\fifo_in.FIFO[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net382),
    .Q(\fifo_in.FIFO[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net396),
    .Q(\fifo_in.FIFO[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net428),
    .Q(\fifo_in.FIFO[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net304),
    .Q(\fifo_in.FIFO[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net424),
    .Q(\fifo_in.FIFO[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net399),
    .Q(\fifo_in.FIFO[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net350),
    .Q(\fifo_in.FIFO[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net472),
    .Q(\fifo_in.FIFO[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net651),
    .Q(\fifo_in.FIFO[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net677),
    .Q(\fifo_in.FIFO[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net581),
    .Q(\fifo_in.FIFO[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net522),
    .Q(\fifo_in.FIFO[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net322),
    .Q(\fifo_in.FIFO[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net573),
    .Q(\fifo_in.FIFO[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net571),
    .Q(\fifo_in.FIFO[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net553),
    .Q(\fifo_in.FIFO[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net520),
    .Q(\fifo_in.FIFO[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net436),
    .Q(\fifo_in.FIFO[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net418),
    .Q(\fifo_in.FIFO[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net446),
    .Q(\fifo_in.FIFO[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net671),
    .Q(\fifo_in.FIFO[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net624),
    .Q(\fifo_in.FIFO[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net647),
    .Q(\fifo_in.FIFO[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net497),
    .Q(\fifo_in.FIFO[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net388),
    .Q(\fifo_in.FIFO[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net298),
    .Q(\fifo_in.FIFO[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net358),
    .Q(\fifo_in.FIFO[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net639),
    .Q(\fifo_in.FIFO[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net283),
    .Q(\fifo_in.FIFO[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net219),
    .Q(\fifo_in.FIFO[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net565),
    .Q(\fifo_in.FIFO[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net508),
    .Q(\fifo_in.FIFO[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net354),
    .Q(\fifo_in.FIFO[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net368),
    .Q(\fifo_in.FIFO[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net330),
    .Q(\fifo_in.FIFO[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net202),
    .Q(\fifo_in.FIFO[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net426),
    .Q(\fifo_in.FIFO[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net663),
    .Q(\fifo_in.FIFO[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net167),
    .Q(\fifo_in.FIFO[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net459),
    .Q(\fifo_in.FIFO[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net653),
    .Q(\fifo_in.FIFO[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net661),
    .Q(\fifo_in.FIFO[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net192),
    .Q(\fifo_in.FIFO[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net180),
    .Q(\fifo_in.FIFO[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net585),
    .Q(\fifo_in.FIFO[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net561),
    .Q(\fifo_in.FIFO[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net583),
    .Q(\fifo_in.FIFO[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net171),
    .Q(\fifo_in.FIFO[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net334),
    .Q(\fifo_in.FIFO[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net150),
    .Q(\fifo_in.FIFO[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net194),
    .Q(\fifo_in.FIFO[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net241),
    .Q(\fifo_in.FIFO[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net461),
    .Q(\fifo_in.FIFO[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net679),
    .Q(\fifo_in.FIFO[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net539),
    .Q(\fifo_in.FIFO[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net285),
    .Q(\fifo_in.FIFO[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net264),
    .Q(\fifo_in.FIFO[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net291),
    .Q(\fifo_in.FIFO[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net239),
    .Q(\fifo_in.FIFO[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net528),
    .Q(\fifo_in.FIFO[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net274),
    .Q(\fifo_in.FIFO[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net235),
    .Q(\fifo_in.FIFO[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net475),
    .Q(\fifo_in.FIFO[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net416),
    .Q(\fifo_in.FIFO[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net340),
    .Q(\fifo_in.FIFO[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net346),
    .Q(\fifo_in.FIFO[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net277),
    .Q(\fifo_in.FIFO[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net200),
    .Q(\fifo_in.FIFO[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net403),
    .Q(\fifo_in.FIFO[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net616),
    .Q(\fifo_in.FIFO[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net178),
    .Q(\fifo_in.FIFO[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net420),
    .Q(\fifo_in.FIFO[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net665),
    .Q(\fifo_in.FIFO[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net669),
    .Q(\fifo_in.FIFO[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net196),
    .Q(\fifo_in.FIFO[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net165),
    .Q(\fifo_in.FIFO[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net567),
    .Q(\fifo_in.FIFO[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net510),
    .Q(\fifo_in.FIFO[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net549),
    .Q(\fifo_in.FIFO[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1327_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net153),
    .Q(\fifo_in.FIFO[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net306),
    .Q(\fifo_in.FIFO[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net148),
    .Q(\fifo_in.FIFO[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net190),
    .Q(\fifo_in.FIFO[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net213),
    .Q(\fifo_in.FIFO[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net455),
    .Q(\fifo_in.FIFO[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1333_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net657),
    .Q(\fifo_in.FIFO[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1334_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net634),
    .Q(\fifo_in.FIFO[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1335_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net247),
    .Q(\fifo_in.FIFO[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1336_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net223),
    .Q(\fifo_in.FIFO[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1337_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net254),
    .Q(\fifo_in.FIFO[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1338_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net328),
    .Q(\fifo_in.FIFO[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1339_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net466),
    .Q(\fifo_in.FIFO[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1340_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net302),
    .Q(\fifo_in.FIFO[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1341_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net225),
    .Q(\fifo_in.FIFO[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1342_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net518),
    .Q(\fifo_in.FIFO[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1343_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net479),
    .Q(\fifo_in.FIFO[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1344_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net512),
    .Q(\fifo_in.FIFO[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1345_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net618),
    .Q(\fifo_in.FIFO[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1346_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net314),
    .Q(\fifo_in.FIFO[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1347_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net198),
    .Q(\fifo_in.FIFO[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1348_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net438),
    .Q(\fifo_in.FIFO[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1349_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net675),
    .Q(\fifo_in.FIFO[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1350_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net158),
    .Q(\fifo_in.FIFO[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1351_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net491),
    .Q(\fifo_in.FIFO[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1352_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net632),
    .Q(\fifo_in.FIFO[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1353_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net673),
    .Q(\fifo_in.FIFO[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1354_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net215),
    .Q(\fifo_in.FIFO[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1355_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net182),
    .Q(\fifo_in.FIFO[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1356_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net516),
    .Q(\fifo_in.FIFO[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1357_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net555),
    .Q(\fifo_in.FIFO[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1358_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net575),
    .Q(\fifo_in.FIFO[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1359_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net162),
    .Q(\fifo_in.FIFO[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1360_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net342),
    .Q(\fifo_in.FIFO[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1361_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net173),
    .Q(\fifo_in.FIFO[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1362_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net217),
    .Q(\fifo_in.FIFO[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1363_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net266),
    .Q(\fifo_in.FIFO[0][23] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_8 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_0395_),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(_0419_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_0397_),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(_0396_),
    .X(net108));
 sky130_fd_sc_hd__buf_8 fanout109 (.A(_0396_),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_8 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(_0516_),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(_0418_),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_16 fanout118 (.A(_0417_),
    .X(net118));
 sky130_fd_sc_hd__buf_8 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(_0416_),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(_0401_),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(net799),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(net799),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net129),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net129),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net129),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net851),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(net134),
    .X(net131));
 sky130_fd_sc_hd__buf_8 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(\fifo_in.read_addr[0] ),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(_0360_),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(_0360_),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net1),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net1),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wbs_adr_i[0]),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\fifo_in.FIFO[2][21] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0272_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\fifo_in.FIFO[2][23] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0265_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(wbs_dat_i[8]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 hold104 (.A(net65),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0086_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(wbs_dat_i[27]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 hold107 (.A(net54),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0301_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\fifo_in.FIFO[6][28] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0263_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0042_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\fifo_in.FIFO[4][28] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0106_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(wbs_dat_i[29]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 hold114 (.A(net56),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0303_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\fifo_in.FIFO[3][29] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0171_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\fifo_in.FIFO[5][21] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0067_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(wbs_dat_i[19]),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\fifo_in.FIFO[0][28] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0004_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\fifo_in.FIFO[3][30] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0172_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\fifo_in.FIFO[2][28] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0270_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\fifo_in.FIFO[0][23] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0329_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(wbs_dat_i[16]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 hold129 (.A(net42),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 hold13 (.A(net45),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0062_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\fifo_in.FIFO[5][7] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0053_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(wbs_dat_i[0]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 hold134 (.A(net35),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0274_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(wbs_dat_i[6]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 hold137 (.A(net63),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0280_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\fifo_in.FIFO[6][8] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0293_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0022_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\fifo_in.FIFO[4][22] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0100_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\fifo_in.FIFO[2][0] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0242_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\fifo_in.FIFO[2][27] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0269_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\fifo_in.FIFO[3][6] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0148_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\fifo_in.FIFO[4][21] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\fifo_in.FIFO[3][19] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0099_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\fifo_in.FIFO[2][29] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0271_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\fifo_in.FIFO[0][29] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0005_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(wbs_dat_i[20]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 hold156 (.A(net47),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0162_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\fifo_in.FIFO[7][29] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0239_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0161_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\fifo_in.FIFO[6][21] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0035_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\fifo_in.FIFO[0][0] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0306_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\fifo_in.FIFO[7][7] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0217_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\fifo_in.FIFO[1][20] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0294_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\fifo_in.FIFO[4][11] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0089_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(wbs_dat_i[10]),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\fifo_in.FIFO[5][29] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0075_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\fifo_in.FIFO[6][7] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0021_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\fifo_in.FIFO[0][6] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0312_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\fifo_in.FIFO[3][0] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0142_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\fifo_in.FIFO[6][29] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0043_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 hold18 (.A(net36),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\fifo_in.FIFO[6][16] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0030_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\fifo_in.FIFO[7][16] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0226_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\fifo_in.FIFO[5][1] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0047_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\fifo_in.FIFO[5][30] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0076_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\fifo_in.FIFO[1][30] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0304_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0316_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\fifo_in.FIFO[2][6] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0248_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\fifo_in.FIFO[4][16] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0094_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\fifo_in.FIFO[2][20] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0262_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(wbs_dat_i[5]),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 hold197 (.A(net62),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0147_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(wbs_dat_i[4]),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net2),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\fifo_in.FIFO[3][10] ),
    .X(net159));
 sky130_fd_sc_hd__buf_2 hold200 (.A(net61),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0278_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\fifo_in.FIFO[0][20] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0326_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\fifo_in.FIFO[4][29] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0107_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\fifo_in.FIFO[1][5] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0279_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\fifo_in.FIFO[3][4] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0146_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0152_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\fifo_in.FIFO[7][10] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0220_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\fifo_in.FIFO[4][30] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0108_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\fifo_in.FIFO[2][4] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0246_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\fifo_in.FIFO[6][10] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0024_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\fifo_in.FIFO[7][30] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0240_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\fifo_in.FIFO[0][19] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\fifo_in.FIFO[6][30] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0044_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\fifo_in.FIFO[6][5] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0019_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\fifo_in.FIFO[7][1] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0211_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\fifo_in.FIFO[5][4] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0050_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\fifo_in.FIFO[2][5] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0247_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0325_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\fifo_in.FIFO[5][23] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0069_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\fifo_in.FIFO[6][4] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0018_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\fifo_in.FIFO[3][27] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0169_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\fifo_in.FIFO[4][4] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0082_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\fifo_in.FIFO[4][23] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0101_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(wbs_dat_i[15]),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\fifo_in.FIFO[4][10] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0088_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\fifo_in.FIFO[7][4] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0214_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\fifo_in.FIFO[0][27] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0003_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\fifo_in.FIFO[5][22] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_0068_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\fifo_in.FIFO[7][28] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0238_),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 hold25 (.A(net41),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\fifo_in.FIFO[6][23] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0037_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\fifo_in.FIFO[3][8] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0150_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\fifo_in.FIFO[4][5] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0083_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\fifo_in.FIFO[7][5] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0215_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(wbs_dat_i[9]),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 hold259 (.A(net66),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0289_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0219_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\fifo_in.FIFO[5][27] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0073_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\fifo_in.FIFO[1][8] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0282_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\fifo_in.FIFO[6][27] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0041_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\fifo_in.FIFO[4][27] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0105_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\fifo_in.FIFO[6][22] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fifo_in.FIFO[2][10] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0036_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\fifo_in.FIFO[5][0] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0046_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\fifo_in.FIFO[6][9] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0023_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(wbs_dat_i[3]),
    .X(net414));
 sky130_fd_sc_hd__buf_2 hold276 (.A(net60),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0277_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\fifo_in.FIFO[7][22] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0232_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0252_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\fifo_in.FIFO[1][11] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0285_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\fifo_in.FIFO[5][3] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0049_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\fifo_in.FIFO[7][8] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0218_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\fifo_in.FIFO[2][8] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0250_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\fifo_in.FIFO[7][6] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0216_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fifo_in.FIFO[3][15] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\fifo_in.FIFO[5][8] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0054_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\fifo_in.FIFO[4][0] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0078_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\fifo_in.FIFO[5][19] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0065_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\fifo_in.FIFO[7][21] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0231_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\fifo_in.FIFO[0][8] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0314_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0361_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0157_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\fifo_in.FIFO[4][7] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0085_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\fifo_in.FIFO[3][3] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0145_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\fifo_in.FIFO[4][6] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0084_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\fifo_in.FIFO[7][23] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0233_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\fifo_in.FIFO[3][11] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0153_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\fifo_in.FIFO[2][19] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\fifo_in.FIFO[6][0] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0014_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(wbs_dat_i[24]),
    .X(net451));
 sky130_fd_sc_hd__buf_2 hold313 (.A(net51),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0000_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\fifo_in.FIFO[1][24] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0298_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\fifo_in.FIFO[5][20] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0066_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\fifo_in.FIFO[2][11] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0261_),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0253_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\fifo_in.FIFO[2][24] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0266_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\fifo_in.FIFO[4][3] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0081_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(wbs_dat_i[31]),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_2 hold326 (.A(net59),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0305_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\fifo_in.FIFO[6][20] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0034_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fifo_in.FIFO[0][21] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\fifo_in.FIFO[6][19] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0033_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\fifo_in.FIFO[7][11] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0221_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(wbs_dat_i[2]),
    .X(net473));
 sky130_fd_sc_hd__buf_2 hold335 (.A(net57),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0276_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\fifo_in.FIFO[4][19] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0097_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\fifo_in.FIFO[0][3] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0327_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0309_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\fifo_in.FIFO[3][24] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0166_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\fifo_in.FIFO[6][11] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0025_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\fifo_in.FIFO[3][31] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0173_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\fifo_in.FIFO[5][15] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0061_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\fifo_in.FIFO[4][20] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(wbs_dat_i[14]),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0098_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\fifo_in.FIFO[0][11] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0317_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\fifo_in.FIFO[6][3] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0017_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\fifo_in.FIFO[3][2] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0144_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\fifo_in.FIFO[7][27] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0237_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\fifo_in.FIFO[6][6] ),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_2 hold36 (.A(net40),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0020_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(wbs_dat_i[17]),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_2 hold362 (.A(net43),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0159_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\fifo_in.FIFO[5][10] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_0056_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\fifo_in.FIFO[7][0] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_0210_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\fifo_in.FIFO[2][3] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0245_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0156_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\fifo_in.FIFO[1][17] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_0291_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\fifo_in.FIFO[0][4] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_0310_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\fifo_in.FIFO[5][6] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_0052_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\fifo_in.FIFO[0][16] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_0322_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\fifo_in.FIFO[0][2] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_0308_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fifo_in.FIFO[1][10] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\fifo_in.FIFO[7][20] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0230_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\fifo_in.FIFO[7][15] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0225_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\fifo_in.FIFO[6][15] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0029_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\fifo_in.FIFO[0][31] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_0007_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\fifo_in.FIFO[2][31] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_0273_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0284_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\fifo_in.FIFO[7][2] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0212_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\fifo_in.FIFO[6][17] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0031_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\fifo_in.FIFO[5][17] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0063_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\fifo_in.FIFO[5][2] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_0048_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(wbs_dat_i[26]),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_2 hold399 (.A(net53),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0177_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\fifo_in.FIFO[2][15] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0268_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(wbs_dat_i[25]),
    .X(net540));
 sky130_fd_sc_hd__buf_2 hold402 (.A(net52),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_0001_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\fifo_in.FIFO[4][2] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0080_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\fifo_in.FIFO[7][3] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0213_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(wbs_dat_i[18]),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_2 hold409 (.A(net44),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0257_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0292_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\fifo_in.FIFO[4][17] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0095_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\fifo_in.FIFO[7][19] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0229_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\fifo_in.FIFO[0][17] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0323_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\fifo_in.FIFO[4][14] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0092_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\fifo_in.FIFO[0][26] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\fifo_in.FIFO[0][15] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0002_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\fifo_in.FIFO[2][17] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0259_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\fifo_in.FIFO[3][9] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0151_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\fifo_in.FIFO[2][2] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0244_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\fifo_in.FIFO[1][16] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0290_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\fifo_in.FIFO[4][15] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0321_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0093_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\fifo_in.FIFO[7][18] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0228_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\fifo_in.FIFO[7][17] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0227_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\fifo_in.FIFO[0][18] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0324_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\fifo_in.FIFO[6][18] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0032_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\fifo_in.FIFO[5][25] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(wbs_dat_i[22]),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0071_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\fifo_in.FIFO[7][14] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0224_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\fifo_in.FIFO[2][18] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0260_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\fifo_in.FIFO[2][16] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0258_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\fifo_in.FIFO[5][31] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0077_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\fifo_in.FIFO[6][2] ),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 hold45 (.A(net49),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0016_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\fifo_in.FIFO[3][18] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0160_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\fifo_in.FIFO[3][26] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0168_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\fifo_in.FIFO[6][25] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0039_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\fifo_in.FIFO[6][14] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0028_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\fifo_in.FIFO[6][31] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0164_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0045_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\fifo_in.FIFO[5][24] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0070_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\fifo_in.FIFO[5][14] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0060_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\fifo_in.FIFO[4][25] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0103_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\fifo_in.FIFO[3][16] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0158_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(wbs_dat_i[12]),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(wbs_dat_i[7]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 hold470 (.A(net38),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0154_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\fifo_in.FIFO[4][26] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0104_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\fifo_in.FIFO[5][5] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0051_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\fifo_in.FIFO[1][9] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0283_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\fifo_in.FIFO[0][5] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0311_),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 hold48 (.A(net64),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\fifo_in.FIFO[5][9] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0055_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\fifo_in.FIFO[6][26] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0040_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\fifo_in.FIFO[7][25] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0235_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\fifo_in.FIFO[6][12] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0026_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\fifo_in.FIFO[4][31] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0109_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0149_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\fifo_in.FIFO[4][12] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0090_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\fifo_in.FIFO[0][12] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0318_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\fifo_in.FIFO[1][26] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0300_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(wbs_dat_i[13]),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_2 hold497 (.A(net39),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0155_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\fifo_in.FIFO[7][31] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(wbs_dat_i[21]),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\fifo_in.FIFO[1][22] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0241_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\fifo_in.FIFO[5][26] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0072_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\fifo_in.FIFO[4][24] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0102_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\fifo_in.FIFO[6][24] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0038_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\fifo_in.FIFO[7][26] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0236_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\fifo_in.FIFO[5][12] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0296_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0058_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\fifo_in.FIFO[7][12] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0222_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\fifo_in.FIFO[2][12] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0254_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\fifo_in.FIFO[6][13] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0027_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\fifo_in.FIFO[1][25] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0299_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\fifo_in.FIFO[3][25] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\fifo_in.FIFO[2][14] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0167_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\fifo_in.FIFO[2][13] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0255_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\fifo_in.FIFO[2][9] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0251_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\fifo_in.FIFO[1][12] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0286_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\fifo_in.FIFO[5][13] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0059_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\fifo_in.FIFO[1][13] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0256_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0287_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\fifo_in.FIFO[7][24] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0234_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\fifo_in.FIFO[0][13] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0319_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\fifo_in.FIFO[0][9] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0315_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\fifo_in.FIFO[7][13] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0223_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\fifo_in.FIFO[2][25] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\fifo_in.FIFO[2][22] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0267_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\fifo_in.FIFO[4][9] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0087_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\fifo_in.FIFO[4][13] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0091_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\fifo_in.FIFO[5][18] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0064_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\fifo_in.FIFO[4][18] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0096_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(wbs_adr_i[6]),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0264_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net30),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0354_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0358_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0359_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0209_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(wbs_adr_i[22]),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(net16),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0349_),
    .X(net696));
 sky130_fd_sc_hd__buf_1 hold558 (.A(_0353_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0363_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\fifo_in.FIFO[1][14] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0367_),
    .X(net699));
 sky130_fd_sc_hd__buf_1 hold561 (.A(net860),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0368_),
    .X(net701));
 sky130_fd_sc_hd__buf_1 hold563 (.A(net862),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0366_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\fifo_in.data_o[1] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0364_),
    .X(net705));
 sky130_fd_sc_hd__buf_1 hold567 (.A(net857),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0365_),
    .X(net707));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold569 (.A(\fifo_in.data_o[6] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0288_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0369_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\fifo_in.data_o[19] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0382_),
    .X(net711));
 sky130_fd_sc_hd__buf_1 hold573 (.A(net863),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0388_),
    .X(net713));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold575 (.A(\fifo_in.data_o[17] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0380_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\fifo_in.data_o[30] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0393_),
    .X(net717));
 sky130_fd_sc_hd__buf_1 hold579 (.A(net861),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\fifo_in.FIFO[0][7] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0394_),
    .X(net719));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold581 (.A(\fifo_in.data_o[20] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0383_),
    .X(net721));
 sky130_fd_sc_hd__buf_1 hold583 (.A(net856),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0389_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\fifo_in.data_o[21] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0384_),
    .X(net725));
 sky130_fd_sc_hd__buf_1 hold587 (.A(net858),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0372_),
    .X(net727));
 sky130_fd_sc_hd__buf_1 hold589 (.A(net859),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0313_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0387_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\fifo_in.data_o[23] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0386_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\fifo_in.data_o[14] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0377_),
    .X(net733));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold595 (.A(\fifo_in.data_o[18] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0381_),
    .X(net735));
 sky130_fd_sc_hd__buf_1 hold597 (.A(net855),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0375_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\fifo_in.data_o[28] ),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_2 hold6 (.A(net48),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\fifo_in.FIFO[1][7] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0391_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\fifo_in.data_o[29] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0392_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\fifo_in.data_o[22] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0385_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\fifo_in.data_o[27] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0390_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\fifo_in.data_o[8] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0371_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\fifo_in.data_o[11] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0281_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0374_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\fifo_in.data_o[7] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0370_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\fifo_in.data_o[10] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0373_),
    .X(net753));
 sky130_fd_sc_hd__buf_1 hold615 (.A(net864),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0376_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\fifo_in.data_o[16] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0379_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\fifo_in.data_o[15] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\fifo_in.FIFO[2][7] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0378_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\fifo_in.count[0] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0174_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\fifo_in.FIFO[3][14] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0464_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_0124_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\fifo_in.FIFO[3][7] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_0443_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0117_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\fifo_in.FIFO[1][19] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0249_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0479_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_0129_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\fifo_in.count[2] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_0176_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\fifo_in.count[1] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_0175_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\fifo_in.FIFO[1][15] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_0467_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0125_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\fifo_in.FIFO[3][22] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(wbs_dat_i[28]),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0488_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_0132_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\fifo_in.FIFO[5][28] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_0506_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0138_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\fifo_in.FIFO[3][21] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0485_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_0131_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\fifo_in.FIFO[0][10] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_0452_),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 hold65 (.A(net55),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0120_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\fifo_in.FIFO[0][30] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0512_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(_0140_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\fifo_in.FIFO[1][29] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(_0509_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0139_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\fifo_in.FIFO[3][1] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_0425_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0111_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0074_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 hold660 (.A(net849),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_0446_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_0118_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\fifo_in.FIFO[5][11] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0455_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\fifo_in.data_o[0] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0110_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\fifo_in.FIFO[1][27] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0503_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\fifo_in.FIFO[1][6] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\fifo_in.FIFO[3][28] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_0440_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\fifo_in.FIFO[5][16] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0470_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\fifo_in.FIFO[1][23] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0491_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\fifo_in.FIFO[3][20] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_0482_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\fifo_in.FIFO[1][18] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_0476_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\fifo_in.FIFO[3][12] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0170_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\fifo_in.FIFO[1][2] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_0428_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\fifo_in.FIFO[3][17] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_0473_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\fifo_in.FIFO[7][9] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\fifo_in.FIFO[0][24] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_0494_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\fifo_in.FIFO[2][26] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_0499_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0500_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(wbs_dat_i[1]),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\fifo_in.FIFO[3][5] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_0436_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\fifo_in.FIFO[3][13] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_0461_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\fifo_in.FIFO[1][31] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_0515_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\fifo_in.data_o[4] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_0114_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\fifo_in.FIFO[1][3] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_0431_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0163_),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 hold70 (.A(net46),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\fifo_in.FIFO[0][25] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_0497_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\fifo_in.write_addr[1] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_0009_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(wbs_we_i),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_0403_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0008_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\fifo_in.write_addr[2] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_0407_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_0010_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0143_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\fifo_in.read_addr[2] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_0013_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\fifo_in.read_addr[1] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\fifo_in.FIFO[4][8] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\fifo_in.FIFO[1][4] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\fifo_in.FIFO[1][0] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\fifo_in.data_o[12] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\fifo_in.data_o[26] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\fifo_in.data_o[2] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\fifo_in.data_o[9] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(wbs_dat_i[23]),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\fifo_in.data_o[24] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\fifo_in.data_o[5] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\fifo_in.data_o[31] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\fifo_in.data_o[3] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\fifo_in.data_o[25] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\fifo_in.data_o[13] ),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 hold73 (.A(net50),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0297_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\fifo_in.FIFO[0][14] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0320_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\fifo_in.FIFO[0][22] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0328_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\fifo_in.FIFO[2][1] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\fifo_in.FIFO[1][21] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0243_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\fifo_in.FIFO[6][1] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0015_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\fifo_in.FIFO[1][28] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0302_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\fifo_in.FIFO[0][1] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0307_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(wbs_dat_i[11]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 hold88 (.A(net37),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0057_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0295_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(wbs_dat_i[30]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 hold91 (.A(net58),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0006_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\fifo_in.FIFO[4][1] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0079_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\fifo_in.FIFO[1][1] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0275_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\fifo_in.FIFO[3][23] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0165_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\fifo_in.FIFO[2][30] ),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(wbs_adr_i[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wbs_adr_i[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(wbs_adr_i[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(wbs_adr_i[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(wbs_adr_i[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(wbs_adr_i[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net694),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(wbs_adr_i[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(wbs_adr_i[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(wbs_adr_i[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net140),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(wbs_adr_i[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(wbs_adr_i[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(wbs_adr_i[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(wbs_adr_i[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(wbs_adr_i[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(wbs_adr_i[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(wbs_adr_i[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(wbs_adr_i[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(wbs_adr_i[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(wbs_adr_i[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(wbs_adr_i[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net688),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(wbs_adr_i[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(wbs_adr_i[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(wbs_adr_i[9]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(wbs_cyc_i),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(net272),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(net156),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net226),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net608),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(net635),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(wbs_adr_i[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net174),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net163),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net267),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net500),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net547),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net151),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(net208),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net294),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net144),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(net183),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(wbs_adr_i[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net211),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(net451),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net540),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(net537),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net245),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(net203),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(net252),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(net473),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(net229),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(net464),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(wbs_adr_i[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(net414),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(net338),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(net335),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(net275),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net186),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(net242),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(net397),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(wbs_stb_i),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(net843),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(wbs_adr_i[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(wbs_adr_i[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(wbs_adr_i[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__clkbuf_2 wire112 (.A(net698),
    .X(net112));
endmodule

