magic
tech sky130A
magscale 1 2
timestamp 1725547226
<< nwell >>
rect 1066 27461 58918 27782
rect 1066 26373 58918 26939
rect 1066 25285 58918 25851
rect 1066 24197 58918 24763
rect 1066 23109 58918 23675
rect 1066 22021 58918 22587
rect 1066 20933 58918 21499
rect 1066 19845 58918 20411
rect 1066 18757 58918 19323
rect 1066 17669 58918 18235
rect 1066 16581 58918 17147
rect 1066 15493 58918 16059
rect 1066 14405 58918 14971
rect 1066 13317 58918 13883
rect 1066 12229 58918 12795
rect 1066 11141 58918 11707
rect 1066 10053 58918 10619
rect 1066 8965 58918 9531
rect 1066 7877 58918 8443
rect 1066 6789 58918 7355
rect 1066 5701 58918 6267
rect 1066 4613 58918 5179
rect 1066 3525 58918 4091
rect 1066 2437 58918 3003
<< obsli1 >>
rect 1104 2159 58880 27761
<< obsm1 >>
rect 1104 2048 59040 27792
<< metal2 >>
rect 1398 0 1454 800
rect 2226 0 2282 800
rect 3054 0 3110 800
rect 3882 0 3938 800
rect 4710 0 4766 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 8022 0 8078 800
rect 8850 0 8906 800
rect 9678 0 9734 800
rect 10506 0 10562 800
rect 11334 0 11390 800
rect 12162 0 12218 800
rect 12990 0 13046 800
rect 13818 0 13874 800
rect 14646 0 14702 800
rect 15474 0 15530 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19614 0 19670 800
rect 20442 0 20498 800
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 57702 0 57758 800
rect 58530 0 58586 800
<< obsm2 >>
rect 1398 856 59034 27781
rect 1510 734 2170 856
rect 2338 734 2998 856
rect 3166 734 3826 856
rect 3994 734 4654 856
rect 4822 734 5482 856
rect 5650 734 6310 856
rect 6478 734 7138 856
rect 7306 734 7966 856
rect 8134 734 8794 856
rect 8962 734 9622 856
rect 9790 734 10450 856
rect 10618 734 11278 856
rect 11446 734 12106 856
rect 12274 734 12934 856
rect 13102 734 13762 856
rect 13930 734 14590 856
rect 14758 734 15418 856
rect 15586 734 16246 856
rect 16414 734 17074 856
rect 17242 734 17902 856
rect 18070 734 18730 856
rect 18898 734 19558 856
rect 19726 734 20386 856
rect 20554 734 21214 856
rect 21382 734 22042 856
rect 22210 734 22870 856
rect 23038 734 23698 856
rect 23866 734 24526 856
rect 24694 734 25354 856
rect 25522 734 26182 856
rect 26350 734 27010 856
rect 27178 734 27838 856
rect 28006 734 28666 856
rect 28834 734 29494 856
rect 29662 734 30322 856
rect 30490 734 31150 856
rect 31318 734 31978 856
rect 32146 734 32806 856
rect 32974 734 33634 856
rect 33802 734 34462 856
rect 34630 734 35290 856
rect 35458 734 36118 856
rect 36286 734 36946 856
rect 37114 734 37774 856
rect 37942 734 38602 856
rect 38770 734 39430 856
rect 39598 734 40258 856
rect 40426 734 41086 856
rect 41254 734 41914 856
rect 42082 734 42742 856
rect 42910 734 43570 856
rect 43738 734 44398 856
rect 44566 734 45226 856
rect 45394 734 46054 856
rect 46222 734 46882 856
rect 47050 734 47710 856
rect 47878 734 48538 856
rect 48706 734 49366 856
rect 49534 734 50194 856
rect 50362 734 51022 856
rect 51190 734 51850 856
rect 52018 734 52678 856
rect 52846 734 53506 856
rect 53674 734 54334 856
rect 54502 734 55162 856
rect 55330 734 55990 856
rect 56158 734 56818 856
rect 56986 734 57646 856
rect 57814 734 58474 856
rect 58642 734 59034 856
<< obsm3 >>
rect 1393 2143 59038 27777
<< metal4 >>
rect 8166 2128 8486 27792
rect 15388 2128 15708 27792
rect 22610 2128 22930 27792
rect 29832 2128 30152 27792
rect 37054 2128 37374 27792
rect 44276 2128 44596 27792
rect 51498 2128 51818 27792
rect 58720 2128 59040 27792
<< obsm4 >>
rect 6683 3979 8086 20773
rect 8566 3979 15308 20773
rect 15788 3979 22530 20773
rect 23010 3979 29752 20773
rect 30232 3979 36974 20773
rect 37454 3979 42445 20773
<< labels >>
rlabel metal4 s 8166 2128 8486 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 22610 2128 22930 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 37054 2128 37374 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 51498 2128 51818 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 15388 2128 15708 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 29832 2128 30152 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 44276 2128 44596 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 58720 2128 59040 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal2 s 1398 0 1454 800 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wb_rst_i
port 4 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 5 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_cyc_i
port 6 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[0]
port 7 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[10]
port 8 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[11]
port 9 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[12]
port 10 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[13]
port 11 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_i[14]
port 12 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[15]
port 13 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[16]
port 14 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[17]
port 15 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[18]
port 16 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[19]
port 17 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_i[1]
port 18 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[20]
port 19 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[21]
port 20 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[22]
port 21 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[23]
port 22 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_i[24]
port 23 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_i[25]
port 24 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[26]
port 25 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_i[27]
port 26 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[28]
port 27 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[29]
port 28 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[2]
port 29 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[30]
port 30 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_i[31]
port 31 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[3]
port 32 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[4]
port 33 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[5]
port 34 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[6]
port 35 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[7]
port 36 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[8]
port 37 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[9]
port 38 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[0]
port 39 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[10]
port 40 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[11]
port 41 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[12]
port 42 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[13]
port 43 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[14]
port 44 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[15]
port 45 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_o[16]
port 46 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[17]
port 47 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[18]
port 48 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[19]
port 49 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[1]
port 50 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[20]
port 51 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[21]
port 52 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[22]
port 53 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[23]
port 54 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[24]
port 55 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[25]
port 56 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_o[26]
port 57 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[27]
port 58 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_o[28]
port 59 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[29]
port 60 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[2]
port 61 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[30]
port 62 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_o[31]
port 63 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[3]
port 64 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[4]
port 65 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[5]
port 66 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[6]
port 67 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[7]
port 68 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_o[8]
port 69 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[9]
port 70 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_stb_i
port 71 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_we_i
port 72 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3833726
string GDS_FILE /home/jelmer/Documents/stage/efabless/caravel_user_project/openlane/wishbone_nn/runs/24_09_05_16_39/results/signoff/wishbone_nn.magic.gds
string GDS_START 369158
<< end >>

