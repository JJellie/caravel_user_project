// This is the unpowered netlist.
module wishbone_nn (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_dat_i,
    wbs_dat_o);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \fifo_in.FIFO[0][0] ;
 wire \fifo_in.FIFO[0][10] ;
 wire \fifo_in.FIFO[0][11] ;
 wire \fifo_in.FIFO[0][12] ;
 wire \fifo_in.FIFO[0][13] ;
 wire \fifo_in.FIFO[0][14] ;
 wire \fifo_in.FIFO[0][15] ;
 wire \fifo_in.FIFO[0][16] ;
 wire \fifo_in.FIFO[0][17] ;
 wire \fifo_in.FIFO[0][18] ;
 wire \fifo_in.FIFO[0][19] ;
 wire \fifo_in.FIFO[0][1] ;
 wire \fifo_in.FIFO[0][20] ;
 wire \fifo_in.FIFO[0][21] ;
 wire \fifo_in.FIFO[0][22] ;
 wire \fifo_in.FIFO[0][23] ;
 wire \fifo_in.FIFO[0][24] ;
 wire \fifo_in.FIFO[0][25] ;
 wire \fifo_in.FIFO[0][26] ;
 wire \fifo_in.FIFO[0][27] ;
 wire \fifo_in.FIFO[0][28] ;
 wire \fifo_in.FIFO[0][29] ;
 wire \fifo_in.FIFO[0][2] ;
 wire \fifo_in.FIFO[0][30] ;
 wire \fifo_in.FIFO[0][31] ;
 wire \fifo_in.FIFO[0][3] ;
 wire \fifo_in.FIFO[0][4] ;
 wire \fifo_in.FIFO[0][5] ;
 wire \fifo_in.FIFO[0][6] ;
 wire \fifo_in.FIFO[0][7] ;
 wire \fifo_in.FIFO[0][8] ;
 wire \fifo_in.FIFO[0][9] ;
 wire \fifo_in.FIFO[1][0] ;
 wire \fifo_in.FIFO[1][10] ;
 wire \fifo_in.FIFO[1][11] ;
 wire \fifo_in.FIFO[1][12] ;
 wire \fifo_in.FIFO[1][13] ;
 wire \fifo_in.FIFO[1][14] ;
 wire \fifo_in.FIFO[1][15] ;
 wire \fifo_in.FIFO[1][16] ;
 wire \fifo_in.FIFO[1][17] ;
 wire \fifo_in.FIFO[1][18] ;
 wire \fifo_in.FIFO[1][19] ;
 wire \fifo_in.FIFO[1][1] ;
 wire \fifo_in.FIFO[1][20] ;
 wire \fifo_in.FIFO[1][21] ;
 wire \fifo_in.FIFO[1][22] ;
 wire \fifo_in.FIFO[1][23] ;
 wire \fifo_in.FIFO[1][24] ;
 wire \fifo_in.FIFO[1][25] ;
 wire \fifo_in.FIFO[1][26] ;
 wire \fifo_in.FIFO[1][27] ;
 wire \fifo_in.FIFO[1][28] ;
 wire \fifo_in.FIFO[1][29] ;
 wire \fifo_in.FIFO[1][2] ;
 wire \fifo_in.FIFO[1][30] ;
 wire \fifo_in.FIFO[1][31] ;
 wire \fifo_in.FIFO[1][3] ;
 wire \fifo_in.FIFO[1][4] ;
 wire \fifo_in.FIFO[1][5] ;
 wire \fifo_in.FIFO[1][6] ;
 wire \fifo_in.FIFO[1][7] ;
 wire \fifo_in.FIFO[1][8] ;
 wire \fifo_in.FIFO[1][9] ;
 wire \fifo_in.FIFO[2][0] ;
 wire \fifo_in.FIFO[2][10] ;
 wire \fifo_in.FIFO[2][11] ;
 wire \fifo_in.FIFO[2][12] ;
 wire \fifo_in.FIFO[2][13] ;
 wire \fifo_in.FIFO[2][14] ;
 wire \fifo_in.FIFO[2][15] ;
 wire \fifo_in.FIFO[2][16] ;
 wire \fifo_in.FIFO[2][17] ;
 wire \fifo_in.FIFO[2][18] ;
 wire \fifo_in.FIFO[2][19] ;
 wire \fifo_in.FIFO[2][1] ;
 wire \fifo_in.FIFO[2][20] ;
 wire \fifo_in.FIFO[2][21] ;
 wire \fifo_in.FIFO[2][22] ;
 wire \fifo_in.FIFO[2][23] ;
 wire \fifo_in.FIFO[2][24] ;
 wire \fifo_in.FIFO[2][25] ;
 wire \fifo_in.FIFO[2][26] ;
 wire \fifo_in.FIFO[2][27] ;
 wire \fifo_in.FIFO[2][28] ;
 wire \fifo_in.FIFO[2][29] ;
 wire \fifo_in.FIFO[2][2] ;
 wire \fifo_in.FIFO[2][30] ;
 wire \fifo_in.FIFO[2][31] ;
 wire \fifo_in.FIFO[2][3] ;
 wire \fifo_in.FIFO[2][4] ;
 wire \fifo_in.FIFO[2][5] ;
 wire \fifo_in.FIFO[2][6] ;
 wire \fifo_in.FIFO[2][7] ;
 wire \fifo_in.FIFO[2][8] ;
 wire \fifo_in.FIFO[2][9] ;
 wire \fifo_in.FIFO[3][0] ;
 wire \fifo_in.FIFO[3][10] ;
 wire \fifo_in.FIFO[3][11] ;
 wire \fifo_in.FIFO[3][12] ;
 wire \fifo_in.FIFO[3][13] ;
 wire \fifo_in.FIFO[3][14] ;
 wire \fifo_in.FIFO[3][15] ;
 wire \fifo_in.FIFO[3][16] ;
 wire \fifo_in.FIFO[3][17] ;
 wire \fifo_in.FIFO[3][18] ;
 wire \fifo_in.FIFO[3][19] ;
 wire \fifo_in.FIFO[3][1] ;
 wire \fifo_in.FIFO[3][20] ;
 wire \fifo_in.FIFO[3][21] ;
 wire \fifo_in.FIFO[3][22] ;
 wire \fifo_in.FIFO[3][23] ;
 wire \fifo_in.FIFO[3][24] ;
 wire \fifo_in.FIFO[3][25] ;
 wire \fifo_in.FIFO[3][26] ;
 wire \fifo_in.FIFO[3][27] ;
 wire \fifo_in.FIFO[3][28] ;
 wire \fifo_in.FIFO[3][29] ;
 wire \fifo_in.FIFO[3][2] ;
 wire \fifo_in.FIFO[3][30] ;
 wire \fifo_in.FIFO[3][31] ;
 wire \fifo_in.FIFO[3][3] ;
 wire \fifo_in.FIFO[3][4] ;
 wire \fifo_in.FIFO[3][5] ;
 wire \fifo_in.FIFO[3][6] ;
 wire \fifo_in.FIFO[3][7] ;
 wire \fifo_in.FIFO[3][8] ;
 wire \fifo_in.FIFO[3][9] ;
 wire \fifo_in.FIFO[4][0] ;
 wire \fifo_in.FIFO[4][10] ;
 wire \fifo_in.FIFO[4][11] ;
 wire \fifo_in.FIFO[4][12] ;
 wire \fifo_in.FIFO[4][13] ;
 wire \fifo_in.FIFO[4][14] ;
 wire \fifo_in.FIFO[4][15] ;
 wire \fifo_in.FIFO[4][16] ;
 wire \fifo_in.FIFO[4][17] ;
 wire \fifo_in.FIFO[4][18] ;
 wire \fifo_in.FIFO[4][19] ;
 wire \fifo_in.FIFO[4][1] ;
 wire \fifo_in.FIFO[4][20] ;
 wire \fifo_in.FIFO[4][21] ;
 wire \fifo_in.FIFO[4][22] ;
 wire \fifo_in.FIFO[4][23] ;
 wire \fifo_in.FIFO[4][24] ;
 wire \fifo_in.FIFO[4][25] ;
 wire \fifo_in.FIFO[4][26] ;
 wire \fifo_in.FIFO[4][27] ;
 wire \fifo_in.FIFO[4][28] ;
 wire \fifo_in.FIFO[4][29] ;
 wire \fifo_in.FIFO[4][2] ;
 wire \fifo_in.FIFO[4][30] ;
 wire \fifo_in.FIFO[4][31] ;
 wire \fifo_in.FIFO[4][3] ;
 wire \fifo_in.FIFO[4][4] ;
 wire \fifo_in.FIFO[4][5] ;
 wire \fifo_in.FIFO[4][6] ;
 wire \fifo_in.FIFO[4][7] ;
 wire \fifo_in.FIFO[4][8] ;
 wire \fifo_in.FIFO[4][9] ;
 wire \fifo_in.FIFO[5][0] ;
 wire \fifo_in.FIFO[5][10] ;
 wire \fifo_in.FIFO[5][11] ;
 wire \fifo_in.FIFO[5][12] ;
 wire \fifo_in.FIFO[5][13] ;
 wire \fifo_in.FIFO[5][14] ;
 wire \fifo_in.FIFO[5][15] ;
 wire \fifo_in.FIFO[5][16] ;
 wire \fifo_in.FIFO[5][17] ;
 wire \fifo_in.FIFO[5][18] ;
 wire \fifo_in.FIFO[5][19] ;
 wire \fifo_in.FIFO[5][1] ;
 wire \fifo_in.FIFO[5][20] ;
 wire \fifo_in.FIFO[5][21] ;
 wire \fifo_in.FIFO[5][22] ;
 wire \fifo_in.FIFO[5][23] ;
 wire \fifo_in.FIFO[5][24] ;
 wire \fifo_in.FIFO[5][25] ;
 wire \fifo_in.FIFO[5][26] ;
 wire \fifo_in.FIFO[5][27] ;
 wire \fifo_in.FIFO[5][28] ;
 wire \fifo_in.FIFO[5][29] ;
 wire \fifo_in.FIFO[5][2] ;
 wire \fifo_in.FIFO[5][30] ;
 wire \fifo_in.FIFO[5][31] ;
 wire \fifo_in.FIFO[5][3] ;
 wire \fifo_in.FIFO[5][4] ;
 wire \fifo_in.FIFO[5][5] ;
 wire \fifo_in.FIFO[5][6] ;
 wire \fifo_in.FIFO[5][7] ;
 wire \fifo_in.FIFO[5][8] ;
 wire \fifo_in.FIFO[5][9] ;
 wire \fifo_in.FIFO[6][0] ;
 wire \fifo_in.FIFO[6][10] ;
 wire \fifo_in.FIFO[6][11] ;
 wire \fifo_in.FIFO[6][12] ;
 wire \fifo_in.FIFO[6][13] ;
 wire \fifo_in.FIFO[6][14] ;
 wire \fifo_in.FIFO[6][15] ;
 wire \fifo_in.FIFO[6][16] ;
 wire \fifo_in.FIFO[6][17] ;
 wire \fifo_in.FIFO[6][18] ;
 wire \fifo_in.FIFO[6][19] ;
 wire \fifo_in.FIFO[6][1] ;
 wire \fifo_in.FIFO[6][20] ;
 wire \fifo_in.FIFO[6][21] ;
 wire \fifo_in.FIFO[6][22] ;
 wire \fifo_in.FIFO[6][23] ;
 wire \fifo_in.FIFO[6][24] ;
 wire \fifo_in.FIFO[6][25] ;
 wire \fifo_in.FIFO[6][26] ;
 wire \fifo_in.FIFO[6][27] ;
 wire \fifo_in.FIFO[6][28] ;
 wire \fifo_in.FIFO[6][29] ;
 wire \fifo_in.FIFO[6][2] ;
 wire \fifo_in.FIFO[6][30] ;
 wire \fifo_in.FIFO[6][31] ;
 wire \fifo_in.FIFO[6][3] ;
 wire \fifo_in.FIFO[6][4] ;
 wire \fifo_in.FIFO[6][5] ;
 wire \fifo_in.FIFO[6][6] ;
 wire \fifo_in.FIFO[6][7] ;
 wire \fifo_in.FIFO[6][8] ;
 wire \fifo_in.FIFO[6][9] ;
 wire \fifo_in.FIFO[7][0] ;
 wire \fifo_in.FIFO[7][10] ;
 wire \fifo_in.FIFO[7][11] ;
 wire \fifo_in.FIFO[7][12] ;
 wire \fifo_in.FIFO[7][13] ;
 wire \fifo_in.FIFO[7][14] ;
 wire \fifo_in.FIFO[7][15] ;
 wire \fifo_in.FIFO[7][16] ;
 wire \fifo_in.FIFO[7][17] ;
 wire \fifo_in.FIFO[7][18] ;
 wire \fifo_in.FIFO[7][19] ;
 wire \fifo_in.FIFO[7][1] ;
 wire \fifo_in.FIFO[7][20] ;
 wire \fifo_in.FIFO[7][21] ;
 wire \fifo_in.FIFO[7][22] ;
 wire \fifo_in.FIFO[7][23] ;
 wire \fifo_in.FIFO[7][24] ;
 wire \fifo_in.FIFO[7][25] ;
 wire \fifo_in.FIFO[7][26] ;
 wire \fifo_in.FIFO[7][27] ;
 wire \fifo_in.FIFO[7][28] ;
 wire \fifo_in.FIFO[7][29] ;
 wire \fifo_in.FIFO[7][2] ;
 wire \fifo_in.FIFO[7][30] ;
 wire \fifo_in.FIFO[7][31] ;
 wire \fifo_in.FIFO[7][3] ;
 wire \fifo_in.FIFO[7][4] ;
 wire \fifo_in.FIFO[7][5] ;
 wire \fifo_in.FIFO[7][6] ;
 wire \fifo_in.FIFO[7][7] ;
 wire \fifo_in.FIFO[7][8] ;
 wire \fifo_in.FIFO[7][9] ;
 wire \fifo_in.count[0] ;
 wire \fifo_in.count[1] ;
 wire \fifo_in.count[2] ;
 wire \fifo_in.read_addr[0] ;
 wire \fifo_in.read_addr[1] ;
 wire \fifo_in.read_addr[2] ;
 wire \fifo_in.write_addr[0] ;
 wire \fifo_in.write_addr[1] ;
 wire \fifo_in.write_addr[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__0444__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0445__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0446__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0447__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0448__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0449__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0450__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0451__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0452__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0456__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0457__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0459__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0460__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0461__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0462__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0463__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0464__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0467__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0468__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0470__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0471__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0472__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0473__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0475__S (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0479__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0480__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0482__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0488__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0489__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0490__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0491__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0495__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0496__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0499__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0500__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0503__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0504__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__S (.DIODE(_0355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0509__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0512__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__A_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0516__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0539__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0547__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0549__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0551__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0552__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0553__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0559__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0563__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__S (.DIODE(_0376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0578__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__S (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0616__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0624__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__S (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__S (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__S (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__S1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__S (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0951__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(_0354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_0376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_0355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold625_A (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _0437_ (.A(net36),
    .Y(_0349_));
 sky130_fd_sc_hd__and2_1 _0438_ (.A(net2),
    .B(net35),
    .X(_0000_));
 sky130_fd_sc_hd__and3_1 _0439_ (.A(net719),
    .B(net36),
    .C(net2),
    .X(_0350_));
 sky130_fd_sc_hd__nand3_2 _0440_ (.A(net719),
    .B(net36),
    .C(net2),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _0441_ (.A(net722),
    .B(_0350_),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_1 _0442_ (.A(net702),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_4 _0443_ (.A(net1),
    .B(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _0444_ (.A0(net555),
    .A1(net569),
    .S(net71),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0445_ (.A0(net252),
    .A1(net367),
    .S(net71),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0446_ (.A0(net106),
    .A1(net113),
    .S(net71),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0447_ (.A0(net427),
    .A1(net489),
    .S(net71),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0448_ (.A0(net510),
    .A1(net528),
    .S(net71),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0449_ (.A0(net600),
    .A1(net618),
    .S(net71),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0450_ (.A0(net200),
    .A1(net748),
    .S(net71),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0451_ (.A0(net473),
    .A1(net477),
    .S(net71),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0452_ (.A0(net101),
    .A1(net103),
    .S(net71),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0453_ (.A0(net308),
    .A1(net409),
    .S(net71),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0454_ (.A0(net461),
    .A1(net624),
    .S(net71),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0455_ (.A0(net258),
    .A1(net305),
    .S(net71),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0456_ (.A0(net151),
    .A1(net750),
    .S(net71),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0457_ (.A0(net396),
    .A1(net565),
    .S(net71),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0458_ (.A0(net116),
    .A1(net159),
    .S(net70),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0459_ (.A0(net303),
    .A1(net431),
    .S(net70),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0460_ (.A0(net503),
    .A1(net585),
    .S(net70),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0461_ (.A0(net313),
    .A1(net738),
    .S(net70),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0462_ (.A0(net247),
    .A1(net274),
    .S(net70),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0463_ (.A0(net139),
    .A1(net218),
    .S(net70),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0464_ (.A0(net456),
    .A1(net571),
    .S(net70),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0465_ (.A0(net321),
    .A1(net393),
    .S(net70),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0466_ (.A0(net424),
    .A1(net546),
    .S(net70),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0467_ (.A0(net111),
    .A1(net206),
    .S(net70),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0468_ (.A0(net123),
    .A1(net191),
    .S(net70),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0469_ (.A0(net494),
    .A1(net577),
    .S(net70),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0470_ (.A0(net318),
    .A1(net371),
    .S(net70),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0471_ (.A0(net464),
    .A1(net740),
    .S(net70),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0472_ (.A0(net126),
    .A1(net165),
    .S(net70),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0473_ (.A0(net144),
    .A1(net148),
    .S(net70),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0474_ (.A0(net255),
    .A1(net288),
    .S(net71),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0475_ (.A0(net405),
    .A1(net447),
    .S(_0354_),
    .X(_0032_));
 sky130_fd_sc_hd__or4bb_4 _0476_ (.A(net1),
    .B(_0351_),
    .C_N(\fifo_in.write_addr[2] ),
    .D_N(\fifo_in.write_addr[1] ),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _0477_ (.A0(net555),
    .A1(net559),
    .S(net87),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0478_ (.A0(net252),
    .A1(net419),
    .S(net87),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0479_ (.A0(net106),
    .A1(net270),
    .S(net87),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0480_ (.A0(net427),
    .A1(net731),
    .S(net87),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0481_ (.A0(net510),
    .A1(net516),
    .S(net87),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0482_ (.A0(net600),
    .A1(net614),
    .S(net87),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0483_ (.A0(net200),
    .A1(net353),
    .S(net87),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0484_ (.A0(net473),
    .A1(net735),
    .S(net87),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0485_ (.A0(net101),
    .A1(net118),
    .S(net87),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0486_ (.A0(net308),
    .A1(net379),
    .S(net87),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0487_ (.A0(net461),
    .A1(net475),
    .S(net87),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0488_ (.A0(net258),
    .A1(net266),
    .S(net87),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0489_ (.A0(net151),
    .A1(net179),
    .S(net87),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0490_ (.A0(net396),
    .A1(net407),
    .S(net87),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0491_ (.A0(net116),
    .A1(net130),
    .S(net87),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0492_ (.A0(net303),
    .A1(net754),
    .S(net86),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0493_ (.A0(net503),
    .A1(net756),
    .S(net86),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0494_ (.A0(net313),
    .A1(net385),
    .S(net86),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0495_ (.A0(net247),
    .A1(net292),
    .S(net86),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0496_ (.A0(net139),
    .A1(net747),
    .S(net86),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0497_ (.A0(net456),
    .A1(net507),
    .S(net86),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0498_ (.A0(net321),
    .A1(net755),
    .S(net86),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0499_ (.A0(net424),
    .A1(net752),
    .S(net86),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0500_ (.A0(net111),
    .A1(net220),
    .S(net86),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0501_ (.A0(net123),
    .A1(net153),
    .S(net86),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0502_ (.A0(net494),
    .A1(net536),
    .S(net86),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0503_ (.A0(net318),
    .A1(net753),
    .S(net86),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0504_ (.A0(net464),
    .A1(net481),
    .S(net86),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0505_ (.A0(net126),
    .A1(net163),
    .S(net86),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0506_ (.A0(net144),
    .A1(net173),
    .S(net86),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0507_ (.A0(net255),
    .A1(net262),
    .S(net86),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0508_ (.A0(net405),
    .A1(net413),
    .S(_0355_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2b_1 _0509_ (.A_N(\fifo_in.write_addr[0] ),
    .B(net95),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2b_1 _0510_ (.A_N(net95),
    .B(\fifo_in.write_addr[0] ),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_2 _0511_ (.A(_0356_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2b_1 _0512_ (.A_N(net90),
    .B(\fifo_in.write_addr[1] ),
    .X(_0359_));
 sky130_fd_sc_hd__xnor2_2 _0513_ (.A(net90),
    .B(\fifo_in.write_addr[1] ),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2b_1 _0515_ (.A_N(net88),
    .B(\fifo_in.write_addr[2] ),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2b_1 _0516_ (.A_N(\fifo_in.write_addr[2] ),
    .B(net88),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_1 _0517_ (.A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor4_1 _0518_ (.A(net1),
    .B(_0358_),
    .C(_0361_),
    .D(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21o_1 _0519_ (.A1(net646),
    .A2(_0365_),
    .B1(_0358_),
    .X(_0065_));
 sky130_fd_sc_hd__xor2_1 _0520_ (.A(_0356_),
    .B(_0360_),
    .X(_0366_));
 sky130_fd_sc_hd__a21oi_1 _0521_ (.A1(_0356_),
    .A2(_0360_),
    .B1(_0359_),
    .Y(_0367_));
 sky130_fd_sc_hd__or2_1 _0522_ (.A(_0364_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__a31o_1 _0523_ (.A1(_0358_),
    .A2(_0362_),
    .A3(_0368_),
    .B1(_0366_),
    .X(_0369_));
 sky130_fd_sc_hd__nand4_1 _0524_ (.A(_0358_),
    .B(_0362_),
    .C(_0366_),
    .D(_0368_),
    .Y(_0370_));
 sky130_fd_sc_hd__a22o_1 _0525_ (.A1(net650),
    .A2(_0365_),
    .B1(_0369_),
    .B2(_0370_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _0526_ (.A(_0364_),
    .B(_0367_),
    .Y(_0371_));
 sky130_fd_sc_hd__o221a_1 _0527_ (.A1(_0358_),
    .A2(_0361_),
    .B1(_0364_),
    .B2(_0367_),
    .C1(_0362_),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _0528_ (.A(_0371_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a21o_1 _0529_ (.A1(_0368_),
    .A2(_0371_),
    .B1(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _0530_ (.A1(net648),
    .A2(_0365_),
    .B1(_0373_),
    .B2(_0374_),
    .X(_0067_));
 sky130_fd_sc_hd__and4bb_1 _0531_ (.A_N(\fifo_in.write_addr[0] ),
    .B_N(net1),
    .C(net2),
    .D(net36),
    .X(_0375_));
 sky130_fd_sc_hd__and3b_4 _0532_ (.A_N(\fifo_in.write_addr[1] ),
    .B(_0375_),
    .C(\fifo_in.write_addr[2] ),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0533_ (.A0(net595),
    .A1(net555),
    .S(net85),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0534_ (.A0(net402),
    .A1(net252),
    .S(net85),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0535_ (.A0(net310),
    .A1(net106),
    .S(net85),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0536_ (.A0(net491),
    .A1(net427),
    .S(net85),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0537_ (.A0(net579),
    .A1(net510),
    .S(net85),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0538_ (.A0(net636),
    .A1(net600),
    .S(net85),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(net373),
    .A1(net200),
    .S(net85),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0540_ (.A0(net583),
    .A1(net473),
    .S(net85),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0541_ (.A0(net128),
    .A1(net101),
    .S(net85),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0542_ (.A0(net417),
    .A1(net308),
    .S(net85),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0543_ (.A0(net505),
    .A1(net461),
    .S(net85),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0544_ (.A0(net284),
    .A1(net258),
    .S(net85),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0545_ (.A0(net222),
    .A1(net151),
    .S(net85),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0546_ (.A0(net445),
    .A1(net396),
    .S(net85),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0547_ (.A0(net189),
    .A1(net116),
    .S(net85),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0548_ (.A0(net337),
    .A1(net303),
    .S(net84),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0549_ (.A0(net604),
    .A1(net503),
    .S(net84),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0550_ (.A0(net387),
    .A1(net313),
    .S(net84),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(net278),
    .A1(net247),
    .S(net84),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0552_ (.A0(net177),
    .A1(net139),
    .S(net84),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0553_ (.A0(net470),
    .A1(net456),
    .S(net84),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0554_ (.A0(net365),
    .A1(net321),
    .S(net84),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0555_ (.A0(net518),
    .A1(net424),
    .S(net84),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(net232),
    .A1(net111),
    .S(net84),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0557_ (.A0(net187),
    .A1(net123),
    .S(net84),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net552),
    .A1(net494),
    .S(net84),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0559_ (.A0(net329),
    .A1(net318),
    .S(net84),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(net557),
    .A1(net464),
    .S(net84),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0561_ (.A0(net214),
    .A1(net126),
    .S(net84),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0562_ (.A0(net181),
    .A1(net144),
    .S(net84),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(net282),
    .A1(net255),
    .S(net84),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0564_ (.A0(net468),
    .A1(net405),
    .S(_0376_),
    .X(_0099_));
 sky130_fd_sc_hd__and3b_2 _0565_ (.A_N(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0375_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(net626),
    .A1(net555),
    .S(net83),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0567_ (.A0(net415),
    .A1(net252),
    .S(net83),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0568_ (.A0(net136),
    .A1(net106),
    .S(net83),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0569_ (.A0(net514),
    .A1(net427),
    .S(net83),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(net550),
    .A1(net510),
    .S(net83),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0571_ (.A0(net632),
    .A1(net600),
    .S(net83),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(net453),
    .A1(net200),
    .S(net83),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0573_ (.A0(net530),
    .A1(net473),
    .S(net83),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(net120),
    .A1(net101),
    .S(net83),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0575_ (.A0(net437),
    .A1(net308),
    .S(net83),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0576_ (.A0(net642),
    .A1(net461),
    .S(net83),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0577_ (.A0(net400),
    .A1(net258),
    .S(net83),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(net195),
    .A1(net151),
    .S(net83),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(net602),
    .A1(net396),
    .S(net83),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0580_ (.A0(net161),
    .A1(net116),
    .S(net82),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0581_ (.A0(net369),
    .A1(net303),
    .S(net82),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0582_ (.A0(net608),
    .A1(net503),
    .S(net82),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0583_ (.A0(net383),
    .A1(net313),
    .S(net82),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net315),
    .A1(net247),
    .S(net82),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(net240),
    .A1(net139),
    .S(net82),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net589),
    .A1(net456),
    .S(net82),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(net361),
    .A1(net321),
    .S(_0377_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0588_ (.A0(net540),
    .A1(net424),
    .S(net82),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(net204),
    .A1(net111),
    .S(net82),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net193),
    .A1(net123),
    .S(net82),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net573),
    .A1(net494),
    .S(net82),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(net351),
    .A1(net318),
    .S(net82),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net520),
    .A1(net464),
    .S(net82),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net234),
    .A1(net126),
    .S(net82),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(net212),
    .A1(net144),
    .S(net82),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net300),
    .A1(net255),
    .S(net82),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net729),
    .A1(net405),
    .S(net83),
    .X(_0131_));
 sky130_fd_sc_hd__or4_4 _0598_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(net1),
    .D(_0351_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net555),
    .A1(net728),
    .S(net81),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net252),
    .A1(net363),
    .S(net81),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(net106),
    .A1(net745),
    .S(net81),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net427),
    .A1(net496),
    .S(net81),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0603_ (.A0(net510),
    .A1(net727),
    .S(net81),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(net600),
    .A1(net628),
    .S(net81),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(net200),
    .A1(net238),
    .S(net81),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0606_ (.A0(net473),
    .A1(net526),
    .S(net81),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(net101),
    .A1(net734),
    .S(net81),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0608_ (.A0(net308),
    .A1(net347),
    .S(net81),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0609_ (.A0(net461),
    .A1(net638),
    .S(net81),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(net258),
    .A1(net381),
    .S(net81),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0611_ (.A0(net151),
    .A1(net157),
    .S(net81),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0612_ (.A0(net396),
    .A1(net591),
    .S(net81),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0613_ (.A0(net116),
    .A1(net134),
    .S(net80),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(net303),
    .A1(net331),
    .S(net80),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0615_ (.A0(net503),
    .A1(net593),
    .S(net80),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0616_ (.A0(net313),
    .A1(net345),
    .S(net80),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(net247),
    .A1(net280),
    .S(net80),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(net139),
    .A1(net185),
    .S(net80),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(net456),
    .A1(net587),
    .S(net80),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(net321),
    .A1(net341),
    .S(net81),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(net424),
    .A1(net498),
    .S(net80),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(net111),
    .A1(net167),
    .S(net80),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(net123),
    .A1(net742),
    .S(net80),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(net494),
    .A1(net522),
    .S(net80),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0625_ (.A0(net318),
    .A1(net398),
    .S(net80),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(net464),
    .A1(net483),
    .S(net80),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(net126),
    .A1(net746),
    .S(net80),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(net144),
    .A1(net183),
    .S(net80),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(net255),
    .A1(net260),
    .S(net80),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(net405),
    .A1(net466),
    .S(_0378_),
    .X(_0163_));
 sky130_fd_sc_hd__nor3b_4 _0631_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C_N(_0375_),
    .Y(_0379_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(net597),
    .A1(net555),
    .S(net79),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(net739),
    .A1(net252),
    .S(net79),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(net294),
    .A1(net106),
    .S(net79),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(net538),
    .A1(net427),
    .S(net79),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net610),
    .A1(net510),
    .S(net79),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _0637_ (.A0(net630),
    .A1(net600),
    .S(net79),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(net236),
    .A1(net200),
    .S(net79),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(net485),
    .A1(net473),
    .S(net79),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0640_ (.A0(net108),
    .A1(net101),
    .S(net79),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _0641_ (.A0(net736),
    .A1(net308),
    .S(net79),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(net640),
    .A1(net461),
    .S(net79),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(net298),
    .A1(net258),
    .S(net79),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _0644_ (.A0(net197),
    .A1(net151),
    .S(net79),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0645_ (.A0(net606),
    .A1(net396),
    .S(net79),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net132),
    .A1(net116),
    .S(net79),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(net333),
    .A1(net303),
    .S(net78),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0648_ (.A0(net634),
    .A1(net503),
    .S(net78),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(net411),
    .A1(net313),
    .S(net78),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _0650_ (.A0(net327),
    .A1(net247),
    .S(net78),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _0651_ (.A0(net272),
    .A1(net139),
    .S(net78),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(net612),
    .A1(net456),
    .S(net78),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _0653_ (.A0(net335),
    .A1(net321),
    .S(net78),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(net544),
    .A1(net424),
    .S(net78),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(net224),
    .A1(net111),
    .S(net78),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(net226),
    .A1(net123),
    .S(net78),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _0657_ (.A0(net542),
    .A1(net494),
    .S(net78),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(net441),
    .A1(net318),
    .S(net78),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(net500),
    .A1(net464),
    .S(net78),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net210),
    .A1(net126),
    .S(net78),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(net208),
    .A1(net144),
    .S(net78),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(net276),
    .A1(net255),
    .S(net78),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _0663_ (.A0(net451),
    .A1(net405),
    .S(_0379_),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_1 _0664_ (.A1(net36),
    .A2(net2),
    .B1(net719),
    .X(_0380_));
 sky130_fd_sc_hd__and3b_1 _0665_ (.A_N(net1),
    .B(_0351_),
    .C(net720),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _0666_ (.A(net722),
    .B(_0350_),
    .X(_0381_));
 sky130_fd_sc_hd__and3b_1 _0667_ (.A_N(net1),
    .B(_0352_),
    .C(_0381_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _0668_ (.A(net702),
    .B(_0352_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_1 _0669_ (.A1(_0353_),
    .A2(net703),
    .B1(net1),
    .Y(_0198_));
 sky130_fd_sc_hd__o311a_2 _0670_ (.A1(net650),
    .A2(net646),
    .A3(net648),
    .B1(_0349_),
    .C1(net2),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(net95),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nor2_1 _0672_ (.A(net1),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__o21a_1 _0673_ (.A1(net95),
    .A2(_0383_),
    .B1(_0385_),
    .X(_0199_));
 sky130_fd_sc_hd__a21oi_1 _0674_ (.A1(net90),
    .A2(_0384_),
    .B1(net1),
    .Y(_0386_));
 sky130_fd_sc_hd__o21a_1 _0675_ (.A1(net90),
    .A2(_0384_),
    .B1(_0386_),
    .X(_0200_));
 sky130_fd_sc_hd__and3_1 _0676_ (.A(net88),
    .B(net90),
    .C(_0384_),
    .X(_0387_));
 sky130_fd_sc_hd__a21oi_1 _0677_ (.A1(net90),
    .A2(_0384_),
    .B1(net88),
    .Y(_0388_));
 sky130_fd_sc_hd__nor3_1 _0678_ (.A(net1),
    .B(_0387_),
    .C(_0388_),
    .Y(_0201_));
 sky130_fd_sc_hd__and3_2 _0679_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0375_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _0680_ (.A0(net620),
    .A1(net555),
    .S(net77),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _0681_ (.A0(net433),
    .A1(net252),
    .S(net77),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0682_ (.A0(net290),
    .A1(net106),
    .S(net77),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _0683_ (.A0(net449),
    .A1(net427),
    .S(net77),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(net561),
    .A1(net510),
    .S(net77),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0685_ (.A0(net622),
    .A1(net600),
    .S(net77),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _0686_ (.A0(net359),
    .A1(net200),
    .S(net77),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(net567),
    .A1(net473),
    .S(net77),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(net155),
    .A1(net101),
    .S(net77),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0689_ (.A0(net429),
    .A1(net308),
    .S(net77),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(net487),
    .A1(net461),
    .S(net77),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(net296),
    .A1(net258),
    .S(net77),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(net228),
    .A1(net151),
    .S(net77),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(net439),
    .A1(net396),
    .S(net77),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(net169),
    .A1(net116),
    .S(net77),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(net343),
    .A1(net303),
    .S(net76),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(net616),
    .A1(net503),
    .S(net76),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(net349),
    .A1(net313),
    .S(net76),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(net733),
    .A1(net247),
    .S(net76),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(net242),
    .A1(net139),
    .S(net76),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(net581),
    .A1(net456),
    .S(net76),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(net375),
    .A1(net321),
    .S(net76),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(net443),
    .A1(net424),
    .S(_0389_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(net230),
    .A1(net111),
    .S(net76),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(net175),
    .A1(net123),
    .S(net76),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(net532),
    .A1(net494),
    .S(net76),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0706_ (.A0(net357),
    .A1(net318),
    .S(net76),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(net563),
    .A1(net464),
    .S(net76),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(net249),
    .A1(net126),
    .S(net76),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0709_ (.A0(net732),
    .A1(net144),
    .S(net76),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(net286),
    .A1(net255),
    .S(net76),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(net435),
    .A1(net405),
    .S(net76),
    .X(_0233_));
 sky130_fd_sc_hd__or4b_4 _0712_ (.A(\fifo_in.write_addr[1] ),
    .B(net1),
    .C(_0351_),
    .D_N(\fifo_in.write_addr[2] ),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(net555),
    .A1(net575),
    .S(net74),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(net252),
    .A1(net389),
    .S(net74),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(net106),
    .A1(net268),
    .S(net74),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(net427),
    .A1(net458),
    .S(net74),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(net510),
    .A1(net534),
    .S(net74),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(net600),
    .A1(net726),
    .S(net74),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(net200),
    .A1(net355),
    .S(net74),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(net473),
    .A1(net512),
    .S(net74),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(net101),
    .A1(net216),
    .S(net74),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(net308),
    .A1(net391),
    .S(net74),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(net461),
    .A1(net741),
    .S(net74),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(net258),
    .A1(net730),
    .S(net74),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0725_ (.A0(net151),
    .A1(net244),
    .S(net74),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(net396),
    .A1(net751),
    .S(net74),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(net116),
    .A1(net749),
    .S(net74),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net303),
    .A1(net325),
    .S(net74),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(net503),
    .A1(net548),
    .S(net75),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(net313),
    .A1(net377),
    .S(net75),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(net247),
    .A1(net264),
    .S(net75),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net139),
    .A1(net171),
    .S(net75),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0733_ (.A0(net456),
    .A1(net743),
    .S(net75),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(net321),
    .A1(net323),
    .S(net75),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(net424),
    .A1(net524),
    .S(net75),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net111),
    .A1(net737),
    .S(net75),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0737_ (.A0(net123),
    .A1(net141),
    .S(net75),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net494),
    .A1(net725),
    .S(net75),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(net318),
    .A1(net339),
    .S(net75),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net464),
    .A1(net479),
    .S(net75),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(net126),
    .A1(net202),
    .S(net75),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(net144),
    .A1(net146),
    .S(net75),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(net255),
    .A1(net744),
    .S(net75),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(net405),
    .A1(net421),
    .S(net75),
    .X(_0265_));
 sky130_fd_sc_hd__nand2b_4 _0745_ (.A_N(net1),
    .B(_0383_),
    .Y(_0391_));
 sky130_fd_sc_hd__mux4_1 _0746_ (.A0(net595),
    .A1(net575),
    .A2(net620),
    .A3(net559),
    .S0(net95),
    .S1(net90),
    .X(_0392_));
 sky130_fd_sc_hd__mux4_1 _0747_ (.A0(net597),
    .A1(\fifo_in.FIFO[1][0] ),
    .A2(net626),
    .A3(net569),
    .S0(net96),
    .S1(net90),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(_0393_),
    .A1(_0392_),
    .S(net88),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _0749_ (.A0(_0394_),
    .A1(net694),
    .S(net73),
    .X(_0266_));
 sky130_fd_sc_hd__mux4_1 _0750_ (.A0(net402),
    .A1(net389),
    .A2(net433),
    .A3(net419),
    .S0(net95),
    .S1(net90),
    .X(_0395_));
 sky130_fd_sc_hd__mux4_1 _0751_ (.A0(\fifo_in.FIFO[0][1] ),
    .A1(net363),
    .A2(net415),
    .A3(net367),
    .S0(net95),
    .S1(net90),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(_0396_),
    .A1(_0395_),
    .S(net88),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _0753_ (.A0(_0397_),
    .A1(net678),
    .S(net73),
    .X(_0267_));
 sky130_fd_sc_hd__mux4_1 _0754_ (.A0(net310),
    .A1(net268),
    .A2(net290),
    .A3(net270),
    .S0(net95),
    .S1(net90),
    .X(_0398_));
 sky130_fd_sc_hd__mux4_1 _0755_ (.A0(net294),
    .A1(\fifo_in.FIFO[1][2] ),
    .A2(net136),
    .A3(net113),
    .S0(net95),
    .S1(net90),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(_0399_),
    .A1(_0398_),
    .S(net88),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _0757_ (.A0(_0400_),
    .A1(net698),
    .S(net73),
    .X(_0268_));
 sky130_fd_sc_hd__mux4_1 _0758_ (.A0(net491),
    .A1(net458),
    .A2(net449),
    .A3(\fifo_in.FIFO[7][3] ),
    .S0(net96),
    .S1(net90),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _0759_ (.A0(net538),
    .A1(net496),
    .A2(net514),
    .A3(net489),
    .S0(net95),
    .S1(net90),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(_0402_),
    .A1(_0401_),
    .S(net88),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(_0403_),
    .A1(net668),
    .S(net73),
    .X(_0269_));
 sky130_fd_sc_hd__mux4_1 _0762_ (.A0(net579),
    .A1(net534),
    .A2(net561),
    .A3(net516),
    .S0(net95),
    .S1(net91),
    .X(_0404_));
 sky130_fd_sc_hd__mux4_1 _0763_ (.A0(net610),
    .A1(\fifo_in.FIFO[1][4] ),
    .A2(net550),
    .A3(net528),
    .S0(net95),
    .S1(net91),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(_0405_),
    .A1(_0404_),
    .S(net88),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(_0406_),
    .A1(net674),
    .S(net73),
    .X(_0270_));
 sky130_fd_sc_hd__mux4_1 _0766_ (.A0(net636),
    .A1(\fifo_in.FIFO[5][5] ),
    .A2(net622),
    .A3(net614),
    .S0(net95),
    .S1(net94),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _0767_ (.A0(net630),
    .A1(net628),
    .A2(net632),
    .A3(net618),
    .S0(net95),
    .S1(net91),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(_0408_),
    .A1(_0407_),
    .S(net88),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(_0409_),
    .A1(net700),
    .S(net73),
    .X(_0271_));
 sky130_fd_sc_hd__mux4_1 _0770_ (.A0(net373),
    .A1(net355),
    .A2(net359),
    .A3(net353),
    .S0(net95),
    .S1(net90),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _0771_ (.A0(net236),
    .A1(net238),
    .A2(net453),
    .A3(\fifo_in.FIFO[3][6] ),
    .S0(net95),
    .S1(net90),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(_0411_),
    .A1(_0410_),
    .S(net88),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(_0412_),
    .A1(net692),
    .S(net73),
    .X(_0272_));
 sky130_fd_sc_hd__mux4_1 _0774_ (.A0(net583),
    .A1(net512),
    .A2(net567),
    .A3(\fifo_in.FIFO[7][7] ),
    .S0(net96),
    .S1(net91),
    .X(_0413_));
 sky130_fd_sc_hd__mux4_1 _0775_ (.A0(net485),
    .A1(net526),
    .A2(net530),
    .A3(net477),
    .S0(net96),
    .S1(net91),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(_0414_),
    .A1(_0413_),
    .S(net88),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(_0415_),
    .A1(net705),
    .S(net73),
    .X(_0273_));
 sky130_fd_sc_hd__mux4_1 _0778_ (.A0(net128),
    .A1(net216),
    .A2(net155),
    .A3(net118),
    .S0(net96),
    .S1(net91),
    .X(_0416_));
 sky130_fd_sc_hd__mux4_1 _0779_ (.A0(net108),
    .A1(\fifo_in.FIFO[1][8] ),
    .A2(net120),
    .A3(net103),
    .S0(net99),
    .S1(net91),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(_0417_),
    .A1(_0416_),
    .S(net88),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(_0418_),
    .A1(net684),
    .S(net73),
    .X(_0274_));
 sky130_fd_sc_hd__mux4_1 _0782_ (.A0(net417),
    .A1(net391),
    .A2(net429),
    .A3(net379),
    .S0(net96),
    .S1(net91),
    .X(_0419_));
 sky130_fd_sc_hd__mux4_1 _0783_ (.A0(\fifo_in.FIFO[0][9] ),
    .A1(net347),
    .A2(net437),
    .A3(net409),
    .S0(net96),
    .S1(net91),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(_0420_),
    .A1(_0419_),
    .S(net88),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(_0421_),
    .A1(net660),
    .S(net73),
    .X(_0275_));
 sky130_fd_sc_hd__mux4_1 _0786_ (.A0(net505),
    .A1(\fifo_in.FIFO[5][10] ),
    .A2(net487),
    .A3(net475),
    .S0(net96),
    .S1(net91),
    .X(_0422_));
 sky130_fd_sc_hd__mux4_1 _0787_ (.A0(net640),
    .A1(net638),
    .A2(net642),
    .A3(net624),
    .S0(net96),
    .S1(net91),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(_0423_),
    .A1(_0422_),
    .S(net88),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(_0424_),
    .A1(net713),
    .S(net73),
    .X(_0276_));
 sky130_fd_sc_hd__mux4_1 _0790_ (.A0(net284),
    .A1(\fifo_in.FIFO[5][11] ),
    .A2(net296),
    .A3(net266),
    .S0(net96),
    .S1(net91),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _0791_ (.A0(net298),
    .A1(net381),
    .A2(net400),
    .A3(net305),
    .S0(net96),
    .S1(net91),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(_0426_),
    .A1(_0425_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(_0427_),
    .A1(net670),
    .S(net73),
    .X(_0277_));
 sky130_fd_sc_hd__mux4_1 _0794_ (.A0(net222),
    .A1(net244),
    .A2(net228),
    .A3(net179),
    .S0(net96),
    .S1(net91),
    .X(_0428_));
 sky130_fd_sc_hd__mux4_1 _0795_ (.A0(net197),
    .A1(net157),
    .A2(net195),
    .A3(\fifo_in.FIFO[3][12] ),
    .S0(net96),
    .S1(net91),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(_0429_),
    .A1(_0428_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(_0430_),
    .A1(net664),
    .S(net73),
    .X(_0278_));
 sky130_fd_sc_hd__mux4_1 _0798_ (.A0(net445),
    .A1(\fifo_in.FIFO[5][13] ),
    .A2(net439),
    .A3(net407),
    .S0(net96),
    .S1(net94),
    .X(_0431_));
 sky130_fd_sc_hd__mux4_1 _0799_ (.A0(net606),
    .A1(net591),
    .A2(net602),
    .A3(net565),
    .S0(net96),
    .S1(net94),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(_0432_),
    .A1(_0431_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(_0433_),
    .A1(net711),
    .S(net73),
    .X(_0279_));
 sky130_fd_sc_hd__mux4_1 _0802_ (.A0(net189),
    .A1(\fifo_in.FIFO[5][14] ),
    .A2(net169),
    .A3(net130),
    .S0(net98),
    .S1(net93),
    .X(_0434_));
 sky130_fd_sc_hd__mux4_1 _0803_ (.A0(net132),
    .A1(net134),
    .A2(net161),
    .A3(net159),
    .S0(net98),
    .S1(net93),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(_0435_),
    .A1(_0434_),
    .S(net88),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(_0436_),
    .A1(net658),
    .S(net73),
    .X(_0280_));
 sky130_fd_sc_hd__mux4_1 _0806_ (.A0(net337),
    .A1(net325),
    .A2(net343),
    .A3(\fifo_in.FIFO[7][15] ),
    .S0(net98),
    .S1(net93),
    .X(_0298_));
 sky130_fd_sc_hd__mux4_1 _0807_ (.A0(net333),
    .A1(net331),
    .A2(net369),
    .A3(net431),
    .S0(net98),
    .S1(net93),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(_0299_),
    .A1(_0298_),
    .S(net89),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(_0300_),
    .A1(net656),
    .S(net72),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_1 _0810_ (.A0(net604),
    .A1(net548),
    .A2(net616),
    .A3(\fifo_in.FIFO[7][16] ),
    .S0(net98),
    .S1(net93),
    .X(_0301_));
 sky130_fd_sc_hd__mux4_1 _0811_ (.A0(net634),
    .A1(net593),
    .A2(net608),
    .A3(net585),
    .S0(net98),
    .S1(net93),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(_0302_),
    .A1(_0301_),
    .S(net89),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(_0303_),
    .A1(net666),
    .S(net72),
    .X(_0282_));
 sky130_fd_sc_hd__mux4_1 _0814_ (.A0(net387),
    .A1(net377),
    .A2(net349),
    .A3(net385),
    .S0(net98),
    .S1(net93),
    .X(_0304_));
 sky130_fd_sc_hd__mux4_1 _0815_ (.A0(net411),
    .A1(net345),
    .A2(net383),
    .A3(\fifo_in.FIFO[3][17] ),
    .S0(net98),
    .S1(net93),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(_0305_),
    .A1(_0304_),
    .S(net89),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _0817_ (.A0(_0306_),
    .A1(net652),
    .S(net72),
    .X(_0283_));
 sky130_fd_sc_hd__mux4_1 _0818_ (.A0(net278),
    .A1(net264),
    .A2(\fifo_in.FIFO[6][18] ),
    .A3(net292),
    .S0(net98),
    .S1(net93),
    .X(_0307_));
 sky130_fd_sc_hd__mux4_1 _0819_ (.A0(net327),
    .A1(net280),
    .A2(net315),
    .A3(net274),
    .S0(net98),
    .S1(net93),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(_0308_),
    .A1(_0307_),
    .S(net89),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _0821_ (.A0(_0309_),
    .A1(net696),
    .S(net72),
    .X(_0284_));
 sky130_fd_sc_hd__mux4_1 _0822_ (.A0(net177),
    .A1(net171),
    .A2(net242),
    .A3(\fifo_in.FIFO[7][19] ),
    .S0(net98),
    .S1(net93),
    .X(_0310_));
 sky130_fd_sc_hd__mux4_1 _0823_ (.A0(net272),
    .A1(net185),
    .A2(net240),
    .A3(net218),
    .S0(net98),
    .S1(net93),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(_0311_),
    .A1(_0310_),
    .S(net89),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(_0312_),
    .A1(net682),
    .S(net72),
    .X(_0285_));
 sky130_fd_sc_hd__mux4_1 _0826_ (.A0(net470),
    .A1(\fifo_in.FIFO[5][20] ),
    .A2(net581),
    .A3(net507),
    .S0(net98),
    .S1(net93),
    .X(_0313_));
 sky130_fd_sc_hd__mux4_1 _0827_ (.A0(net612),
    .A1(net587),
    .A2(net589),
    .A3(net571),
    .S0(net98),
    .S1(net93),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(_0314_),
    .A1(_0313_),
    .S(net89),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(_0315_),
    .A1(net717),
    .S(net72),
    .X(_0286_));
 sky130_fd_sc_hd__mux4_1 _0830_ (.A0(net365),
    .A1(net323),
    .A2(net375),
    .A3(\fifo_in.FIFO[7][21] ),
    .S0(net98),
    .S1(net93),
    .X(_0316_));
 sky130_fd_sc_hd__mux4_1 _0831_ (.A0(net335),
    .A1(net341),
    .A2(net361),
    .A3(net393),
    .S0(net98),
    .S1(net93),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(_0317_),
    .A1(_0316_),
    .S(net89),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _0833_ (.A0(_0318_),
    .A1(net662),
    .S(net72),
    .X(_0287_));
 sky130_fd_sc_hd__mux4_1 _0834_ (.A0(net518),
    .A1(net524),
    .A2(net443),
    .A3(\fifo_in.FIFO[7][22] ),
    .S0(net99),
    .S1(net92),
    .X(_0319_));
 sky130_fd_sc_hd__mux4_1 _0835_ (.A0(net544),
    .A1(net498),
    .A2(net540),
    .A3(net546),
    .S0(net97),
    .S1(net92),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _0836_ (.A0(_0320_),
    .A1(_0319_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(_0321_),
    .A1(net709),
    .S(net72),
    .X(_0288_));
 sky130_fd_sc_hd__mux4_1 _0838_ (.A0(net232),
    .A1(\fifo_in.FIFO[5][23] ),
    .A2(net230),
    .A3(net220),
    .S0(net97),
    .S1(net92),
    .X(_0322_));
 sky130_fd_sc_hd__mux4_1 _0839_ (.A0(net224),
    .A1(net167),
    .A2(net204),
    .A3(net206),
    .S0(net97),
    .S1(net92),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(_0323_),
    .A1(_0322_),
    .S(net89),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _0841_ (.A0(_0324_),
    .A1(net686),
    .S(net72),
    .X(_0289_));
 sky130_fd_sc_hd__mux4_1 _0842_ (.A0(net187),
    .A1(net141),
    .A2(net175),
    .A3(net153),
    .S0(net97),
    .S1(net92),
    .X(_0325_));
 sky130_fd_sc_hd__mux4_1 _0843_ (.A0(net226),
    .A1(\fifo_in.FIFO[1][24] ),
    .A2(net193),
    .A3(net191),
    .S0(net97),
    .S1(net92),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(_0326_),
    .A1(_0325_),
    .S(net89),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(_0327_),
    .A1(net654),
    .S(net72),
    .X(_0290_));
 sky130_fd_sc_hd__mux4_1 _0846_ (.A0(net552),
    .A1(\fifo_in.FIFO[5][25] ),
    .A2(net532),
    .A3(net536),
    .S0(net99),
    .S1(net92),
    .X(_0328_));
 sky130_fd_sc_hd__mux4_1 _0847_ (.A0(net542),
    .A1(net522),
    .A2(net573),
    .A3(net577),
    .S0(net99),
    .S1(net94),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0329_),
    .A1(_0328_),
    .S(net89),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(_0330_),
    .A1(net688),
    .S(net72),
    .X(_0291_));
 sky130_fd_sc_hd__mux4_1 _0850_ (.A0(net329),
    .A1(net339),
    .A2(net357),
    .A3(\fifo_in.FIFO[7][26] ),
    .S0(net97),
    .S1(net92),
    .X(_0331_));
 sky130_fd_sc_hd__mux4_1 _0851_ (.A0(net441),
    .A1(net398),
    .A2(net351),
    .A3(net371),
    .S0(net99),
    .S1(net94),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(_0332_),
    .A1(_0331_),
    .S(net89),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _0853_ (.A0(_0333_),
    .A1(net672),
    .S(net72),
    .X(_0292_));
 sky130_fd_sc_hd__mux4_1 _0854_ (.A0(net557),
    .A1(net479),
    .A2(net563),
    .A3(net481),
    .S0(net97),
    .S1(net92),
    .X(_0334_));
 sky130_fd_sc_hd__mux4_1 _0855_ (.A0(net500),
    .A1(net483),
    .A2(net520),
    .A3(\fifo_in.FIFO[3][27] ),
    .S0(net97),
    .S1(net92),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(_0335_),
    .A1(_0334_),
    .S(net89),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _0857_ (.A0(_0336_),
    .A1(net715),
    .S(net72),
    .X(_0293_));
 sky130_fd_sc_hd__mux4_1 _0858_ (.A0(net214),
    .A1(net202),
    .A2(net249),
    .A3(net163),
    .S0(net97),
    .S1(net92),
    .X(_0337_));
 sky130_fd_sc_hd__mux4_1 _0859_ (.A0(net210),
    .A1(\fifo_in.FIFO[1][28] ),
    .A2(net234),
    .A3(net165),
    .S0(net97),
    .S1(net92),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(_0338_),
    .A1(_0337_),
    .S(net89),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _0861_ (.A0(_0339_),
    .A1(net690),
    .S(net72),
    .X(_0294_));
 sky130_fd_sc_hd__mux4_1 _0862_ (.A0(net181),
    .A1(net146),
    .A2(\fifo_in.FIFO[6][29] ),
    .A3(net173),
    .S0(net97),
    .S1(net92),
    .X(_0340_));
 sky130_fd_sc_hd__mux4_1 _0863_ (.A0(net208),
    .A1(net183),
    .A2(net212),
    .A3(net148),
    .S0(net97),
    .S1(net92),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(_0341_),
    .A1(_0340_),
    .S(net89),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _0865_ (.A0(_0342_),
    .A1(net680),
    .S(net72),
    .X(_0295_));
 sky130_fd_sc_hd__mux4_1 _0866_ (.A0(net282),
    .A1(\fifo_in.FIFO[5][30] ),
    .A2(net286),
    .A3(net262),
    .S0(net97),
    .S1(net92),
    .X(_0343_));
 sky130_fd_sc_hd__mux4_1 _0867_ (.A0(net276),
    .A1(net260),
    .A2(net300),
    .A3(net288),
    .S0(net97),
    .S1(net92),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _0868_ (.A0(_0344_),
    .A1(_0343_),
    .S(net89),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _0869_ (.A0(_0345_),
    .A1(net676),
    .S(net72),
    .X(_0296_));
 sky130_fd_sc_hd__mux4_1 _0870_ (.A0(net468),
    .A1(net421),
    .A2(net435),
    .A3(net413),
    .S0(net97),
    .S1(net94),
    .X(_0346_));
 sky130_fd_sc_hd__mux4_1 _0871_ (.A0(net451),
    .A1(net466),
    .A2(\fifo_in.FIFO[2][31] ),
    .A3(net447),
    .S0(net97),
    .S1(net94),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _0872_ (.A0(_0347_),
    .A1(_0346_),
    .S(net89),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _0873_ (.A0(_0348_),
    .A1(net707),
    .S(_0391_),
    .X(_0297_));
 sky130_fd_sc_hd__dfxtp_1 _0874_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net645),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _0875_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net570),
    .Q(\fifo_in.FIFO[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0876_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net368),
    .Q(\fifo_in.FIFO[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0877_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net114),
    .Q(\fifo_in.FIFO[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0878_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net490),
    .Q(\fifo_in.FIFO[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0879_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net529),
    .Q(\fifo_in.FIFO[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0880_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net619),
    .Q(\fifo_in.FIFO[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0881_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net201),
    .Q(\fifo_in.FIFO[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0882_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net478),
    .Q(\fifo_in.FIFO[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0883_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net104),
    .Q(\fifo_in.FIFO[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0884_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net410),
    .Q(\fifo_in.FIFO[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0885_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net625),
    .Q(\fifo_in.FIFO[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0886_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net306),
    .Q(\fifo_in.FIFO[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0887_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net152),
    .Q(\fifo_in.FIFO[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0888_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net566),
    .Q(\fifo_in.FIFO[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0889_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net160),
    .Q(\fifo_in.FIFO[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0890_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net432),
    .Q(\fifo_in.FIFO[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0891_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net586),
    .Q(\fifo_in.FIFO[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0892_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net314),
    .Q(\fifo_in.FIFO[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0893_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net275),
    .Q(\fifo_in.FIFO[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0894_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net219),
    .Q(\fifo_in.FIFO[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0895_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net572),
    .Q(\fifo_in.FIFO[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net394),
    .Q(\fifo_in.FIFO[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net547),
    .Q(\fifo_in.FIFO[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net207),
    .Q(\fifo_in.FIFO[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net192),
    .Q(\fifo_in.FIFO[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0900_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net578),
    .Q(\fifo_in.FIFO[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net372),
    .Q(\fifo_in.FIFO[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net465),
    .Q(\fifo_in.FIFO[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net166),
    .Q(\fifo_in.FIFO[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net149),
    .Q(\fifo_in.FIFO[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net289),
    .Q(\fifo_in.FIFO[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net448),
    .Q(\fifo_in.FIFO[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net560),
    .Q(\fifo_in.FIFO[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net420),
    .Q(\fifo_in.FIFO[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net271),
    .Q(\fifo_in.FIFO[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net428),
    .Q(\fifo_in.FIFO[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net517),
    .Q(\fifo_in.FIFO[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net615),
    .Q(\fifo_in.FIFO[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net354),
    .Q(\fifo_in.FIFO[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net474),
    .Q(\fifo_in.FIFO[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0915_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net119),
    .Q(\fifo_in.FIFO[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0916_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net380),
    .Q(\fifo_in.FIFO[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0917_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net476),
    .Q(\fifo_in.FIFO[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0918_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net267),
    .Q(\fifo_in.FIFO[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0919_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net180),
    .Q(\fifo_in.FIFO[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0920_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net408),
    .Q(\fifo_in.FIFO[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0921_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net131),
    .Q(\fifo_in.FIFO[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0922_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net304),
    .Q(\fifo_in.FIFO[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net504),
    .Q(\fifo_in.FIFO[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0924_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net386),
    .Q(\fifo_in.FIFO[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0925_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net293),
    .Q(\fifo_in.FIFO[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net140),
    .Q(\fifo_in.FIFO[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net508),
    .Q(\fifo_in.FIFO[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0928_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net322),
    .Q(\fifo_in.FIFO[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net425),
    .Q(\fifo_in.FIFO[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net221),
    .Q(\fifo_in.FIFO[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0931_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net154),
    .Q(\fifo_in.FIFO[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net537),
    .Q(\fifo_in.FIFO[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net319),
    .Q(\fifo_in.FIFO[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net482),
    .Q(\fifo_in.FIFO[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net164),
    .Q(\fifo_in.FIFO[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net174),
    .Q(\fifo_in.FIFO[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net263),
    .Q(\fifo_in.FIFO[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net414),
    .Q(\fifo_in.FIFO[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net647),
    .Q(\fifo_in.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net651),
    .Q(\fifo_in.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net649),
    .Q(\fifo_in.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net596),
    .Q(\fifo_in.FIFO[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net403),
    .Q(\fifo_in.FIFO[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net311),
    .Q(\fifo_in.FIFO[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net492),
    .Q(\fifo_in.FIFO[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net580),
    .Q(\fifo_in.FIFO[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net637),
    .Q(\fifo_in.FIFO[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net374),
    .Q(\fifo_in.FIFO[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net584),
    .Q(\fifo_in.FIFO[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net129),
    .Q(\fifo_in.FIFO[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net418),
    .Q(\fifo_in.FIFO[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net506),
    .Q(\fifo_in.FIFO[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net285),
    .Q(\fifo_in.FIFO[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net223),
    .Q(\fifo_in.FIFO[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net446),
    .Q(\fifo_in.FIFO[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net190),
    .Q(\fifo_in.FIFO[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net338),
    .Q(\fifo_in.FIFO[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net605),
    .Q(\fifo_in.FIFO[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net388),
    .Q(\fifo_in.FIFO[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net279),
    .Q(\fifo_in.FIFO[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net178),
    .Q(\fifo_in.FIFO[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net471),
    .Q(\fifo_in.FIFO[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net366),
    .Q(\fifo_in.FIFO[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net519),
    .Q(\fifo_in.FIFO[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net233),
    .Q(\fifo_in.FIFO[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net188),
    .Q(\fifo_in.FIFO[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net553),
    .Q(\fifo_in.FIFO[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net330),
    .Q(\fifo_in.FIFO[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net558),
    .Q(\fifo_in.FIFO[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net215),
    .Q(\fifo_in.FIFO[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net182),
    .Q(\fifo_in.FIFO[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net283),
    .Q(\fifo_in.FIFO[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net469),
    .Q(\fifo_in.FIFO[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net627),
    .Q(\fifo_in.FIFO[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net416),
    .Q(\fifo_in.FIFO[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net137),
    .Q(\fifo_in.FIFO[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net515),
    .Q(\fifo_in.FIFO[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net551),
    .Q(\fifo_in.FIFO[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net633),
    .Q(\fifo_in.FIFO[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net454),
    .Q(\fifo_in.FIFO[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net531),
    .Q(\fifo_in.FIFO[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net121),
    .Q(\fifo_in.FIFO[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net438),
    .Q(\fifo_in.FIFO[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net643),
    .Q(\fifo_in.FIFO[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net401),
    .Q(\fifo_in.FIFO[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net196),
    .Q(\fifo_in.FIFO[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net603),
    .Q(\fifo_in.FIFO[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net162),
    .Q(\fifo_in.FIFO[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net370),
    .Q(\fifo_in.FIFO[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net609),
    .Q(\fifo_in.FIFO[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net384),
    .Q(\fifo_in.FIFO[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net316),
    .Q(\fifo_in.FIFO[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net241),
    .Q(\fifo_in.FIFO[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net590),
    .Q(\fifo_in.FIFO[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net362),
    .Q(\fifo_in.FIFO[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net541),
    .Q(\fifo_in.FIFO[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net205),
    .Q(\fifo_in.FIFO[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net194),
    .Q(\fifo_in.FIFO[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net574),
    .Q(\fifo_in.FIFO[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net352),
    .Q(\fifo_in.FIFO[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net521),
    .Q(\fifo_in.FIFO[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net235),
    .Q(\fifo_in.FIFO[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net213),
    .Q(\fifo_in.FIFO[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net301),
    .Q(\fifo_in.FIFO[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net406),
    .Q(\fifo_in.FIFO[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net556),
    .Q(\fifo_in.FIFO[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net364),
    .Q(\fifo_in.FIFO[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net107),
    .Q(\fifo_in.FIFO[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net497),
    .Q(\fifo_in.FIFO[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net511),
    .Q(\fifo_in.FIFO[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net629),
    .Q(\fifo_in.FIFO[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net239),
    .Q(\fifo_in.FIFO[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net527),
    .Q(\fifo_in.FIFO[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net102),
    .Q(\fifo_in.FIFO[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net348),
    .Q(\fifo_in.FIFO[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net639),
    .Q(\fifo_in.FIFO[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net382),
    .Q(\fifo_in.FIFO[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net158),
    .Q(\fifo_in.FIFO[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net592),
    .Q(\fifo_in.FIFO[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net135),
    .Q(\fifo_in.FIFO[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net332),
    .Q(\fifo_in.FIFO[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net594),
    .Q(\fifo_in.FIFO[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net346),
    .Q(\fifo_in.FIFO[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net281),
    .Q(\fifo_in.FIFO[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net186),
    .Q(\fifo_in.FIFO[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net588),
    .Q(\fifo_in.FIFO[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net342),
    .Q(\fifo_in.FIFO[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net499),
    .Q(\fifo_in.FIFO[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net168),
    .Q(\fifo_in.FIFO[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net124),
    .Q(\fifo_in.FIFO[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net523),
    .Q(\fifo_in.FIFO[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net399),
    .Q(\fifo_in.FIFO[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net484),
    .Q(\fifo_in.FIFO[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net127),
    .Q(\fifo_in.FIFO[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net184),
    .Q(\fifo_in.FIFO[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net261),
    .Q(\fifo_in.FIFO[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net467),
    .Q(\fifo_in.FIFO[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net598),
    .Q(\fifo_in.FIFO[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net253),
    .Q(\fifo_in.FIFO[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net295),
    .Q(\fifo_in.FIFO[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net539),
    .Q(\fifo_in.FIFO[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net611),
    .Q(\fifo_in.FIFO[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net631),
    .Q(\fifo_in.FIFO[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net237),
    .Q(\fifo_in.FIFO[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net486),
    .Q(\fifo_in.FIFO[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net109),
    .Q(\fifo_in.FIFO[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net309),
    .Q(\fifo_in.FIFO[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net641),
    .Q(\fifo_in.FIFO[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net299),
    .Q(\fifo_in.FIFO[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net198),
    .Q(\fifo_in.FIFO[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net607),
    .Q(\fifo_in.FIFO[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net133),
    .Q(\fifo_in.FIFO[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net334),
    .Q(\fifo_in.FIFO[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net635),
    .Q(\fifo_in.FIFO[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net412),
    .Q(\fifo_in.FIFO[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net328),
    .Q(\fifo_in.FIFO[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net273),
    .Q(\fifo_in.FIFO[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net613),
    .Q(\fifo_in.FIFO[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net336),
    .Q(\fifo_in.FIFO[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net545),
    .Q(\fifo_in.FIFO[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net225),
    .Q(\fifo_in.FIFO[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net227),
    .Q(\fifo_in.FIFO[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net543),
    .Q(\fifo_in.FIFO[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net442),
    .Q(\fifo_in.FIFO[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net501),
    .Q(\fifo_in.FIFO[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net211),
    .Q(\fifo_in.FIFO[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net209),
    .Q(\fifo_in.FIFO[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net277),
    .Q(\fifo_in.FIFO[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net452),
    .Q(\fifo_in.FIFO[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net721),
    .Q(\fifo_in.write_addr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1071_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0197_),
    .Q(\fifo_in.write_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1072_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net704),
    .Q(\fifo_in.write_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0199_),
    .Q(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0200_),
    .Q(\fifo_in.read_addr[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1075_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0201_),
    .Q(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net621),
    .Q(\fifo_in.FIFO[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net434),
    .Q(\fifo_in.FIFO[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net291),
    .Q(\fifo_in.FIFO[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net450),
    .Q(\fifo_in.FIFO[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net562),
    .Q(\fifo_in.FIFO[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net623),
    .Q(\fifo_in.FIFO[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net360),
    .Q(\fifo_in.FIFO[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net568),
    .Q(\fifo_in.FIFO[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net156),
    .Q(\fifo_in.FIFO[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net430),
    .Q(\fifo_in.FIFO[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net488),
    .Q(\fifo_in.FIFO[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net297),
    .Q(\fifo_in.FIFO[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net229),
    .Q(\fifo_in.FIFO[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net440),
    .Q(\fifo_in.FIFO[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net170),
    .Q(\fifo_in.FIFO[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net344),
    .Q(\fifo_in.FIFO[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net617),
    .Q(\fifo_in.FIFO[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net350),
    .Q(\fifo_in.FIFO[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net248),
    .Q(\fifo_in.FIFO[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net243),
    .Q(\fifo_in.FIFO[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net582),
    .Q(\fifo_in.FIFO[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net376),
    .Q(\fifo_in.FIFO[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net444),
    .Q(\fifo_in.FIFO[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net231),
    .Q(\fifo_in.FIFO[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net176),
    .Q(\fifo_in.FIFO[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net533),
    .Q(\fifo_in.FIFO[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net358),
    .Q(\fifo_in.FIFO[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net564),
    .Q(\fifo_in.FIFO[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net250),
    .Q(\fifo_in.FIFO[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net145),
    .Q(\fifo_in.FIFO[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net287),
    .Q(\fifo_in.FIFO[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net436),
    .Q(\fifo_in.FIFO[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net576),
    .Q(\fifo_in.FIFO[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net390),
    .Q(\fifo_in.FIFO[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net269),
    .Q(\fifo_in.FIFO[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net459),
    .Q(\fifo_in.FIFO[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net535),
    .Q(\fifo_in.FIFO[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net601),
    .Q(\fifo_in.FIFO[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net356),
    .Q(\fifo_in.FIFO[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net513),
    .Q(\fifo_in.FIFO[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net217),
    .Q(\fifo_in.FIFO[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net392),
    .Q(\fifo_in.FIFO[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net462),
    .Q(\fifo_in.FIFO[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net259),
    .Q(\fifo_in.FIFO[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net245),
    .Q(\fifo_in.FIFO[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net397),
    .Q(\fifo_in.FIFO[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net117),
    .Q(\fifo_in.FIFO[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net326),
    .Q(\fifo_in.FIFO[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net549),
    .Q(\fifo_in.FIFO[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net378),
    .Q(\fifo_in.FIFO[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net265),
    .Q(\fifo_in.FIFO[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net172),
    .Q(\fifo_in.FIFO[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net457),
    .Q(\fifo_in.FIFO[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net324),
    .Q(\fifo_in.FIFO[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net525),
    .Q(\fifo_in.FIFO[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net112),
    .Q(\fifo_in.FIFO[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net142),
    .Q(\fifo_in.FIFO[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net495),
    .Q(\fifo_in.FIFO[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net340),
    .Q(\fifo_in.FIFO[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net480),
    .Q(\fifo_in.FIFO[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net203),
    .Q(\fifo_in.FIFO[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net147),
    .Q(\fifo_in.FIFO[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net256),
    .Q(\fifo_in.FIFO[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net422),
    .Q(\fifo_in.FIFO[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net695),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net679),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net699),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net669),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net675),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net701),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net693),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net706),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net685),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net661),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net714),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net671),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net665),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net712),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net659),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net657),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net667),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net653),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net697),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net683),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net718),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net663),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net710),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net687),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net655),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net689),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net673),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net716),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net691),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net681),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net677),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net708),
    .Q(net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_8 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_8 fanout71 (.A(_0354_),
    .X(net71));
 sky130_fd_sc_hd__buf_6 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_0391_),
    .X(net73));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(_0390_),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(_0390_),
    .X(net75));
 sky130_fd_sc_hd__buf_8 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_8 fanout77 (.A(_0389_),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(_0379_),
    .X(net79));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout81 (.A(_0378_),
    .X(net81));
 sky130_fd_sc_hd__buf_8 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(_0377_),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_8 fanout85 (.A(_0376_),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_8 fanout87 (.A(_0355_),
    .X(net87));
 sky130_fd_sc_hd__buf_6 fanout88 (.A(net724),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(\fifo_in.read_addr[2] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout91 (.A(net94),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_8 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(\fifo_in.read_addr[1] ),
    .X(net94));
 sky130_fd_sc_hd__buf_6 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(net99),
    .X(net96));
 sky130_fd_sc_hd__buf_8 fanout97 (.A(net99),
    .X(net97));
 sky130_fd_sc_hd__buf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(\fifo_in.read_addr[0] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wbs_dat_i[8]),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0172_),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(wbs_dat_i[6]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 hold101 (.A(net31),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0007_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\fifo_in.FIFO[5][28] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0262_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\fifo_in.FIFO[2][23] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0123_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\fifo_in.FIFO[3][23] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0024_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\fifo_in.FIFO[0][29] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(wbs_dat_i[23]),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0193_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\fifo_in.FIFO[0][28] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0192_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\fifo_in.FIFO[2][29] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0129_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\fifo_in.FIFO[4][28] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0096_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\fifo_in.FIFO[5][8] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0242_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\fifo_in.FIFO[3][19] ),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 hold12 (.A(net18),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0020_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\fifo_in.FIFO[7][23] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0056_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\fifo_in.FIFO[4][12] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0080_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\fifo_in.FIFO[0][23] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0187_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\fifo_in.FIFO[0][24] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0188_),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\fifo_in.FIFO[6][12] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0257_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0214_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\fifo_in.FIFO[6][23] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0225_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\fifo_in.FIFO[4][23] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0091_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\fifo_in.FIFO[2][28] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0128_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\fifo_in.FIFO[0][6] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0170_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\fifo_in.FIFO[1][6] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\fifo_in.FIFO[3][2] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0138_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\fifo_in.FIFO[2][19] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0119_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\fifo_in.FIFO[6][19] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0221_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\fifo_in.FIFO[5][12] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0246_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(wbs_dat_i[18]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 hold148 (.A(net12),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0220_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0003_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\fifo_in.FIFO[6][28] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0230_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(wbs_dat_i[1]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 hold153 (.A(net14),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0165_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(wbs_dat_i[30]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 hold156 (.A(net26),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0264_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(wbs_dat_i[11]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 hold159 (.A(net5),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(wbs_dat_i[14]),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0245_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\fifo_in.FIFO[1][30] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0162_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\fifo_in.FIFO[7][30] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0063_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\fifo_in.FIFO[5][18] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0252_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\fifo_in.FIFO[7][11] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0044_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\fifo_in.FIFO[5][2] ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 hold17 (.A(net8),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0236_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\fifo_in.FIFO[7][2] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0035_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\fifo_in.FIFO[0][19] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0183_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\fifo_in.FIFO[3][18] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0019_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\fifo_in.FIFO[0][30] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0194_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\fifo_in.FIFO[4][18] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0248_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0086_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\fifo_in.FIFO[1][18] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0150_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\fifo_in.FIFO[4][30] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0098_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\fifo_in.FIFO[4][11] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0079_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\fifo_in.FIFO[6][30] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0232_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\fifo_in.FIFO[3][30] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\fifo_in.FIFO[7][8] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0031_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\fifo_in.FIFO[6][2] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0204_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\fifo_in.FIFO[7][18] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0051_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\fifo_in.FIFO[0][2] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0166_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\fifo_in.FIFO[6][11] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0213_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\fifo_in.FIFO[0][11] ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 hold2 (.A(net33),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0041_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0175_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\fifo_in.FIFO[2][30] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0130_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(wbs_dat_i[15]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 hold204 (.A(net9),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0048_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\fifo_in.FIFO[3][11] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0012_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(wbs_dat_i[9]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 hold209 (.A(net34),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\fifo_in.FIFO[2][8] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0173_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\fifo_in.FIFO[4][2] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0070_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(wbs_dat_i[17]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 hold214 (.A(net11),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0018_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\fifo_in.FIFO[2][18] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0118_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(wbs_dat_i[26]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 hold219 (.A(net21),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0108_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0059_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(wbs_dat_i[21]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 hold222 (.A(net16),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0054_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\fifo_in.FIFO[5][21] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0255_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\fifo_in.FIFO[5][15] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0249_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\fifo_in.FIFO[0][18] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0182_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(wbs_dat_i[24]),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\fifo_in.FIFO[4][26] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0094_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\fifo_in.FIFO[1][15] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0147_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\fifo_in.FIFO[0][15] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0179_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\fifo_in.FIFO[0][21] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0185_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\fifo_in.FIFO[4][15] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0083_),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 hold24 (.A(net19),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\fifo_in.FIFO[5][26] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0260_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\fifo_in.FIFO[1][21] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0153_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\fifo_in.FIFO[6][15] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0217_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\fifo_in.FIFO[1][17] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_0149_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\fifo_in.FIFO[1][9] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0141_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0156_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\fifo_in.FIFO[6][17] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0219_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\fifo_in.FIFO[2][26] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0126_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\fifo_in.FIFO[7][6] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0039_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\fifo_in.FIFO[5][6] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0240_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\fifo_in.FIFO[6][26] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0228_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(wbs_dat_i[28]),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\fifo_in.FIFO[6][6] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0208_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\fifo_in.FIFO[2][21] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0121_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\fifo_in.FIFO[1][1] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0133_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\fifo_in.FIFO[4][21] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0089_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\fifo_in.FIFO[3][1] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0002_),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 hold27 (.A(net23),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\fifo_in.FIFO[2][15] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0115_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\fifo_in.FIFO[3][26] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0027_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\fifo_in.FIFO[4][6] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0074_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\fifo_in.FIFO[6][21] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0223_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\fifo_in.FIFO[5][17] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0251_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0160_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\fifo_in.FIFO[7][9] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0042_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\fifo_in.FIFO[1][11] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0143_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\fifo_in.FIFO[2][17] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0117_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\fifo_in.FIFO[7][17] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0050_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\fifo_in.FIFO[4][17] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0085_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fifo_in.FIFO[4][8] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\fifo_in.FIFO[5][1] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0235_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\fifo_in.FIFO[5][9] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0243_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\fifo_in.FIFO[3][21] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0022_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(wbs_dat_i[13]),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 hold297 (.A(net7),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0247_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\fifo_in.FIFO[1][26] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0140_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0076_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0158_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\fifo_in.FIFO[2][11] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0111_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\fifo_in.FIFO[4][1] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0069_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(wbs_dat_i[31]),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 hold306 (.A(net27),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0131_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\fifo_in.FIFO[7][13] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0046_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\fifo_in.FIFO[7][14] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\fifo_in.FIFO[3][9] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0010_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\fifo_in.FIFO[0][17] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0181_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\fifo_in.FIFO[7][31] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0064_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\fifo_in.FIFO[2][1] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0101_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\fifo_in.FIFO[4][9] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0077_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0047_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\fifo_in.FIFO[7][1] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0034_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\fifo_in.FIFO[5][31] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0265_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(wbs_dat_i[22]),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 hold325 (.A(net17),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0055_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(wbs_dat_i[3]),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 hold328 (.A(net28),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0036_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fifo_in.FIFO[0][14] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\fifo_in.FIFO[6][9] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0211_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\fifo_in.FIFO[3][15] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0016_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\fifo_in.FIFO[6][1] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0203_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\fifo_in.FIFO[6][31] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0233_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\fifo_in.FIFO[2][9] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0109_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0178_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\fifo_in.FIFO[6][13] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0215_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\fifo_in.FIFO[0][26] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_0190_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\fifo_in.FIFO[6][22] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0224_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\fifo_in.FIFO[4][13] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0081_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\fifo_in.FIFO[3][31] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0032_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\fifo_in.FIFO[1][14] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\fifo_in.FIFO[6][3] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_0205_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\fifo_in.FIFO[0][31] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_0195_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\fifo_in.FIFO[2][6] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0106_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(wbs_dat_i[20]),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 hold357 (.A(net15),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0254_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\fifo_in.FIFO[5][3] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0146_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0237_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(wbs_dat_i[10]),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 hold362 (.A(net4),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0244_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(wbs_dat_i[27]),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 hold365 (.A(net22),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0028_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\fifo_in.FIFO[1][31] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0163_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\fifo_in.FIFO[4][31] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\fifo_in.FIFO[2][2] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0099_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\fifo_in.FIFO[4][20] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0088_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(wbs_dat_i[7]),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_2 hold374 (.A(net32),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_0040_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\fifo_in.FIFO[7][10] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_0043_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\fifo_in.FIFO[3][7] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_0008_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0102_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\fifo_in.FIFO[5][27] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0261_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\fifo_in.FIFO[7][27] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0060_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\fifo_in.FIFO[1][27] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0159_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\fifo_in.FIFO[0][7] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_0171_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\fifo_in.FIFO[6][10] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_0212_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(wbs_dat_i[19]),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\fifo_in.FIFO[3][3] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0004_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\fifo_in.FIFO[4][3] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0071_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(wbs_dat_i[25]),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_2 hold395 (.A(net20),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0259_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\fifo_in.FIFO[1][3] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0135_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\fifo_in.FIFO[1][22] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\fifo_in.FIFO[3][8] ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 hold40 (.A(net13),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0154_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\fifo_in.FIFO[0][27] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0191_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(wbs_dat_i[16]),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_2 hold404 (.A(net10),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0049_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\fifo_in.FIFO[4][10] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0078_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\fifo_in.FIFO[7][20] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_0053_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0052_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(wbs_dat_i[4]),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_2 hold411 (.A(net29),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0136_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\fifo_in.FIFO[5][7] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0241_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\fifo_in.FIFO[2][3] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0103_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\fifo_in.FIFO[7][4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0037_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\fifo_in.FIFO[4][22] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\fifo_in.FIFO[5][24] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0090_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\fifo_in.FIFO[2][27] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0127_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\fifo_in.FIFO[1][25] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0157_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\fifo_in.FIFO[5][22] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0256_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\fifo_in.FIFO[1][7] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0139_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\fifo_in.FIFO[3][4] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0258_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0005_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\fifo_in.FIFO[2][7] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0107_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\fifo_in.FIFO[6][25] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0227_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\fifo_in.FIFO[5][4] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0238_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\fifo_in.FIFO[7][25] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0058_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\fifo_in.FIFO[0][3] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(wbs_dat_i[29]),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0167_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\fifo_in.FIFO[2][22] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0122_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\fifo_in.FIFO[0][25] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0189_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\fifo_in.FIFO[0][22] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0186_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\fifo_in.FIFO[3][22] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0023_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\fifo_in.FIFO[5][16] ),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_2 hold45 (.A(net24),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0250_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\fifo_in.FIFO[2][4] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0104_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\fifo_in.FIFO[4][25] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0093_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(wbs_dat_i[0]),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_2 hold456 (.A(net3),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_0132_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\fifo_in.FIFO[4][27] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_0095_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0231_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\fifo_in.FIFO[7][0] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0033_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\fifo_in.FIFO[6][4] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_0206_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\fifo_in.FIFO[6][27] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0229_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\fifo_in.FIFO[3][13] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0014_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\fifo_in.FIFO[6][7] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_0209_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\fifo_in.FIFO[5][29] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\fifo_in.FIFO[3][0] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0001_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\fifo_in.FIFO[3][20] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0021_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\fifo_in.FIFO[2][25] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0125_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\fifo_in.FIFO[5][0] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0234_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\fifo_in.FIFO[3][25] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0026_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0263_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\fifo_in.FIFO[4][4] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0072_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\fifo_in.FIFO[6][20] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0222_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\fifo_in.FIFO[4][7] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0075_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\fifo_in.FIFO[3][16] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0017_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\fifo_in.FIFO[1][20] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0152_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\fifo_in.FIFO[3][29] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\fifo_in.FIFO[2][20] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0120_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\fifo_in.FIFO[1][13] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0145_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\fifo_in.FIFO[1][16] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0148_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\fifo_in.FIFO[4][0] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0068_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\fifo_in.FIFO[0][0] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0164_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0009_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0030_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(wbs_dat_i[5]),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_2 hold501 (.A(net30),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0239_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\fifo_in.FIFO[2][13] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0113_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\fifo_in.FIFO[4][16] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0084_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\fifo_in.FIFO[0][13] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0177_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\fifo_in.FIFO[2][16] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(wbs_dat_i[12]),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0116_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\fifo_in.FIFO[0][4] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0168_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\fifo_in.FIFO[0][20] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0184_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\fifo_in.FIFO[7][5] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0038_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\fifo_in.FIFO[6][16] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0218_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\fifo_in.FIFO[3][5] ),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 hold52 (.A(net6),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0006_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\fifo_in.FIFO[6][0] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0202_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\fifo_in.FIFO[6][5] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0207_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\fifo_in.FIFO[3][10] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0011_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\fifo_in.FIFO[2][0] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0100_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\fifo_in.FIFO[1][5] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0013_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0137_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\fifo_in.FIFO[0][5] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0169_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\fifo_in.FIFO[2][5] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0105_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\fifo_in.FIFO[0][16] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0180_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\fifo_in.FIFO[4][5] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0073_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\fifo_in.FIFO[1][10] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\fifo_in.FIFO[7][24] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0142_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\fifo_in.FIFO[0][10] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0174_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\fifo_in.FIFO[2][10] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0110_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(wbs_cyc_i),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0000_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\fifo_in.count[0] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0065_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\fifo_in.count[2] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0057_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0067_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\fifo_in.count[1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0066_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net46),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0283_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(net54),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0290_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(net44),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0281_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net43),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\fifo_in.FIFO[6][8] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0280_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net69),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0275_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(net51),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0287_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net41),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0278_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(net45),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0282_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(net63),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0210_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0269_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(net40),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0277_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(net56),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0292_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net64),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0270_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(net61),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0296_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net49),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\fifo_in.FIFO[1][12] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0267_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net59),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0295_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net48),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0285_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(net68),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0274_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(net53),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0289_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(net55),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0144_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0291_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net58),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0294_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(net66),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0272_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net38),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0266_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net47),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0284_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(net60),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(wbs_dat_i[2]),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\fifo_in.FIFO[3][14] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0268_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(net65),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0271_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\fifo_in.write_addr[2] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0382_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_0198_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net67),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_0273_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(net62),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_0297_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0015_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net52),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_0288_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net42),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_0279_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(net39),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_0276_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net57),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_0293_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(net50),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_0286_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\fifo_in.FIFO[2][14] ),
    .X(net161));
 sky130_fd_sc_hd__buf_1 hold620 (.A(\fifo_in.write_addr[0] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(_0380_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0196_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\fifo_in.write_addr[1] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(wbs_we_i),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\fifo_in.read_addr[2] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\fifo_in.FIFO[5][25] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\fifo_in.FIFO[5][5] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\fifo_in.FIFO[1][4] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\fifo_in.FIFO[1][0] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0114_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\fifo_in.FIFO[2][31] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\fifo_in.FIFO[5][11] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\fifo_in.FIFO[7][3] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\fifo_in.FIFO[6][29] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\fifo_in.FIFO[6][18] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\fifo_in.FIFO[1][8] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\fifo_in.FIFO[7][7] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\fifo_in.FIFO[0][9] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\fifo_in.FIFO[5][23] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\fifo_in.FIFO[3][17] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\fifo_in.FIFO[7][28] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\fifo_in.FIFO[0][1] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\fifo_in.FIFO[3][27] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\fifo_in.FIFO[5][10] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\fifo_in.FIFO[1][24] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\fifo_in.FIFO[5][20] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\fifo_in.FIFO[5][30] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\fifo_in.FIFO[1][2] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\fifo_in.FIFO[1][28] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\fifo_in.FIFO[7][19] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\fifo_in.FIFO[3][6] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0061_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\fifo_in.FIFO[5][14] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\fifo_in.FIFO[3][12] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\fifo_in.FIFO[5][13] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\fifo_in.FIFO[7][22] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\fifo_in.FIFO[7][26] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\fifo_in.FIFO[7][15] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\fifo_in.FIFO[7][21] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\fifo_in.FIFO[7][16] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\fifo_in.FIFO[3][28] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0029_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\fifo_in.FIFO[1][23] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0155_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 hold7 (.A(net25),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\fifo_in.FIFO[6][14] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0216_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\fifo_in.FIFO[5][19] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0253_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\fifo_in.FIFO[7][29] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0062_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\fifo_in.FIFO[6][24] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0226_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\fifo_in.FIFO[4][19] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0087_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0134_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\fifo_in.FIFO[7][12] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0045_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\fifo_in.FIFO[4][29] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0097_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\fifo_in.FIFO[1][29] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0161_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\fifo_in.FIFO[1][19] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0151_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\fifo_in.FIFO[4][24] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0092_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fifo_in.FIFO[0][8] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\fifo_in.FIFO[4][14] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0082_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\fifo_in.FIFO[3][24] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0025_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\fifo_in.FIFO[2][24] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0124_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\fifo_in.FIFO[2][12] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0112_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\fifo_in.FIFO[0][12] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0176_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net502),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net312),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net246),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net138),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(net251),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net455),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net320),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net423),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net110),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(net122),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(net644),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(net493),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(net317),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(net463),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net125),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(net143),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(net105),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(net254),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net404),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net426),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(net509),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net554),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net599),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net199),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(net472),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(net100),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(net307),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(wbs_stb_i),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(net723),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net460),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net257),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net150),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net395),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net115),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net302),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wbs_dat_o[9]));
endmodule

